-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive := 8;
            DATA_LENGTH:  positive := 13);
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0));

end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin
	bank <= (
		0 => "0000100101110",
		1 => "0000010111000",
		141 => "0000010100001",
		6 => "0000000000110",
		85 => "0000000011000",
		206 => "0000010101010",
		35 => "0000001001101",
		138 => "0000000101111",
		220 => "0000100101111",
		137 => "0000011011000",
		13 => "0000001110101",
		14 => "0000001000110",
		207 => "0000011000000",
		16 => "0000010010000",
		252 => "0000001110100",
		19 => "0000001110011",
		192 => "0000000100110",
		20 => "0000000110000",
		21 => "0000001001011",
		111 => "0000100101010",
		23 => "0000001001111",
		24 => "0000010011101",
		25 => "0000000001101",
		26 => "0000001001000",
		27 => "0000001111100",
		28 => "0000000000111",
		29 => "0000011110100",
		30 => "0000010100110",
		31 => "0000001001100",
		32 => "0000001111000",
		34 => "0000001110111",
		36 => "0000010110010",
		37 => "0000001101010",
		38 => "0000001110110",
		5 => "0000001101000",
		56 => "0000011100010",
		41 => "0000100010111",
		43 => "0000100010100",
		44 => "0000010000000",
		45 => "0000010010100",
		39 => "0000001011011",
		48 => "0000000100001",
		49 => "0000000111000",
		253 => "0000001111110",
		52 => "0000000010110",
		255 => "0000000011010",
		119 => "0000000010111",
		148 => "0000000101110",
		55 => "0000011110111",
		40 => "0000101010011",
		214 => "0000101000111",
		59 => "0000010000001",
		60 => "0000000001110",
		61 => "0000001000000",
		62 => "0000100001111",
		58 => "0000010010011",
		178 => "0000011110010",
		64 => "0000001010101",
		65 => "0000010100000",
		67 => "0000001111101",
		128 => "0000000100111",
		63 => "0000011011010",
		69 => "0000100100111",
		71 => "0000010010111",
		72 => "0000010101101",
		73 => "0000001100110",
		74 => "0000010001110",
		70 => "0000010111110",
		78 => "0000010001111",
		3 => "0000010101110",
		80 => "0000010011011",
		82 => "0000001100111",
		83 => "0000010100101",
		84 => "0000100111111",
		86 => "0000011101001",
		33 => "0000010110001",
		143 => "0000000000100",
		89 => "0000011001101",
		204 => "0000000101010",
		90 => "0000100111010",
		91 => "0000000011100",
		92 => "0000001010110",
		94 => "0000000100010",
		248 => "0000001010000",
		96 => "0000000011110",
		177 => "0000011001000",
		98 => "0000011100101",
		99 => "0000000010010",
		100 => "0000000001001",
		101 => "0000100011101",
		2 => "0000010111111",
		103 => "0000000110110",
		66 => "0000010110000",
		238 => "0000000111110",
		105 => "0000100101100",
		108 => "0000010001010",
		109 => "0000000010001",
		110 => "0000010010001",
		68 => "0000010001101",
		113 => "0000100000010",
		114 => "0000010000011",
		156 => "0000001101100",
		115 => "0000011011111",
		116 => "0000010111011",
		118 => "0000011111111",
		102 => "0000011000010",
		120 => "0000010010010",
		121 => "0000000001010",
		87 => "0000000011001",
		122 => "0000010100010",
		123 => "0000011100111",
		125 => "0000011111010",
		57 => "0000000100110",
		127 => "0000011100100",
		147 => "0000000011000",
		112 => "0000010111010",
		129 => "0000000100101",
		131 => "0000101001100",
		132 => "0000100100101",
		209 => "0000001101011",
		133 => "0000010101100",
		134 => "0000000001011",
		229 => "0000001001001",
		135 => "0000011110000",
		230 => "0000000010100",
		198 => "0000010000101",
		53 => "0000001111010",
		54 => "0000001111111",
		190 => "0000000110011",
		139 => "0000010011000",
		140 => "0000101011000",
		166 => "0000001100101",
		186 => "0000011101011",
		142 => "0000000101000",
		88 => "0000010100100",
		232 => "0000010001001",
		191 => "0000100001010",
		145 => "0000000011101",
		146 => "0000000011011",
		81 => "0000011001100",
		97 => "0000010010110",
		149 => "0000000101101",
		151 => "0000001101111",
		203 => "0000000110100",
		152 => "0000000001100",
		153 => "0000000000101",
		154 => "0000101000001",
		155 => "0000001001110",
		107 => "0000000101011",
		157 => "0000100010001",
		237 => "0000100000011",
		160 => "0000100000110",
		162 => "0000010010101",
		164 => "0000101001001",
		165 => "0000100110001",
		159 => "0000001011100",
		216 => "0000010000010",
		167 => "0000001000001",
		179 => "0000100110101",
		168 => "0000001010010",
		169 => "0000000010101",
		170 => "0000100001100",
		77 => "0000011010011",
		171 => "0000010101001",
		172 => "0000010110110",
		215 => "0000100100010",
		173 => "0000001011101",
		174 => "0000101000110",
		176 => "0000000110101",
		9 => "0000011001010",
		76 => "0000010011111",
		163 => "0000001011110",
		243 => "0000100110111",
		180 => "0000100011001",
		181 => "0000011001001",
		182 => "0000011010110",
		242 => "0000000011111",
		183 => "0000010110101",
		184 => "0000011101101",
		150 => "0000000110111",
		17 => "0000010000100",
		187 => "0000000010011",
		201 => "0000100101000",
		188 => "0000001011111",
		189 => "0000011000100",
		11 => "0000011001111",
		79 => "0000011010000",
		75 => "0000000110010",
		193 => "0000010011110",
		194 => "0000100011011",
		235 => "0000010110100",
		195 => "0000001000011",
		196 => "0000000101001",
		197 => "0000011111101",
		130 => "0000011000110",
		199 => "0000000111111",
		212 => "0000010101111",
		200 => "0000001110001",
		124 => "0000000001000",
		95 => "0000010111100",
		136 => "0000000111001",
		18 => "0000000111010",
		205 => "0000001000101",
		104 => "0000001101110",
		15 => "0000000111011",
		208 => "0000000010000",
		161 => "0000000100000",
		210 => "0000000101100",
		211 => "0000011000111",
		106 => "0000100011111",
		213 => "0000010111101",
		4 => "0000010101011",
		185 => "0000100101101",
		42 => "0000011001011",
		217 => "0000010001011",
		244 => "0000101001111",
		219 => "0000001011000",
		10 => "0000100101011",
		50 => "0000000100100",
		222 => "0000100110010",
		223 => "0000001010001",
		224 => "0000001101001",
		225 => "0000010110111",
		226 => "0000010100111",
		202 => "0000000011010",
		227 => "0000001000100",
		228 => "0000010011001",
		12 => "0000000100010",
		51 => "0000100011110",
		231 => "0000011011011",
		144 => "0000000111101",
		233 => "0000010001000",
		234 => "0000101000011",
		218 => "0000000011111",
		236 => "0000100111100",
		93 => "0000001111011",
		175 => "0000010101000",
		239 => "0000001110010",
		221 => "0000100000111",
		240 => "0000001100000",
		241 => "0000001110000",
		47 => "0000010111001",
		22 => "0000000111100",
		158 => "0000011000011",
		245 => "0000010000110",
		246 => "0000000100011",
		247 => "0000000001111",
		117 => "0000001010100",
		249 => "0000001011010",
		250 => "0000000110001",
		126 => "0000100110000",
		251 => "0000100100001",
		46 => "0000001000111",
		8 => "0000001100001",
		254 => "0000001100011",
		7 => "0000011011101",
		others => (others => '0')
	);

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
