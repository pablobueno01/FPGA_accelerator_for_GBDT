-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive := 8;
            DATA_LENGTH:  positive := 13);
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0));

end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin
	bank <= (
		0 => "0000100101110",
		1 => "0000010111000",
		2 => "0000010100001",
		3 => "0000000000110",
		4 => "0000000011000",
		5 => "0000010101010",
		6 => "0000001001101",
		7 => "0000000101111",
		8 => "0000100101111",
		9 => "0000011011000",
		10 => "0000001110101",
		11 => "0000001000110",
		12 => "0000011000000",
		13 => "0000010010000",
		14 => "0000001110100",
		15 => "0000001110011",
		16 => "0000000100110",
		17 => "0000000110000",
		18 => "0000001001011",
		19 => "0000100101010",
		20 => "0000001001111",
		21 => "0000010011101",
		22 => "0000000001101",
		23 => "0000001001000",
		24 => "0000001111100",
		25 => "0000000000111",
		26 => "0000011110100",
		27 => "0000010100110",
		28 => "0000001001100",
		29 => "0000001111000",
		30 => "0000001110111",
		31 => "0000010110010",
		32 => "0000001101010",
		33 => "0000001110110",
		34 => "0000001101000",
		35 => "0000011100010",
		36 => "0000100010111",
		37 => "0000100010100",
		38 => "0000010000000",
		39 => "0000010010100",
		40 => "0000001011011",
		41 => "0000000100001",
		42 => "0000000111000",
		43 => "0000001111110",
		44 => "0000000010110",
		45 => "0000000011010",
		46 => "0000000010111",
		47 => "0000000101110",
		48 => "0000011110111",
		49 => "0000101010011",
		50 => "0000101000111",
		51 => "0000010000001",
		52 => "0000000001110",
		53 => "0000001000000",
		54 => "0000100001111",
		55 => "0000010010011",
		56 => "0000011110010",
		57 => "0000001010101",
		58 => "0000010100000",
		59 => "0000001111101",
		60 => "0000000100111",
		61 => "0000011011010",
		62 => "0000100100111",
		63 => "0000010010111",
		64 => "0000010101101",
		65 => "0000001100110",
		66 => "0000010001110",
		67 => "0000010111110",
		68 => "0000010001111",
		69 => "0000010101110",
		70 => "0000010011011",
		71 => "0000001100111",
		72 => "0000010100101",
		73 => "0000100111111",
		74 => "0000011101001",
		75 => "0000010110001",
		76 => "0000000000100",
		77 => "0000011001101",
		78 => "0000000101010",
		79 => "0000100111010",
		80 => "0000000011100",
		81 => "0000001010110",
		82 => "0000000100010",
		83 => "0000001010000",
		84 => "0000000011110",
		85 => "0000011001000",
		86 => "0000011100101",
		87 => "0000000010010",
		88 => "0000000001001",
		89 => "0000100011101",
		90 => "0000010111111",
		91 => "0000000110110",
		92 => "0000010110000",
		93 => "0000000111110",
		94 => "0000100101100",
		95 => "0000010001010",
		96 => "0000000010001",
		97 => "0000010010001",
		98 => "0000010001101",
		99 => "0000100000010",
		100 => "0000010000011",
		101 => "0000001101100",
		102 => "0000011011111",
		103 => "0000010111011",
		104 => "0000011111111",
		105 => "0000011000010",
		106 => "0000010010010",
		107 => "0000000001010",
		108 => "0000000011001",
		109 => "0000010100010",
		110 => "0000011100111",
		111 => "0000011111010",
		112 => "0000000100110",
		113 => "0000011100100",
		114 => "0000000011000",
		115 => "0000010111010",
		116 => "0000000100101",
		117 => "0000101001100",
		118 => "0000100100101",
		119 => "0000001101011",
		120 => "0000010101100",
		121 => "0000000001011",
		122 => "0000001001001",
		123 => "0000011110000",
		124 => "0000000010100",
		125 => "0000010000101",
		126 => "0000001111010",
		127 => "0000001111111",
		128 => "0000000110011",
		129 => "0000010011000",
		130 => "0000101011000",
		131 => "0000001100101",
		132 => "0000011101011",
		133 => "0000000101000",
		134 => "0000010100100",
		135 => "0000010001001",
		136 => "0000100001010",
		137 => "0000000011101",
		138 => "0000000011011",
		139 => "0000011001100",
		140 => "0000010010110",
		141 => "0000000101101",
		142 => "0000001101111",
		143 => "0000000110100",
		144 => "0000000001100",
		145 => "0000000000101",
		146 => "0000101000001",
		147 => "0000001001110",
		148 => "0000000101011",
		149 => "0000100010001",
		150 => "0000100000011",
		151 => "0000100000110",
		152 => "0000010010101",
		153 => "0000101001001",
		154 => "0000100110001",
		155 => "0000001011100",
		156 => "0000010000010",
		157 => "0000001000001",
		158 => "0000100110101",
		159 => "0000001010010",
		160 => "0000000010101",
		161 => "0000100001100",
		162 => "0000011010011",
		163 => "0000010101001",
		164 => "0000010110110",
		165 => "0000100100010",
		166 => "0000001011101",
		167 => "0000101000110",
		168 => "0000000110101",
		169 => "0000011001010",
		170 => "0000010011111",
		171 => "0000001011110",
		172 => "0000100110111",
		173 => "0000100011001",
		174 => "0000011001001",
		175 => "0000011010110",
		176 => "0000000011111",
		177 => "0000010110101",
		178 => "0000011101101",
		179 => "0000000110111",
		180 => "0000010000100",
		181 => "0000000010011",
		182 => "0000100101000",
		183 => "0000001011111",
		184 => "0000011000100",
		185 => "0000011001111",
		186 => "0000011010000",
		187 => "0000000110010",
		188 => "0000010011110",
		189 => "0000100011011",
		190 => "0000010110100",
		191 => "0000001000011",
		192 => "0000000101001",
		193 => "0000011111101",
		194 => "0000011000110",
		195 => "0000000111111",
		196 => "0000010101111",
		197 => "0000001110001",
		198 => "0000000001000",
		199 => "0000010111100",
		200 => "0000000111001",
		201 => "0000000111010",
		202 => "0000001000101",
		203 => "0000001101110",
		204 => "0000000111011",
		205 => "0000000010000",
		206 => "0000000100000",
		207 => "0000000101100",
		208 => "0000011000111",
		209 => "0000100011111",
		210 => "0000010111101",
		211 => "0000010101011",
		212 => "0000100101101",
		213 => "0000011001011",
		214 => "0000010001011",
		215 => "0000101001111",
		216 => "0000001011000",
		217 => "0000100101011",
		218 => "0000000100100",
		219 => "0000100110010",
		220 => "0000001010001",
		221 => "0000001101001",
		222 => "0000010110111",
		223 => "0000010100111",
		224 => "0000000011010",
		225 => "0000001000100",
		226 => "0000010011001",
		227 => "0000000100010",
		228 => "0000100011110",
		229 => "0000011011011",
		230 => "0000000111101",
		231 => "0000010001000",
		232 => "0000101000011",
		233 => "0000000011111",
		234 => "0000100111100",
		235 => "0000001111011",
		236 => "0000010101000",
		237 => "0000001110010",
		238 => "0000100000111",
		239 => "0000001100000",
		240 => "0000001110000",
		241 => "0000010111001",
		242 => "0000000111100",
		243 => "0000011000011",
		244 => "0000010000110",
		245 => "0000000100011",
		246 => "0000000001111",
		247 => "0000001010100",
		248 => "0000001011010",
		249 => "0000000110001",
		250 => "0000100110000",
		251 => "0000100100001",
		252 => "0000001000111",
		253 => "0000001100001",
		254 => "0000001100011",
		255 => "0000011011101",
		others => (others => '0')
	);

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
