-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive;
            DATA_LENGTH:  positive;
            SELECT_ROM:  integer := 0); -- Select which ROM to use
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0);
         initial_addr_2: out std_logic_vector (ADDRESS_BITS - 1 downto 0);
         initial_addr_3: out std_logic_vector (ADDRESS_BITS - 1 downto 0));
end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin

	gen_rom_0: if SELECT_ROM = 0 generate
		bank <= (
			0 => "0011010111011100001100",
			1 => "0010001111001000000100",
			2 => "1111111000000001011101",
			3 => "0001010101111000000100",
			4 => "0000001000000001011101",
			5 => "1111111000000001011101",
			6 => "0011111010011000000100",
			7 => "1111111000000001011101",
			8 => "0001010101110000011100",
			9 => "0001111100011100010000",
			10 => "0000000100110100000100",
			11 => "0000001000000001011101",
			12 => "0010011010000100000100",
			13 => "1111111000000001011101",
			14 => "0000101111001100000100",
			15 => "0000000000000001011101",
			16 => "0000000000000001011101",
			17 => "0001011011000000001000",
			18 => "0010101111101000000100",
			19 => "0000001000000001011101",
			20 => "0000000000000001011101",
			21 => "0000001000000001011101",
			22 => "1111111000000001011101",
			23 => "0011010111011100010000",
			24 => "0001010101111000001000",
			25 => "0010101000000000000100",
			26 => "0000000000000011101001",
			27 => "0000000000000011101001",
			28 => "0010011111011000000100",
			29 => "0000000000000011101001",
			30 => "0000000000000011101001",
			31 => "0001000110101100011100",
			32 => "0011111010011000000100",
			33 => "0000000000000011101001",
			34 => "0000001010111000010000",
			35 => "0010010110000000000100",
			36 => "0000000000000011101001",
			37 => "0010101111101000000100",
			38 => "0000000000000011101001",
			39 => "0010001111011000000100",
			40 => "0000000000000011101001",
			41 => "0000000000000011101001",
			42 => "0011011101101000000100",
			43 => "0000000000000011101001",
			44 => "0000000000000011101001",
			45 => "0001001001010000001100",
			46 => "0000010101011100001000",
			47 => "0000000110111100000100",
			48 => "0000000000000011101001",
			49 => "0000000000000011101001",
			50 => "0000000000000011101001",
			51 => "0000110011110100001000",
			52 => "0000001110110100000100",
			53 => "0000000000000011101001",
			54 => "0000000000000011101001",
			55 => "0000010111011100000100",
			56 => "0000000000000011101001",
			57 => "0000000000000011101001",
			58 => "0000010110001100100000",
			59 => "0010000000110000010000",
			60 => "0000010011110000000100",
			61 => "1111111000000101110101",
			62 => "0010111010100100001000",
			63 => "0011011010100100000100",
			64 => "1111111000000101110101",
			65 => "0000000000000101110101",
			66 => "1111111000000101110101",
			67 => "0011001001001000001000",
			68 => "0010011010000100000100",
			69 => "0000000000000101110101",
			70 => "0000010000000101110101",
			71 => "0011001001000100000100",
			72 => "0000000000000101110101",
			73 => "1111111000000101110101",
			74 => "0011111101100000001000",
			75 => "0010010011001000000100",
			76 => "0000000000000101110101",
			77 => "1111111000000101110101",
			78 => "0000111010011100011100",
			79 => "0011010101011100000100",
			80 => "0000000000000101110101",
			81 => "0001011000100000010000",
			82 => "0001110011110100001000",
			83 => "0000101111001100000100",
			84 => "0000001000000101110101",
			85 => "1111111000000101110101",
			86 => "0001001000000000000100",
			87 => "0000001000000101110101",
			88 => "0000001000000101110101",
			89 => "0011000101101100000100",
			90 => "0000001000000101110101",
			91 => "0000001000000101110101",
			92 => "1111111000000101110101",
			93 => "0000011110011000111000",
			94 => "0000010110001100100100",
			95 => "0000010011110000001000",
			96 => "0010001111011000000100",
			97 => "1111111000001000011001",
			98 => "1111111000001000011001",
			99 => "0011110100010000001100",
			100 => "0011000101011100001000",
			101 => "0001110011001000000100",
			102 => "1111111000001000011001",
			103 => "0000000000001000011001",
			104 => "1111111000001000011001",
			105 => "0010000000110000001000",
			106 => "0010101001010100000100",
			107 => "0000000000001000011001",
			108 => "1111111000001000011001",
			109 => "0011110110011000000100",
			110 => "0000010000001000011001",
			111 => "0000000000001000011001",
			112 => "0011111101100000001000",
			113 => "0001101010011000000100",
			114 => "1111111000001000011001",
			115 => "0000000000001000011001",
			116 => "0000000110101000000100",
			117 => "0000010000001000011001",
			118 => "0001010011000100000100",
			119 => "1111111000001000011001",
			120 => "0000001000001000011001",
			121 => "0011110011101000001000",
			122 => "0011000011001000000100",
			123 => "0000000000001000011001",
			124 => "1111111000001000011001",
			125 => "0010010011001000000100",
			126 => "0000000000001000011001",
			127 => "0010000011100100000100",
			128 => "0000001000001000011001",
			129 => "0011010101101100000100",
			130 => "0000010000001000011001",
			131 => "0001000011000000000100",
			132 => "0000001000001000011001",
			133 => "0000010000001000011001",
			134 => "0011010101011100010100",
			135 => "0001010101111000001000",
			136 => "0010101000000000000100",
			137 => "0000000000001011001101",
			138 => "0000000000001011001101",
			139 => "0011100101001100001000",
			140 => "0010101000000000000100",
			141 => "0000000000001011001101",
			142 => "0000000000001011001101",
			143 => "0000000000001011001101",
			144 => "0011000110000000011100",
			145 => "0011100100010000010000",
			146 => "0001101110010000001000",
			147 => "0001101010001100000100",
			148 => "0000000000001011001101",
			149 => "0000000000001011001101",
			150 => "0011110010111100000100",
			151 => "0000000000001011001101",
			152 => "0000000000001011001101",
			153 => "0000100101101000000100",
			154 => "0000000000001011001101",
			155 => "0011100001100000000100",
			156 => "0000000000001011001101",
			157 => "0000000000001011001101",
			158 => "0000010111011100011000",
			159 => "0001010011000100001100",
			160 => "0001011011111000001000",
			161 => "0000011110011000000100",
			162 => "0000000000001011001101",
			163 => "0000000000001011001101",
			164 => "0000000000001011001101",
			165 => "0001011010100000001000",
			166 => "0011110111000000000100",
			167 => "0000000000001011001101",
			168 => "0000000000001011001101",
			169 => "0000000000001011001101",
			170 => "0011101010001000001100",
			171 => "0000001010010100001000",
			172 => "0001100110110000000100",
			173 => "0000000000001011001101",
			174 => "0000000000001011001101",
			175 => "0000000000001011001101",
			176 => "0010111101101000000100",
			177 => "0000000000001011001101",
			178 => "0000000000001011001101",
			179 => "0000011110011000110100",
			180 => "0000010110001100100100",
			181 => "0000011101000000011000",
			182 => "0010001111011000010000",
			183 => "0000010011110000000100",
			184 => "1110000000001101111001",
			185 => "0011110100010000000100",
			186 => "1110000000001101111001",
			187 => "0001101010111100000100",
			188 => "1110001000001101111001",
			189 => "1110000000001101111001",
			190 => "0010011100000000000100",
			191 => "1110001000001101111001",
			192 => "1110000000001101111001",
			193 => "0011111101100000000100",
			194 => "1110000000001101111001",
			195 => "0000000000000000000100",
			196 => "1110010000001101111001",
			197 => "1110000000001101111001",
			198 => "0011111101100000001000",
			199 => "0010011100000000000100",
			200 => "1110000000001101111001",
			201 => "1110000000001101111001",
			202 => "0001010011000100000100",
			203 => "1110001000001101111001",
			204 => "1110100000001101111001",
			205 => "0001101100011000001000",
			206 => "0001110001010000000100",
			207 => "1110000000001101111001",
			208 => "1110000000001101111001",
			209 => "0001000011000000001000",
			210 => "0010111001000100000100",
			211 => "1110010000001101111001",
			212 => "1110101000001101111001",
			213 => "0010000011100100000100",
			214 => "1110100000001101111001",
			215 => "0000010111011100001100",
			216 => "0001010011000100000100",
			217 => "1110100000001101111001",
			218 => "0001011010011100000100",
			219 => "1110110000001101111001",
			220 => "1110101000001101111001",
			221 => "1110110000001101111001",
			222 => "0000010110001100100000",
			223 => "0010000000110000010000",
			224 => "0000010011110000000100",
			225 => "1111111000010000000101",
			226 => "0000100101011000001000",
			227 => "0001101001011100000100",
			228 => "1111111000010000000101",
			229 => "0000001000010000000101",
			230 => "1111111000010000000101",
			231 => "0011001001000100001100",
			232 => "0010011010000100000100",
			233 => "0000000000010000000101",
			234 => "0001011100101100000100",
			235 => "0000000000010000000101",
			236 => "0000001000010000000101",
			237 => "1111111000010000000101",
			238 => "0001101010001100000100",
			239 => "1111111000010000000101",
			240 => "0000110000111000100000",
			241 => "0011011101101000010100",
			242 => "0011111100111000000100",
			243 => "0000001000010000000101",
			244 => "0001000011000000001000",
			245 => "0001001010000100000100",
			246 => "0000000000010000000101",
			247 => "1111111000010000000101",
			248 => "0001111001011000000100",
			249 => "0000000000010000000101",
			250 => "0000001000010000000101",
			251 => "0000111001010000001000",
			252 => "0000111001010100000100",
			253 => "0000001000010000000101",
			254 => "0000000000010000000101",
			255 => "0000001000010000000101",
			256 => "1111111000010000000101",
			257 => "0010001111011000100000",
			258 => "0011110111010000011000",
			259 => "0000010011110000000100",
			260 => "0000000000010011000001",
			261 => "0011111101100000001100",
			262 => "0010101100010000001000",
			263 => "0000010110001100000100",
			264 => "0000000000010011000001",
			265 => "0000000000010011000001",
			266 => "0000000000010011000001",
			267 => "0011111010101100000100",
			268 => "0000000000010011000001",
			269 => "0000000000010011000001",
			270 => "0011100101001100000100",
			271 => "0000000000010011000001",
			272 => "0000000000010011000001",
			273 => "0000100000101000100100",
			274 => "0000011100101000011000",
			275 => "0001111011111000001100",
			276 => "0000001110011100001000",
			277 => "0000000111101000000100",
			278 => "0000000000010011000001",
			279 => "0000000000010011000001",
			280 => "0000000000010011000001",
			281 => "0000110000111000001000",
			282 => "0001101100011000000100",
			283 => "0000000000010011000001",
			284 => "0000001000010011000001",
			285 => "0000000000010011000001",
			286 => "0011110110011000001000",
			287 => "0000001010101000000100",
			288 => "0000000000010011000001",
			289 => "0000000000010011000001",
			290 => "0000000000010011000001",
			291 => "0000010101011100010000",
			292 => "0011000101101100000100",
			293 => "0000000000010011000001",
			294 => "0001010011000100000100",
			295 => "0000000000010011000001",
			296 => "0001101110000100000100",
			297 => "0000000000010011000001",
			298 => "0000000000010011000001",
			299 => "0000011100101000000100",
			300 => "0000000000010011000001",
			301 => "0000010101101100000100",
			302 => "0000000000010011000001",
			303 => "0000000000010011000001",
			304 => "0000010110001100100000",
			305 => "0010000000110000010000",
			306 => "0000010011110000000100",
			307 => "1111111000010101010101",
			308 => "0010110111011100001000",
			309 => "0010011001000100000100",
			310 => "1111111000010101010101",
			311 => "0000001000010101010101",
			312 => "1111111000010101010101",
			313 => "0011001001000100001100",
			314 => "0001111101001000000100",
			315 => "1111111000010101010101",
			316 => "0011110110011000000100",
			317 => "0000010000010101010101",
			318 => "0000000000010101010101",
			319 => "1111111000010101010101",
			320 => "0011111111010100001000",
			321 => "0010110101101100000100",
			322 => "0000000000010101010101",
			323 => "1111111000010101010101",
			324 => "0011010101011100000100",
			325 => "0000000000010101010101",
			326 => "0010100000111000011100",
			327 => "0001010011000100001100",
			328 => "0000000110101000000100",
			329 => "0000010000010101010101",
			330 => "0001110011110100000100",
			331 => "0000000000010101010101",
			332 => "0000001000010101010101",
			333 => "0001110000111100001000",
			334 => "0011101101100100000100",
			335 => "0000001000010101010101",
			336 => "0000001000010101010101",
			337 => "0011000110000000000100",
			338 => "0000001000010101010101",
			339 => "0000001000010101010101",
			340 => "0000000000010101010101",
			341 => "0010001111011000100000",
			342 => "0001101010001000011000",
			343 => "0001100010110000010000",
			344 => "0011010101010100000100",
			345 => "0000000000011000000001",
			346 => "0010101111101000001000",
			347 => "0010101000111000000100",
			348 => "0000000000011000000001",
			349 => "0000000000011000000001",
			350 => "0000000000011000000001",
			351 => "0000011001100000000100",
			352 => "0000000000011000000001",
			353 => "0000000000011000000001",
			354 => "0001001100110000000100",
			355 => "0000000000011000000001",
			356 => "0000000000011000000001",
			357 => "0010101100001100101100",
			358 => "0001010011000100100000",
			359 => "0001110011110100011000",
			360 => "0001001010000100001100",
			361 => "0010011000000100000100",
			362 => "0000000000011000000001",
			363 => "0011011101101000000100",
			364 => "0000000000011000000001",
			365 => "0000000000011000000001",
			366 => "0000011110011000000100",
			367 => "0000000000011000000001",
			368 => "0011110110011000000100",
			369 => "0000000000011000000001",
			370 => "0000000000011000000001",
			371 => "0011010011001000000100",
			372 => "0000000000011000000001",
			373 => "0000000000011000000001",
			374 => "0011110000000100001000",
			375 => "0000111011111000000100",
			376 => "0000000000011000000001",
			377 => "0000000000011000000001",
			378 => "0000000000011000000001",
			379 => "0000010101010100001000",
			380 => "0001111010011100000100",
			381 => "0000000000011000000001",
			382 => "0000000000011000000001",
			383 => "0000000000011000000001",
			384 => "0001011100101100100000",
			385 => "0010001000000000011000",
			386 => "0000100000100100001100",
			387 => "0011100010011100000100",
			388 => "0000000000011010111101",
			389 => "0011011010100100000100",
			390 => "0000000000011010111101",
			391 => "0000000000011010111101",
			392 => "0010101000000000001000",
			393 => "0001111101001000000100",
			394 => "0000000000011010111101",
			395 => "0000000000011010111101",
			396 => "0000000000011010111101",
			397 => "0011100110110000000100",
			398 => "0000000000011010111101",
			399 => "0000000000011010111101",
			400 => "0010100000111100100100",
			401 => "0000101111001100011000",
			402 => "0000010011110000000100",
			403 => "0000000000011010111101",
			404 => "0000011100101000001100",
			405 => "0001100010111100001000",
			406 => "0001001001010100000100",
			407 => "0000000000011010111101",
			408 => "0000000000011010111101",
			409 => "0000000000011010111101",
			410 => "0000111111101000000100",
			411 => "0000000000011010111101",
			412 => "0000000000011010111101",
			413 => "0000101001101000001000",
			414 => "0001100000001000000100",
			415 => "0000000000011010111101",
			416 => "0000000000011010111101",
			417 => "0000000000011010111101",
			418 => "0001101110000100011000",
			419 => "0000010111011100010000",
			420 => "0001111011111000001000",
			421 => "0001111111101000000100",
			422 => "0000000000011010111101",
			423 => "0000000000011010111101",
			424 => "0001110011110100000100",
			425 => "0000000000011010111101",
			426 => "0000000000011010111101",
			427 => "0000001111101100000100",
			428 => "0000000000011010111101",
			429 => "0000000000011010111101",
			430 => "0000000000011010111101",
			431 => "0000010110001100011100",
			432 => "0010001111011000010100",
			433 => "0000010011110000000100",
			434 => "1111111000011101011001",
			435 => "0011111101100000000100",
			436 => "1111111000011101011001",
			437 => "0011100001101100000100",
			438 => "0000001000011101011001",
			439 => "0001111011000000000100",
			440 => "1111111000011101011001",
			441 => "0000000000011101011001",
			442 => "0011001001000100000100",
			443 => "0000001000011101011001",
			444 => "1111111000011101011001",
			445 => "0011111101100000001000",
			446 => "0010011111011000000100",
			447 => "0000000000011101011001",
			448 => "1111111000011101011001",
			449 => "0001111100011100011000",
			450 => "0000101111001100010100",
			451 => "0011010101011100000100",
			452 => "0000000000011101011001",
			453 => "0000000110101000001000",
			454 => "0001110011000100000100",
			455 => "0000001000011101011001",
			456 => "0000001000011101011001",
			457 => "0000011110011000000100",
			458 => "0000000000011101011001",
			459 => "0000001000011101011001",
			460 => "1111111000011101011001",
			461 => "0000000011001100000100",
			462 => "0000001000011101011001",
			463 => "0001011011000000001000",
			464 => "0000101011001100000100",
			465 => "0000001000011101011001",
			466 => "0000001000011101011001",
			467 => "0010001000000000000100",
			468 => "0000001000011101011001",
			469 => "0000001000011101011001",
			470 => "0010001111011000011100",
			471 => "0000010011110000000100",
			472 => "1111111000011111011101",
			473 => "0010011001000100000100",
			474 => "1111111000011111011101",
			475 => "0011001100101000001100",
			476 => "0010101001010100000100",
			477 => "0000001000011111011101",
			478 => "0001110001010000000100",
			479 => "1111111000011111011101",
			480 => "0000000000011111011101",
			481 => "0011110011101000000100",
			482 => "1111111000011111011101",
			483 => "0000000000011111011101",
			484 => "0011110000110100000100",
			485 => "1111111000011111011101",
			486 => "0000110000111000100000",
			487 => "0001010011000100010000",
			488 => "0000111000000000000100",
			489 => "0000001000011111011101",
			490 => "0001111110001100001000",
			491 => "0000100100010100000100",
			492 => "0000000000011111011101",
			493 => "0000000000011111011101",
			494 => "0000001000011111011101",
			495 => "0001110000111100001000",
			496 => "0010011100000000000100",
			497 => "0000000000011111011101",
			498 => "0000001000011111011101",
			499 => "0011000110000000000100",
			500 => "0000001000011111011101",
			501 => "0000001000011111011101",
			502 => "1111111000011111011101",
			503 => "0011100010110101001100",
			504 => "0011111100111100110100",
			505 => "0001000101111000011000",
			506 => "0010010110000000001100",
			507 => "0001001010000100000100",
			508 => "0000000000100010100001",
			509 => "0000001011110100000100",
			510 => "0000000000100010100001",
			511 => "0000000000100010100001",
			512 => "0001101010011000000100",
			513 => "0000000000100010100001",
			514 => "0010101111101000000100",
			515 => "0000000000100010100001",
			516 => "0000000000100010100001",
			517 => "0010000011001000010000",
			518 => "0011110010111100001100",
			519 => "0011011001001000000100",
			520 => "0000000000100010100001",
			521 => "0011010101101100000100",
			522 => "0000000000100010100001",
			523 => "0000000000100010100001",
			524 => "0000000000100010100001",
			525 => "0000110000111000001000",
			526 => "0011101100011000000100",
			527 => "0000000000100010100001",
			528 => "0000000000100010100001",
			529 => "0000000000100010100001",
			530 => "0010001000111000010100",
			531 => "0001001001000100001000",
			532 => "0010101101001000000100",
			533 => "0000000000100010100001",
			534 => "0000000000100010100001",
			535 => "0010110101010100001000",
			536 => "0010110111011100000100",
			537 => "0000000000100010100001",
			538 => "0000000000100010100001",
			539 => "0000000000100010100001",
			540 => "0000000000100010100001",
			541 => "0000010111011100010000",
			542 => "0001010011000100001000",
			543 => "0001101110000100000100",
			544 => "0000000000100010100001",
			545 => "0000000000100010100001",
			546 => "0001101110000100000100",
			547 => "0000000000100010100001",
			548 => "0000000000100010100001",
			549 => "0011011101101000000100",
			550 => "0000000000100010100001",
			551 => "0000000000100010100001",
			552 => "0011010111011100001100",
			553 => "0010011111011000000100",
			554 => "1111111000100101000101",
			555 => "0010001001000100000100",
			556 => "0000000000100101000101",
			557 => "0000000000100101000101",
			558 => "0001111110111000111000",
			559 => "0011110110011000100100",
			560 => "0010000011100100011000",
			561 => "0011000101011100001000",
			562 => "0010010110000000000100",
			563 => "1111111000100101000101",
			564 => "0000000000100101000101",
			565 => "0001110001001000001000",
			566 => "0010011111011000000100",
			567 => "1111111000100101000101",
			568 => "0000000000100101000101",
			569 => "0000011101000000000100",
			570 => "0000000000100101000101",
			571 => "0000001000100101000101",
			572 => "0010011101001000001000",
			573 => "0000001010101000000100",
			574 => "0000000000100101000101",
			575 => "0000001000100101000101",
			576 => "1111111000100101000101",
			577 => "0001000011000000001000",
			578 => "0011110100110100000100",
			579 => "1111111000100101000101",
			580 => "0000000000100101000101",
			581 => "0001101101010000000100",
			582 => "0000001000100101000101",
			583 => "0010000011100100000100",
			584 => "1111111000100101000101",
			585 => "0000000000100101000101",
			586 => "0000111001010000001000",
			587 => "0000111001010100000100",
			588 => "0000001000100101000101",
			589 => "1111111000100101000101",
			590 => "0000111010100000000100",
			591 => "0000001000100101000101",
			592 => "0000000000100101000101",
			593 => "0010000011100101000000",
			594 => "0000100110010100101000",
			595 => "0010110110000000100100",
			596 => "0010010110000000001100",
			597 => "0001010101111000001000",
			598 => "0010101000000000000100",
			599 => "0000000000101000010001",
			600 => "0000000000101000010001",
			601 => "0000000000101000010001",
			602 => "0011010111011100001100",
			603 => "0001010011001000000100",
			604 => "0000000000101000010001",
			605 => "0010011111011000000100",
			606 => "0000000000101000010001",
			607 => "0000000000101000010001",
			608 => "0011111010011000000100",
			609 => "0000000000101000010001",
			610 => "0001001100101100000100",
			611 => "0000000000101000010001",
			612 => "0000000000101000010001",
			613 => "0000000000101000010001",
			614 => "0001010001001000010000",
			615 => "0011100101100000001100",
			616 => "0010101111101000001000",
			617 => "0010101000101000000100",
			618 => "0000000000101000010001",
			619 => "0000000000101000010001",
			620 => "0000000000101000010001",
			621 => "0000000000101000010001",
			622 => "0001101010101100000100",
			623 => "0000000000101000010001",
			624 => "0000000000101000010001",
			625 => "0001000011000000010000",
			626 => "0000111000000000001100",
			627 => "0010001000000000000100",
			628 => "0000000000101000010001",
			629 => "0010111000000100000100",
			630 => "0000000000101000010001",
			631 => "0000000000101000010001",
			632 => "0000000000101000010001",
			633 => "0000011110011000001000",
			634 => "0000100011100000000100",
			635 => "0000000000101000010001",
			636 => "0000000000101000010001",
			637 => "0010001001010100001000",
			638 => "0000111110001100000100",
			639 => "0000000000101000010001",
			640 => "0000000000101000010001",
			641 => "0011101010001000000100",
			642 => "0000000000101000010001",
			643 => "0000000000101000010001",
			644 => "0010001111011000100000",
			645 => "0011110111010000011000",
			646 => "0000010011110000000100",
			647 => "0000000000101011011101",
			648 => "0011111101100000001100",
			649 => "0010101100010000001000",
			650 => "0000010110001100000100",
			651 => "0000000000101011011101",
			652 => "0000000000101011011101",
			653 => "0000000000101011011101",
			654 => "0011111010101100000100",
			655 => "0000000000101011011101",
			656 => "0000000000101011011101",
			657 => "0011100101001100000100",
			658 => "0000000000101011011101",
			659 => "0000000000101011011101",
			660 => "0000100000101000110000",
			661 => "0000011100101000100100",
			662 => "0001100001100000011000",
			663 => "0000111001010100001000",
			664 => "0000000000001100000100",
			665 => "0000000000101011011101",
			666 => "0000000000101011011101",
			667 => "0000011110011000001000",
			668 => "0000001000100100000100",
			669 => "0000000000101011011101",
			670 => "0000000000101011011101",
			671 => "0001011100001100000100",
			672 => "0000000000101011011101",
			673 => "0000000000101011011101",
			674 => "0001001011111000001000",
			675 => "0000100100010100000100",
			676 => "0000001000101011011101",
			677 => "0000000000101011011101",
			678 => "0000000000101011011101",
			679 => "0011110110011000001000",
			680 => "0000001010101000000100",
			681 => "0000000000101011011101",
			682 => "0000000000101011011101",
			683 => "0000000000101011011101",
			684 => "0001110011110100001100",
			685 => "0000111001010000000100",
			686 => "0000000000101011011101",
			687 => "0000111111101000000100",
			688 => "0000000000101011011101",
			689 => "0000000000101011011101",
			690 => "0011000011000000000100",
			691 => "0000000000101011011101",
			692 => "0011001111011000000100",
			693 => "0000000000101011011101",
			694 => "0000000000101011011101",
			695 => "0000010110001100100000",
			696 => "0010000000110000010000",
			697 => "0000010011110000000100",
			698 => "1111111000101101111001",
			699 => "0001000110000000000100",
			700 => "1111111000101101111001",
			701 => "0000111100110000000100",
			702 => "0000001000101101111001",
			703 => "1111111000101101111001",
			704 => "0011001001000100001100",
			705 => "0001111101001000000100",
			706 => "1111111000101101111001",
			707 => "0011110100011000000100",
			708 => "0000001000101101111001",
			709 => "0000000000101101111001",
			710 => "1111111000101101111001",
			711 => "0011111010011000000100",
			712 => "1111111000101101111001",
			713 => "0010101110010100101000",
			714 => "0011011101101000010100",
			715 => "0011111100111000000100",
			716 => "0000001000101101111001",
			717 => "0001111001011000001000",
			718 => "0011110000001000000100",
			719 => "0000000000101101111001",
			720 => "1111111000101101111001",
			721 => "0000111100110000000100",
			722 => "0000000000101101111001",
			723 => "0000001000101101111001",
			724 => "0000010111011100001000",
			725 => "0001011000100000000100",
			726 => "0000000000101101111001",
			727 => "0000001000101101111001",
			728 => "0000111001010000001000",
			729 => "0011100001100000000100",
			730 => "0000001000101101111001",
			731 => "0000001000101101111001",
			732 => "0000001000101101111001",
			733 => "1111111000101101111001",
			734 => "0010001111011000110000",
			735 => "0011101110100000101000",
			736 => "0001111000101000011000",
			737 => "0010101100010000010100",
			738 => "0001001010000100001100",
			739 => "0011000111011100000100",
			740 => "0000000000110001001101",
			741 => "0011000101011100000100",
			742 => "0000000000110001001101",
			743 => "0000000000110001001101",
			744 => "0001011001010100000100",
			745 => "0000000000110001001101",
			746 => "0000000000110001001101",
			747 => "0000000000110001001101",
			748 => "0001000110011100001100",
			749 => "0000001000010000001000",
			750 => "0000010011110000000100",
			751 => "0000000000110001001101",
			752 => "0000000000110001001101",
			753 => "0000000000110001001101",
			754 => "0000000000110001001101",
			755 => "0011100101001100000100",
			756 => "1111111000110001001101",
			757 => "0000000000110001001101",
			758 => "0010100000111100100100",
			759 => "0000001010111000011000",
			760 => "0011100110110000001100",
			761 => "0011110100001000001000",
			762 => "0011111010011000000100",
			763 => "0000000000110001001101",
			764 => "0000000000110001001101",
			765 => "0000000000110001001101",
			766 => "0011000110000000000100",
			767 => "0000001000110001001101",
			768 => "0010001000111000000100",
			769 => "0000000000110001001101",
			770 => "0000000000110001001101",
			771 => "0011011101101000000100",
			772 => "0000000000110001001101",
			773 => "0001001000000000000100",
			774 => "0000000000110001001101",
			775 => "0000000000110001001101",
			776 => "0001101110000100010100",
			777 => "0000010111011100001100",
			778 => "0000000110111100001000",
			779 => "0000001101110100000100",
			780 => "0000000000110001001101",
			781 => "0000000000110001001101",
			782 => "0000000000110001001101",
			783 => "0000000010100100000100",
			784 => "0000000000110001001101",
			785 => "0000000000110001001101",
			786 => "0000000000110001001101",
			787 => "0010100000111100111100",
			788 => "0001011000100000110000",
			789 => "0011010011000000101000",
			790 => "0000101111001100011100",
			791 => "0000111000101000010000",
			792 => "0000111100110000001000",
			793 => "0000010011010000000100",
			794 => "0000000000110011110001",
			795 => "0000000000110011110001",
			796 => "0010010011000000000100",
			797 => "0000000000110011110001",
			798 => "0000000000110011110001",
			799 => "0000010111011100001000",
			800 => "0000111011111000000100",
			801 => "0000000000110011110001",
			802 => "0000000000110011110001",
			803 => "0000000000110011110001",
			804 => "0011110000011100000100",
			805 => "0000000000110011110001",
			806 => "0011110111101100000100",
			807 => "0000000000110011110001",
			808 => "0000000000110011110001",
			809 => "0000000010101100000100",
			810 => "0000000000110011110001",
			811 => "0000000000110011110001",
			812 => "0011010111011100000100",
			813 => "0000000000110011110001",
			814 => "0010111111011000000100",
			815 => "0000000000110011110001",
			816 => "0000000000110011110001",
			817 => "0001101110000100010100",
			818 => "0000000101101000010000",
			819 => "0011011001001000000100",
			820 => "0000000000110011110001",
			821 => "0001001110111000001000",
			822 => "0000000011111000000100",
			823 => "0000000000110011110001",
			824 => "0000000000110011110001",
			825 => "0000000000110011110001",
			826 => "0000000000110011110001",
			827 => "0000000000110011110001",
			828 => "0011011001001000110100",
			829 => "0011001100101000100100",
			830 => "0010010011000000011100",
			831 => "0000100000100100010100",
			832 => "0001000011000000001100",
			833 => "0010011001000100000100",
			834 => "0000000000110111010101",
			835 => "0000000110000100000100",
			836 => "0000000000110111010101",
			837 => "0000000000110111010101",
			838 => "0000000000100100000100",
			839 => "0000000000110111010101",
			840 => "0000000000110111010101",
			841 => "0001010001001000000100",
			842 => "0000000000110111010101",
			843 => "0000000000110111010101",
			844 => "0001101101000100000100",
			845 => "0000000000110111010101",
			846 => "0000000000110111010101",
			847 => "0001010001001000000100",
			848 => "0000000000110111010101",
			849 => "0010100000111100000100",
			850 => "0000000000110111010101",
			851 => "0001111000100000000100",
			852 => "0000000000110111010101",
			853 => "0000000000110111010101",
			854 => "0001000011000000011100",
			855 => "0010000011001000001000",
			856 => "0001110100101100000100",
			857 => "0000000000110111010101",
			858 => "0000000000110111010101",
			859 => "0010001100110000010000",
			860 => "0001001100101000001000",
			861 => "0001000101010100000100",
			862 => "0000000000110111010101",
			863 => "0000000000110111010101",
			864 => "0011101111010100000100",
			865 => "0000000000110111010101",
			866 => "0000000000110111010101",
			867 => "0000000000110111010101",
			868 => "0010101100001100011100",
			869 => "0011011010000100001100",
			870 => "0000001000001100001000",
			871 => "0011100010110000000100",
			872 => "0000000000110111010101",
			873 => "0000000000110111010101",
			874 => "0000000000110111010101",
			875 => "0010010110101100001000",
			876 => "0001010011000100000100",
			877 => "0000000000110111010101",
			878 => "0000000000110111010101",
			879 => "0000001100100100000100",
			880 => "0000000000110111010101",
			881 => "0000000000110111010101",
			882 => "0000111100110100000100",
			883 => "0000000000110111010101",
			884 => "0000000000110111010101",
			885 => "0011010111011100001000",
			886 => "0010000000110000000100",
			887 => "1111111000111001001001",
			888 => "0000000000111001001001",
			889 => "0000111100110100110000",
			890 => "0001011000100000100000",
			891 => "0001001100010000011100",
			892 => "0011011101101000010000",
			893 => "0011110000001100001000",
			894 => "0001101010001100000100",
			895 => "1111111000111001001001",
			896 => "0000001000111001001001",
			897 => "0001111011111000000100",
			898 => "1111111000111001001001",
			899 => "0000000000111001001001",
			900 => "0011101010001000001000",
			901 => "0010001100110000000100",
			902 => "0000001000111001001001",
			903 => "0000000000111001001001",
			904 => "0000001000111001001001",
			905 => "1111111000111001001001",
			906 => "0010000000110000000100",
			907 => "1111111000111001001001",
			908 => "0010111001001000000100",
			909 => "0000000000111001001001",
			910 => "0000101010101000000100",
			911 => "0000000000111001001001",
			912 => "0000001000111001001001",
			913 => "1111111000111001001001",
			914 => "0011010111011100010100",
			915 => "0001010011001000001100",
			916 => "0010011001000100000100",
			917 => "0000000000111011110101",
			918 => "0010101000000100000100",
			919 => "0000000000111011110101",
			920 => "0000000000111011110101",
			921 => "0010011111011000000100",
			922 => "0000000000111011110101",
			923 => "0000000000111011110101",
			924 => "0000110011110100111100",
			925 => "0001011000100000101000",
			926 => "0001001000111000100000",
			927 => "0001000011000000010000",
			928 => "0011101111010100001000",
			929 => "0001011100010000000100",
			930 => "0000000000111011110101",
			931 => "0000000000111011110101",
			932 => "0001001010000100000100",
			933 => "0000000000111011110101",
			934 => "0000000000111011110101",
			935 => "0000011110011000001000",
			936 => "0011010101011100000100",
			937 => "0000000000111011110101",
			938 => "0000000000111011110101",
			939 => "0010000110101100000100",
			940 => "0000000000111011110101",
			941 => "0000000000111011110101",
			942 => "0000010111011100000100",
			943 => "0000000000111011110101",
			944 => "0000000000111011110101",
			945 => "0011110000000100001000",
			946 => "0010011000000100000100",
			947 => "0000000000111011110101",
			948 => "0000000000111011110101",
			949 => "0000110000111100001000",
			950 => "0000111000101000000100",
			951 => "0000000000111011110101",
			952 => "0000000000111011110101",
			953 => "0000000000111011110101",
			954 => "0001000110011100000100",
			955 => "0000000000111011110101",
			956 => "0000000000111011110101",
			957 => "0011010011000000110000",
			958 => "0010011001000100000100",
			959 => "1111111000111101100001",
			960 => "0011100101100000101000",
			961 => "0000101111001100011100",
			962 => "0011111101001100010000",
			963 => "0011000101010100001000",
			964 => "0001001101101000000100",
			965 => "0000000000111101100001",
			966 => "0000001000111101100001",
			967 => "0010000000110000000100",
			968 => "1111111000111101100001",
			969 => "0000000000111101100001",
			970 => "0000011110011000000100",
			971 => "0000000000111101100001",
			972 => "0011110000101100000100",
			973 => "0000001000111101100001",
			974 => "0000000000111101100001",
			975 => "0001011000100000001000",
			976 => "0001011000101000000100",
			977 => "0000000000111101100001",
			978 => "1111111000111101100001",
			979 => "0000000000111101100001",
			980 => "0000000000111101100001",
			981 => "0001101000101100000100",
			982 => "0000000000111101100001",
			983 => "0000001000111101100001",
			984 => "0011011101101001010000",
			985 => "0000100100010100101100",
			986 => "0011110000000100100000",
			987 => "0011111100111000011100",
			988 => "0011010101010100010000",
			989 => "0001010011001000001000",
			990 => "0000110011001000000100",
			991 => "0000000001000000111101",
			992 => "0000000001000000111101",
			993 => "0011100010001000000100",
			994 => "0000000001000000111101",
			995 => "0000000001000000111101",
			996 => "0011111010011000000100",
			997 => "0000000001000000111101",
			998 => "0011000110000000000100",
			999 => "0000000001000000111101",
			1000 => "0000000001000000111101",
			1001 => "0000000001000000111101",
			1002 => "0001011001010000000100",
			1003 => "0000000001000000111101",
			1004 => "0001001000000000000100",
			1005 => "0000000001000000111101",
			1006 => "0000000001000000111101",
			1007 => "0001001000000000011000",
			1008 => "0010101101001000001000",
			1009 => "0001011000111000000100",
			1010 => "0000000001000000111101",
			1011 => "0000000001000000111101",
			1012 => "0001010011000100001100",
			1013 => "0001011011111000001000",
			1014 => "0001010100101100000100",
			1015 => "0000000001000000111101",
			1016 => "0000000001000000111101",
			1017 => "0000000001000000111101",
			1018 => "0000000001000000111101",
			1019 => "0000111011000000001000",
			1020 => "0011010101010100000100",
			1021 => "0000000001000000111101",
			1022 => "0000000001000000111101",
			1023 => "0000000001000000111101",
			1024 => "0001000110101100010000",
			1025 => "0010001001010100001000",
			1026 => "0000000001110100000100",
			1027 => "0000000001000000111101",
			1028 => "0000000001000000111101",
			1029 => "0001100101111100000100",
			1030 => "0000000001000000111101",
			1031 => "0000000001000000111101",
			1032 => "0011011010000100000100",
			1033 => "0000000001000000111101",
			1034 => "0000010111011100000100",
			1035 => "0000000001000000111101",
			1036 => "0000000010100100000100",
			1037 => "0000000001000000111101",
			1038 => "0000000001000000111101",
			1039 => "0010001000000001010000",
			1040 => "0011111100111100111000",
			1041 => "0001111100110000010000",
			1042 => "0011010101011100000100",
			1043 => "0000000001000100100001",
			1044 => "0000110011001000001000",
			1045 => "0010100110000000000100",
			1046 => "0000000001000100100001",
			1047 => "0000000001000100100001",
			1048 => "0000000001000100100001",
			1049 => "0000111011000000010100",
			1050 => "0001001100010000010000",
			1051 => "0010101111101000001000",
			1052 => "0011011010100100000100",
			1053 => "0000000001000100100001",
			1054 => "0000000001000100100001",
			1055 => "0000111111101000000100",
			1056 => "0000000001000100100001",
			1057 => "0000000001000100100001",
			1058 => "0000000001000100100001",
			1059 => "0001110011000100001100",
			1060 => "0001111011111000001000",
			1061 => "0001110001010000000100",
			1062 => "0000000001000100100001",
			1063 => "0000000001000100100001",
			1064 => "0000000001000100100001",
			1065 => "0010110011000000000100",
			1066 => "0000000001000100100001",
			1067 => "0000000001000100100001",
			1068 => "0010101011000000001100",
			1069 => "0001001001001000001000",
			1070 => "0001001100101000000100",
			1071 => "0000000001000100100001",
			1072 => "0000000001000100100001",
			1073 => "0000000001000100100001",
			1074 => "0001110000111100001000",
			1075 => "0000111111101000000100",
			1076 => "0000000001000100100001",
			1077 => "0000000001000100100001",
			1078 => "0000000001000100100001",
			1079 => "0011100110110000001100",
			1080 => "0010101111101000000100",
			1081 => "0000000001000100100001",
			1082 => "0001101010001000000100",
			1083 => "0000000001000100100001",
			1084 => "0000000001000100100001",
			1085 => "0000101111001100001000",
			1086 => "0001101101010100000100",
			1087 => "0000000001000100100001",
			1088 => "0000000001000100100001",
			1089 => "0000101110110000000100",
			1090 => "0000000001000100100001",
			1091 => "0001100110011000000100",
			1092 => "0000000001000100100001",
			1093 => "0011110011100000000100",
			1094 => "0000000001000100100001",
			1095 => "0000000001000100100001",
			1096 => "0010001111011000100100",
			1097 => "0001101010001000011100",
			1098 => "0001100010110000010000",
			1099 => "0011010101010100000100",
			1100 => "0000000001000111011101",
			1101 => "0000000110000100000100",
			1102 => "0000000001000111011101",
			1103 => "0011011100101000000100",
			1104 => "0000000001000111011101",
			1105 => "0000000001000111011101",
			1106 => "0001011110010100001000",
			1107 => "0000110011001000000100",
			1108 => "0000000001000111011101",
			1109 => "0000000001000111011101",
			1110 => "0000000001000111011101",
			1111 => "0001001100110000000100",
			1112 => "0000000001000111011101",
			1113 => "0000000001000111011101",
			1114 => "0001110011110100110100",
			1115 => "0000101111001100101100",
			1116 => "0000111111101000011000",
			1117 => "0011011001000100001100",
			1118 => "0011110101111100001000",
			1119 => "0000001110110100000100",
			1120 => "0000000001000111011101",
			1121 => "0000000001000111011101",
			1122 => "0000000001000111011101",
			1123 => "0010011000111000000100",
			1124 => "0000000001000111011101",
			1125 => "0000000001110100000100",
			1126 => "0000000001000111011101",
			1127 => "0000000001000111011101",
			1128 => "0001010011000100000100",
			1129 => "0000000001000111011101",
			1130 => "0000111011000000001000",
			1131 => "0010100011000100000100",
			1132 => "0000000001000111011101",
			1133 => "0000000001000111011101",
			1134 => "0001110011000100000100",
			1135 => "0000000001000111011101",
			1136 => "0000000001000111011101",
			1137 => "0001010110011100000100",
			1138 => "0000000001000111011101",
			1139 => "0000000001000111011101",
			1140 => "0001100100000100000100",
			1141 => "0000000001000111011101",
			1142 => "0000000001000111011101",
			1143 => "0001111100011101010000",
			1144 => "0000101111001101000100",
			1145 => "0010000000110000011000",
			1146 => "0000000100111100010100",
			1147 => "0000100100001000001100",
			1148 => "0010101100010000001000",
			1149 => "0010101000111000000100",
			1150 => "0000000001001010101001",
			1151 => "0000000001001010101001",
			1152 => "0000000001001010101001",
			1153 => "0011111101100000000100",
			1154 => "0000000001001010101001",
			1155 => "0000000001001010101001",
			1156 => "0000000001001010101001",
			1157 => "0010011000000100010100",
			1158 => "0001001010000100001000",
			1159 => "0001111101001000000100",
			1160 => "0000000001001010101001",
			1161 => "0000000001001010101001",
			1162 => "0011101110100100001000",
			1163 => "0000000100011000000100",
			1164 => "0000000001001010101001",
			1165 => "0000000001001010101001",
			1166 => "0000000001001010101001",
			1167 => "0001010011000100010000",
			1168 => "0000111000000000001000",
			1169 => "0011000011000000000100",
			1170 => "0000000001001010101001",
			1171 => "0000000001001010101001",
			1172 => "0011101111010100000100",
			1173 => "0000000001001010101001",
			1174 => "0000000001001010101001",
			1175 => "0000110000111000000100",
			1176 => "0000000001001010101001",
			1177 => "0000000001001010101001",
			1178 => "0011101110010000000100",
			1179 => "0000000001001010101001",
			1180 => "0000111001010100000100",
			1181 => "0000000001001010101001",
			1182 => "0000000001001010101001",
			1183 => "0011000011000000001000",
			1184 => "0010100000111100000100",
			1185 => "0000000001001010101001",
			1186 => "0000000001001010101001",
			1187 => "0011010011000000001000",
			1188 => "0000111011111000000100",
			1189 => "0000000001001010101001",
			1190 => "0000000001001010101001",
			1191 => "0000101011111100000100",
			1192 => "0000000001001010101001",
			1193 => "0000000001001010101001",
			1194 => "0011010111011100001000",
			1195 => "0010000000110000000100",
			1196 => "1111111001001101011101",
			1197 => "0000000001001101011101",
			1198 => "0010011000000100101100",
			1199 => "0000111000101000011000",
			1200 => "0000011110011000010100",
			1201 => "0011100010110000001100",
			1202 => "0010010110000000000100",
			1203 => "1111111001001101011101",
			1204 => "0001101010011000000100",
			1205 => "1111111001001101011101",
			1206 => "0000001001001101011101",
			1207 => "0001001010000100000100",
			1208 => "0000000001001101011101",
			1209 => "1111111001001101011101",
			1210 => "0000001001001101011101",
			1211 => "0010111001001000010000",
			1212 => "0001011000100000000100",
			1213 => "1111111001001101011101",
			1214 => "0010100000111100000100",
			1215 => "0000001001001101011101",
			1216 => "0010010101111000000100",
			1217 => "0000000001001101011101",
			1218 => "1111111001001101011101",
			1219 => "0000001001001101011101",
			1220 => "0001010011000100011100",
			1221 => "0000010111011100010000",
			1222 => "0001011011111000001100",
			1223 => "0000111100110000001000",
			1224 => "0010000011100100000100",
			1225 => "1111111001001101011101",
			1226 => "0000000001001101011101",
			1227 => "0000001001001101011101",
			1228 => "1111111001001101011101",
			1229 => "0000111001010000001000",
			1230 => "0011010101111000000100",
			1231 => "1111111001001101011101",
			1232 => "0000000001001101011101",
			1233 => "0000001001001101011101",
			1234 => "0000110000111000001000",
			1235 => "0010000011001000000100",
			1236 => "0000000001001101011101",
			1237 => "0000001001001101011101",
			1238 => "1111111001001101011101",
			1239 => "0001111100011101011000",
			1240 => "0010000011100101000100",
			1241 => "0000111000101000101000",
			1242 => "0011110101111100010100",
			1243 => "0011111100111000010000",
			1244 => "0010010110000000001000",
			1245 => "0001010101111000000100",
			1246 => "0000000001010000111001",
			1247 => "0000000001010000111001",
			1248 => "0011111010011000000100",
			1249 => "0000000001010000111001",
			1250 => "0000000001010000111001",
			1251 => "0000000001010000111001",
			1252 => "0011110101100100001000",
			1253 => "0001111011111000000100",
			1254 => "0000000001010000111001",
			1255 => "0000000001010000111001",
			1256 => "0000001001101000001000",
			1257 => "0000111100110000000100",
			1258 => "0000000001010000111001",
			1259 => "0000000001010000111001",
			1260 => "0000000001010000111001",
			1261 => "0010100011000100001100",
			1262 => "0000001101011100001000",
			1263 => "0011111110010000000100",
			1264 => "0000000001010000111001",
			1265 => "0000000001010000111001",
			1266 => "1111111001010000111001",
			1267 => "0001011001000000000100",
			1268 => "0000000001010000111001",
			1269 => "0010110101101100000100",
			1270 => "0000000001010000111001",
			1271 => "0010011000111000000100",
			1272 => "0000000001010000111001",
			1273 => "0000000001010000111001",
			1274 => "0011010101101100000100",
			1275 => "0000000001010000111001",
			1276 => "0010101001010100000100",
			1277 => "0000000001010000111001",
			1278 => "0000001110110000001000",
			1279 => "0011000101111000000100",
			1280 => "0000000001010000111001",
			1281 => "0000000001010000111001",
			1282 => "0000000001010000111001",
			1283 => "0011000011000000001000",
			1284 => "0011110100111100000100",
			1285 => "0000000001010000111001",
			1286 => "0000000001010000111001",
			1287 => "0011010011000000001000",
			1288 => "0010011101001000000100",
			1289 => "0000000001010000111001",
			1290 => "0000000001010000111001",
			1291 => "0000101011111100000100",
			1292 => "0000000001010000111001",
			1293 => "0000000001010000111001",
			1294 => "0001110011110101011100",
			1295 => "0000111000101000101000",
			1296 => "0000111100110000011000",
			1297 => "0000010011010000010000",
			1298 => "0010011001000100000100",
			1299 => "0000000001010100001101",
			1300 => "0000001011100100001000",
			1301 => "0000100100001000000100",
			1302 => "0000000001010100001101",
			1303 => "0000000001010100001101",
			1304 => "0000000001010100001101",
			1305 => "0001001001000100000100",
			1306 => "0000000001010100001101",
			1307 => "1111111001010100001101",
			1308 => "0010010011000000000100",
			1309 => "0000000001010100001101",
			1310 => "0001000110000000000100",
			1311 => "0000000001010100001101",
			1312 => "0001010110011100000100",
			1313 => "0000001001010100001101",
			1314 => "0000000001010100001101",
			1315 => "0001011000100000010100",
			1316 => "0010000011100100010000",
			1317 => "0011101110100000001100",
			1318 => "0011111110010000000100",
			1319 => "0000000001010100001101",
			1320 => "0000001011100100000100",
			1321 => "0000000001010100001101",
			1322 => "0000000001010100001101",
			1323 => "1111111001010100001101",
			1324 => "0000000001010100001101",
			1325 => "0000111011000000001000",
			1326 => "0010011010000100000100",
			1327 => "0000000001010100001101",
			1328 => "0000001001010100001101",
			1329 => "0011001101101000001100",
			1330 => "0000001100100100001000",
			1331 => "0000001110110100000100",
			1332 => "0000000001010100001101",
			1333 => "0000000001010100001101",
			1334 => "0000000001010100001101",
			1335 => "0001011010100000001000",
			1336 => "0011101100011000000100",
			1337 => "0000000001010100001101",
			1338 => "0000000001010100001101",
			1339 => "0000000001010100001101",
			1340 => "0011000011000000000100",
			1341 => "0000001001010100001101",
			1342 => "0001011011000000000100",
			1343 => "0000000001010100001101",
			1344 => "0000110101110000000100",
			1345 => "0000000001010100001101",
			1346 => "0000000001010100001101",
			1347 => "0001110011110101010000",
			1348 => "0011110000001100100100",
			1349 => "0001111100010000000100",
			1350 => "1111111001010111010001",
			1351 => "0001000110000000001100",
			1352 => "0010010110000000000100",
			1353 => "0000000001010111010001",
			1354 => "0011001001001000000100",
			1355 => "0000000001010111010001",
			1356 => "0000000001010111010001",
			1357 => "0001000110011100001100",
			1358 => "0000011001100000000100",
			1359 => "0000000001010111010001",
			1360 => "0001101010001100000100",
			1361 => "0000000001010111010001",
			1362 => "0000001001010111010001",
			1363 => "0011110001100000000100",
			1364 => "0000000001010111010001",
			1365 => "0000000001010111010001",
			1366 => "0001111011111000000100",
			1367 => "1111111001010111010001",
			1368 => "0001000011000000010000",
			1369 => "0001001010000100001100",
			1370 => "0010101111101000001000",
			1371 => "0001000101010100000100",
			1372 => "0000000001010111010001",
			1373 => "0000001001010111010001",
			1374 => "0000000001010111010001",
			1375 => "1111111001010111010001",
			1376 => "0001001100000000001000",
			1377 => "0000101111001100000100",
			1378 => "0000001001010111010001",
			1379 => "0000000001010111010001",
			1380 => "0010000011100100001000",
			1381 => "0001011000100000000100",
			1382 => "1111111001010111010001",
			1383 => "0000000001010111010001",
			1384 => "0011011010000100000100",
			1385 => "0000001001010111010001",
			1386 => "0000000001010111010001",
			1387 => "0011000011000000000100",
			1388 => "0000001001010111010001",
			1389 => "0011010011000000001000",
			1390 => "0001011010011100000100",
			1391 => "0000000001010111010001",
			1392 => "0000000001010111010001",
			1393 => "0000101011111100000100",
			1394 => "0000000001010111010001",
			1395 => "0000000001010111010001",
			1396 => "0001111100011101011000",
			1397 => "0000101111001101001100",
			1398 => "0010000000110000100000",
			1399 => "0000000100111100010100",
			1400 => "0000100100001000001100",
			1401 => "0010101100010000001000",
			1402 => "0010101000111000000100",
			1403 => "0000000001011010101101",
			1404 => "0000000001011010101101",
			1405 => "0000000001011010101101",
			1406 => "0011111101100000000100",
			1407 => "0000000001011010101101",
			1408 => "0000000001011010101101",
			1409 => "0001100001000000001000",
			1410 => "0001100110110000000100",
			1411 => "0000000001011010101101",
			1412 => "0000000001011010101101",
			1413 => "0000000001011010101101",
			1414 => "0011011001000100011100",
			1415 => "0011110000000100010000",
			1416 => "0010101001010100001000",
			1417 => "0001111101001000000100",
			1418 => "0000000001011010101101",
			1419 => "0000000001011010101101",
			1420 => "0011010101101100000100",
			1421 => "0000000001011010101101",
			1422 => "0000000001011010101101",
			1423 => "0001111001011000000100",
			1424 => "0000000001011010101101",
			1425 => "0000111111101000000100",
			1426 => "0000000001011010101101",
			1427 => "0000000001011010101101",
			1428 => "0011111001111000001100",
			1429 => "0000110000111000001000",
			1430 => "0001101100011000000100",
			1431 => "0000000001011010101101",
			1432 => "0000000001011010101101",
			1433 => "0000000001011010101101",
			1434 => "0000000001011010101101",
			1435 => "0011101110010000000100",
			1436 => "0000000001011010101101",
			1437 => "0000111001010100000100",
			1438 => "0000000001011010101101",
			1439 => "0000000001011010101101",
			1440 => "0011000011000000001000",
			1441 => "0010100000111100000100",
			1442 => "0000000001011010101101",
			1443 => "0000000001011010101101",
			1444 => "0011010011000000001000",
			1445 => "0000111011111000000100",
			1446 => "0000000001011010101101",
			1447 => "0000000001011010101101",
			1448 => "0000101011111100000100",
			1449 => "0000000001011010101101",
			1450 => "0000000001011010101101",
			1451 => "0010001111001000000100",
			1452 => "1111111001011101001001",
			1453 => "0000001101011100100100",
			1454 => "0001111100010000000100",
			1455 => "1111111001011101001001",
			1456 => "0010101001011000010100",
			1457 => "0001000110000000001100",
			1458 => "0010101000000000001000",
			1459 => "0001011101101000000100",
			1460 => "0000000001011101001001",
			1461 => "0000000001011101001001",
			1462 => "0000000001011101001001",
			1463 => "0001100010110000000100",
			1464 => "0000000001011101001001",
			1465 => "0000001001011101001001",
			1466 => "0001000110101100000100",
			1467 => "0000000001011101001001",
			1468 => "0001000011000100000100",
			1469 => "0000000001011101001001",
			1470 => "0000000001011101001001",
			1471 => "0010001111011000001000",
			1472 => "0000001000001100000100",
			1473 => "1111111001011101001001",
			1474 => "0000000001011101001001",
			1475 => "0010010110101100011000",
			1476 => "0001010011000100001100",
			1477 => "0001010110011100001000",
			1478 => "0011011001000100000100",
			1479 => "0000000001011101001001",
			1480 => "0000000001011101001001",
			1481 => "1111111001011101001001",
			1482 => "0001110000111100001000",
			1483 => "0001010001011000000100",
			1484 => "0000000001011101001001",
			1485 => "0000000001011101001001",
			1486 => "0000001001011101001001",
			1487 => "0011110000001000000100",
			1488 => "0000000001011101001001",
			1489 => "0000001001011101001001",
			1490 => "0010011001000100000100",
			1491 => "1111111001011111100101",
			1492 => "0000111000000000010000",
			1493 => "0001101010011000000100",
			1494 => "0000000001011111100101",
			1495 => "0010001111001000000100",
			1496 => "0000000001011111100101",
			1497 => "0000000110100100000100",
			1498 => "0000001001011111100101",
			1499 => "0000000001011111100101",
			1500 => "0010000000110000010100",
			1501 => "0010111010100100000100",
			1502 => "0000000001011111100101",
			1503 => "0001110001011000001100",
			1504 => "0010101000101000001000",
			1505 => "0000111100110000000100",
			1506 => "0000000001011111100101",
			1507 => "0000000001011111100101",
			1508 => "1111111001011111100101",
			1509 => "0000000001011111100101",
			1510 => "0001000011000000001100",
			1511 => "0001001010000100001000",
			1512 => "0010101111101000000100",
			1513 => "0000001001011111100101",
			1514 => "0000000001011111100101",
			1515 => "1111111001011111100101",
			1516 => "0001111011000000001100",
			1517 => "0001101110010000001000",
			1518 => "0011111010011000000100",
			1519 => "0000000001011111100101",
			1520 => "0000000001011111100101",
			1521 => "1111111001011111100101",
			1522 => "0000100111111000001000",
			1523 => "0000110011000100000100",
			1524 => "0000001001011111100101",
			1525 => "0000000001011111100101",
			1526 => "0000010101011100000100",
			1527 => "0000000001011111100101",
			1528 => "0000001001011111100101",
			1529 => "0011010111011100001000",
			1530 => "0010000000110000000100",
			1531 => "1111111001100010010001",
			1532 => "0000000001100010010001",
			1533 => "0001111100011101000000",
			1534 => "0000101111001100111000",
			1535 => "0010011000000100011000",
			1536 => "0000111100101100010000",
			1537 => "0010010011001000001000",
			1538 => "0001100100011100000100",
			1539 => "0000001001100010010001",
			1540 => "0000000001100010010001",
			1541 => "0000001000100100000100",
			1542 => "0000000001100010010001",
			1543 => "0000001001100010010001",
			1544 => "0000110000111100000100",
			1545 => "1111111001100010010001",
			1546 => "0000000001100010010001",
			1547 => "0001000011000000010000",
			1548 => "0011011101101000001000",
			1549 => "0011000011000000000100",
			1550 => "1111111001100010010001",
			1551 => "0000000001100010010001",
			1552 => "0011000011001000000100",
			1553 => "0000001001100010010001",
			1554 => "0000000001100010010001",
			1555 => "0010000011100100001000",
			1556 => "0011000110000000000100",
			1557 => "0000000001100010010001",
			1558 => "1111111001100010010001",
			1559 => "0011000101111000000100",
			1560 => "0000001001100010010001",
			1561 => "1111111001100010010001",
			1562 => "0001101110000100000100",
			1563 => "1111111001100010010001",
			1564 => "0000000001100010010001",
			1565 => "0001011011000000001000",
			1566 => "0001101100111100000100",
			1567 => "0000001001100010010001",
			1568 => "0000000001100010010001",
			1569 => "0000111010100000000100",
			1570 => "0000001001100010010001",
			1571 => "0000000001100010010001",
			1572 => "0011010011000001000100",
			1573 => "0001111100010000000100",
			1574 => "1111111001100100100101",
			1575 => "0011111100111000011100",
			1576 => "0001100011101100010000",
			1577 => "0011101010011000001100",
			1578 => "0000111000101000001000",
			1579 => "0011001001001000000100",
			1580 => "0000001001100100100101",
			1581 => "0000000001100100100101",
			1582 => "0000000001100100100101",
			1583 => "1111111001100100100101",
			1584 => "0000011001100000000100",
			1585 => "0000000001100100100101",
			1586 => "0001010001111100000100",
			1587 => "0000001001100100100101",
			1588 => "0000000001100100100101",
			1589 => "0001111011111000000100",
			1590 => "1111111001100100100101",
			1591 => "0000111001010000010000",
			1592 => "0010000011001000001000",
			1593 => "0000001100001000000100",
			1594 => "0000000001100100100101",
			1595 => "0000001001100100100101",
			1596 => "0010001000000000000100",
			1597 => "1111111001100100100101",
			1598 => "0000000001100100100101",
			1599 => "0010000011100100001000",
			1600 => "0001001100000000000100",
			1601 => "0000000001100100100101",
			1602 => "0000000001100100100101",
			1603 => "0010101110111000000100",
			1604 => "0000001001100100100101",
			1605 => "0000000001100100100101",
			1606 => "0001101000101100000100",
			1607 => "0000000001100100100101",
			1608 => "0000001001100100100101",
			1609 => "0001111100011101100100",
			1610 => "0010000011100101001100",
			1611 => "0000111000101000110000",
			1612 => "0011101101100100011100",
			1613 => "0011111100111000010000",
			1614 => "0010010110000000001000",
			1615 => "0001010101111000000100",
			1616 => "0000000001101000010001",
			1617 => "0000000001101000010001",
			1618 => "0011111010011000000100",
			1619 => "0000000001101000010001",
			1620 => "0000000001101000010001",
			1621 => "0000011101000000001000",
			1622 => "0000011001100000000100",
			1623 => "0000000001101000010001",
			1624 => "0000000001101000010001",
			1625 => "0000000001101000010001",
			1626 => "0011110101100100001000",
			1627 => "0011000111011100000100",
			1628 => "0000000001101000010001",
			1629 => "0000000001101000010001",
			1630 => "0000001001101000001000",
			1631 => "0000111100110000000100",
			1632 => "0000000001101000010001",
			1633 => "0000000001101000010001",
			1634 => "0000000001101000010001",
			1635 => "0010100011000100001100",
			1636 => "0000001101011100001000",
			1637 => "0011111110010000000100",
			1638 => "0000000001101000010001",
			1639 => "0000000001101000010001",
			1640 => "1111111001101000010001",
			1641 => "0001011001000000000100",
			1642 => "0000000001101000010001",
			1643 => "0010110101101100000100",
			1644 => "0000000001101000010001",
			1645 => "0010011000111000000100",
			1646 => "0000000001101000010001",
			1647 => "0000000001101000010001",
			1648 => "0011010101101100000100",
			1649 => "0000000001101000010001",
			1650 => "0010101001010100000100",
			1651 => "0000000001101000010001",
			1652 => "0001111110111000001100",
			1653 => "0010100001101000001000",
			1654 => "0001001000000000000100",
			1655 => "0000000001101000010001",
			1656 => "0000000001101000010001",
			1657 => "0000000001101000010001",
			1658 => "0000000001101000010001",
			1659 => "0011000011000000000100",
			1660 => "0000000001101000010001",
			1661 => "0011010011000000001000",
			1662 => "0010011101001000000100",
			1663 => "0000000001101000010001",
			1664 => "0000000001101000010001",
			1665 => "0000101011111100000100",
			1666 => "0000000001101000010001",
			1667 => "0000000001101000010001",
			1668 => "0010011001000100000100",
			1669 => "1111111001101011001111",
			1670 => "0000111000000000001100",
			1671 => "0001101010011000000100",
			1672 => "0000000001101011001111",
			1673 => "0010001111001000000100",
			1674 => "0000000001101011001111",
			1675 => "0000001001101011001111",
			1676 => "0001010001001000101100",
			1677 => "0000101111101100011000",
			1678 => "0001011001010100001000",
			1679 => "0010111001001000000100",
			1680 => "0000000001101011001111",
			1681 => "1111111001101011001111",
			1682 => "0011101110100100001000",
			1683 => "0001011000101000000100",
			1684 => "0000001001101011001111",
			1685 => "0000000001101011001111",
			1686 => "0001011011000000000100",
			1687 => "0000001001101011001111",
			1688 => "0000000001101011001111",
			1689 => "0011011001001000000100",
			1690 => "1111111001101011001111",
			1691 => "0000111001010000001000",
			1692 => "0011010011000000000100",
			1693 => "1111111001101011001111",
			1694 => "0000001001101011001111",
			1695 => "0000111111101000000100",
			1696 => "0000001001101011001111",
			1697 => "0000000001101011001111",
			1698 => "0000111011000000001100",
			1699 => "0010011010000100000100",
			1700 => "0000000001101011001111",
			1701 => "0010001111011000000100",
			1702 => "0000000001101011001111",
			1703 => "0000001001101011001111",
			1704 => "0001110000111100010000",
			1705 => "0010111001001000001000",
			1706 => "0001111011111000000100",
			1707 => "0000000001101011001111",
			1708 => "1111111001101011001111",
			1709 => "0011110100110000000100",
			1710 => "0000000001101011001111",
			1711 => "0000000001101011001111",
			1712 => "0000110001010100000100",
			1713 => "0000001001101011001111",
			1714 => "0000000001101011001111",
			1715 => "0000010110001100100000",
			1716 => "0010000000110000010000",
			1717 => "0000010011110000000100",
			1718 => "1111111001101101010001",
			1719 => "0010111010100100001000",
			1720 => "0010111110011000000100",
			1721 => "1111111001101101010001",
			1722 => "0000000001101101010001",
			1723 => "1111111001101101010001",
			1724 => "0011001001001000001000",
			1725 => "0011111101010100000100",
			1726 => "0000010001101101010001",
			1727 => "0000000001101101010001",
			1728 => "0011001001000100000100",
			1729 => "0000000001101101010001",
			1730 => "1111111001101101010001",
			1731 => "0011111110100000001000",
			1732 => "0010011111011000000100",
			1733 => "0000001001101101010001",
			1734 => "1111111001101101010001",
			1735 => "0011010101011100000100",
			1736 => "0000000001101101010001",
			1737 => "0010101100001100010100",
			1738 => "0001011000100000001100",
			1739 => "0000001101011100000100",
			1740 => "0000010001101101010001",
			1741 => "0010000011100100000100",
			1742 => "0000000001101101010001",
			1743 => "0000001001101101010001",
			1744 => "0010000011100100000100",
			1745 => "0000010001101101010001",
			1746 => "0000001001101101010001",
			1747 => "0000001001101101010001",
			1748 => "0000010011110000001000",
			1749 => "0010001111011000000100",
			1750 => "1111111001101111000101",
			1751 => "0000001001101111000101",
			1752 => "0001111100011100100100",
			1753 => "0000101111001100011000",
			1754 => "0001101010001100000100",
			1755 => "1111111001101111000101",
			1756 => "0000000100110100000100",
			1757 => "0000001001101111000101",
			1758 => "0010000011100100001000",
			1759 => "0001001010000100000100",
			1760 => "0000000001101111000101",
			1761 => "0000000001101111000101",
			1762 => "0011000101111000000100",
			1763 => "0000001001101111000101",
			1764 => "1111111001101111000101",
			1765 => "0000001111010000001000",
			1766 => "0011110000101100000100",
			1767 => "1111111001101111000101",
			1768 => "1111111001101111000101",
			1769 => "0000000001101111000101",
			1770 => "0001011011000000001000",
			1771 => "0001111110001100000100",
			1772 => "0000000001101111000101",
			1773 => "0000001001101111000101",
			1774 => "0000111010100000000100",
			1775 => "0000001001101111000101",
			1776 => "1111111001101111000101",
			1777 => "0000011110011000110000",
			1778 => "0000010110001100100000",
			1779 => "0000011101000000010100",
			1780 => "0000010011110000001000",
			1781 => "0010001111011000000100",
			1782 => "1111111001110001101001",
			1783 => "1111111001110001101001",
			1784 => "0011110100010000000100",
			1785 => "1111111001110001101001",
			1786 => "0001100000010000000100",
			1787 => "0000001001110001101001",
			1788 => "1111111001110001101001",
			1789 => "0011111101100000000100",
			1790 => "1111111001110001101001",
			1791 => "0000000000000000000100",
			1792 => "0000001001110001101001",
			1793 => "0000000001110001101001",
			1794 => "0011111101100000001000",
			1795 => "0001101010011000000100",
			1796 => "1111111001110001101001",
			1797 => "0000000001110001101001",
			1798 => "0001010011000100000100",
			1799 => "0000000001110001101001",
			1800 => "0000010001110001101001",
			1801 => "0011110011101000001000",
			1802 => "0010011101001000000100",
			1803 => "0000000001110001101001",
			1804 => "1111111001110001101001",
			1805 => "0010111100101000000100",
			1806 => "0000001001110001101001",
			1807 => "0000111100110000001000",
			1808 => "0011011101101000000100",
			1809 => "0000001001110001101001",
			1810 => "0000011001110001101001",
			1811 => "0000001110110000000100",
			1812 => "0000011001110001101001",
			1813 => "0011101110010000000100",
			1814 => "0000010001110001101001",
			1815 => "0000111000101000000100",
			1816 => "0000010001110001101001",
			1817 => "0000011001110001101001",
			1818 => "0010000011100100110100",
			1819 => "0000100110010100100100",
			1820 => "0000101010101000011000",
			1821 => "0011110000001100010100",
			1822 => "0001111100010000000100",
			1823 => "1111111001110100010101",
			1824 => "0000111000101000001000",
			1825 => "0001000110000000000100",
			1826 => "0000000001110100010101",
			1827 => "0000001001110100010101",
			1828 => "0011111110010000000100",
			1829 => "0000000001110100010101",
			1830 => "0000000001110100010101",
			1831 => "1111111001110100010101",
			1832 => "0001101101010000001000",
			1833 => "0001110100101100000100",
			1834 => "0000000001110100010101",
			1835 => "0000001001110100010101",
			1836 => "1111111001110100010101",
			1837 => "0011011001001000001000",
			1838 => "0001010001001000000100",
			1839 => "1111111001110100010101",
			1840 => "0000000001110100010101",
			1841 => "0011001001000100000100",
			1842 => "0000000001110100010101",
			1843 => "0000000001110100010101",
			1844 => "0010100000111100011000",
			1845 => "0000101111001100010000",
			1846 => "0011101111110100001000",
			1847 => "0001111011000000000100",
			1848 => "0000000001110100010101",
			1849 => "0000000001110100010101",
			1850 => "0001100101111100000100",
			1851 => "0000001001110100010101",
			1852 => "0000000001110100010101",
			1853 => "0000111001010000000100",
			1854 => "0000000001110100010101",
			1855 => "0000001001110100010101",
			1856 => "0001011110111000000100",
			1857 => "1111111001110100010101",
			1858 => "0000110000111000000100",
			1859 => "0000000001110100010101",
			1860 => "0000000001110100010101",
			1861 => "0010101111101000100000",
			1862 => "0010010110000000001100",
			1863 => "0000000000000100001000",
			1864 => "0001100010110000000100",
			1865 => "0000000001110111010001",
			1866 => "0000000001110111010001",
			1867 => "0000000001110111010001",
			1868 => "0001101010011000000100",
			1869 => "0000000001110111010001",
			1870 => "0011010111011100000100",
			1871 => "0000000001110111010001",
			1872 => "0001011011111000001000",
			1873 => "0000101011001100000100",
			1874 => "0000000001110111010001",
			1875 => "0000000001110111010001",
			1876 => "0000000001110111010001",
			1877 => "0001010011000100011100",
			1878 => "0000101100001000010000",
			1879 => "0001101100000100001000",
			1880 => "0001111001010100000100",
			1881 => "0000000001110111010001",
			1882 => "0000000001110111010001",
			1883 => "0010001010000100000100",
			1884 => "0000000001110111010001",
			1885 => "0000000001110111010001",
			1886 => "0010010110101100001000",
			1887 => "0011100101100000000100",
			1888 => "0000000001110111010001",
			1889 => "0000000001110111010001",
			1890 => "0000000001110111010001",
			1891 => "0000111011000000010000",
			1892 => "0010010101111000001000",
			1893 => "0011110111000000000100",
			1894 => "0000000001110111010001",
			1895 => "0000000001110111010001",
			1896 => "0000001111010000000100",
			1897 => "0000000001110111010001",
			1898 => "0000000001110111010001",
			1899 => "0001101110000100010000",
			1900 => "0000010011010000001000",
			1901 => "0010101000100000000100",
			1902 => "0000000001110111010001",
			1903 => "0000000001110111010001",
			1904 => "0010100000111000000100",
			1905 => "0000000001110111010001",
			1906 => "0000000001110111010001",
			1907 => "0000000001110111010001",
			1908 => "0011010111011100001100",
			1909 => "0010001111001000000100",
			1910 => "1111111001111000111101",
			1911 => "0001010101111000000100",
			1912 => "0000001001111000111101",
			1913 => "1111111001111000111101",
			1914 => "0011111010011000000100",
			1915 => "1111111001111000111101",
			1916 => "0000110000111000100100",
			1917 => "0001111100011100010100",
			1918 => "0000101111001100001100",
			1919 => "0000000100110100000100",
			1920 => "0000001001111000111101",
			1921 => "0010011010000100000100",
			1922 => "1111111001111000111101",
			1923 => "0000000001111000111101",
			1924 => "0001101110000100000100",
			1925 => "1111111001111000111101",
			1926 => "0000000001111000111101",
			1927 => "0011111110011100001000",
			1928 => "0010110110000000000100",
			1929 => "0000001001111000111101",
			1930 => "0000001001111000111101",
			1931 => "0001000110101100000100",
			1932 => "0000001001111000111101",
			1933 => "0000000001111000111101",
			1934 => "1111111001111000111101",
			1935 => "0011010111011100010000",
			1936 => "0010011111011000001000",
			1937 => "0010000000110000000100",
			1938 => "1111111001111011010001",
			1939 => "0000000001111011010001",
			1940 => "0001011110001100000100",
			1941 => "0000000001111011010001",
			1942 => "0000000001111011010001",
			1943 => "0010100000111100101000",
			1944 => "0001010001001000100000",
			1945 => "0011010011000000011000",
			1946 => "0000101011001100010000",
			1947 => "0010001000000000001000",
			1948 => "0011000110000000000100",
			1949 => "0000000001111011010001",
			1950 => "1111111001111011010001",
			1951 => "0011100110110000000100",
			1952 => "0000000001111011010001",
			1953 => "0000001001111011010001",
			1954 => "0001111110111000000100",
			1955 => "1111111001111011010001",
			1956 => "0000000001111011010001",
			1957 => "0000000010101100000100",
			1958 => "0000000001111011010001",
			1959 => "0000001001111011010001",
			1960 => "0011110100100000000100",
			1961 => "0000000001111011010001",
			1962 => "0000001001111011010001",
			1963 => "0011101110010000010000",
			1964 => "0000001111001100001100",
			1965 => "0011011001001000000100",
			1966 => "1111111001111011010001",
			1967 => "0000110000111000000100",
			1968 => "0000001001111011010001",
			1969 => "1111111001111011010001",
			1970 => "1111111001111011010001",
			1971 => "0000001001111011010001",
			1972 => "0011010111011100010000",
			1973 => "0010001111001000000100",
			1974 => "1111111001111101000101",
			1975 => "0001010011001000000100",
			1976 => "0000001001111101000101",
			1977 => "0001010110011100000100",
			1978 => "1111111001111101000101",
			1979 => "0000000001111101000101",
			1980 => "0011111010011000000100",
			1981 => "1111111001111101000101",
			1982 => "0001010101110000100100",
			1983 => "0001010011000100010000",
			1984 => "0011110000001100000100",
			1985 => "0000001001111101000101",
			1986 => "0010010011000000000100",
			1987 => "1111111001111101000101",
			1988 => "0001010110011100000100",
			1989 => "0000000001111101000101",
			1990 => "1111111001111101000101",
			1991 => "0001110011000100001100",
			1992 => "0000111100101100000100",
			1993 => "0000000001111101000101",
			1994 => "0000110000111100000100",
			1995 => "1111111001111101000101",
			1996 => "0000000001111101000101",
			1997 => "0010101100001100000100",
			1998 => "0000001001111101000101",
			1999 => "0000000001111101000101",
			2000 => "1111111001111101000101",
			2001 => "0000010110001100100000",
			2002 => "0010000000110000010000",
			2003 => "0000010011110000000100",
			2004 => "1111111001111111011001",
			2005 => "0010110111011100001000",
			2006 => "0010011001000100000100",
			2007 => "1111111001111111011001",
			2008 => "0000001001111111011001",
			2009 => "1111111001111111011001",
			2010 => "0011001001000100001100",
			2011 => "0001111101001000000100",
			2012 => "1111111001111111011001",
			2013 => "0000100110111100000100",
			2014 => "0000001001111111011001",
			2015 => "0000000001111111011001",
			2016 => "1111111001111111011001",
			2017 => "0011111111010100001000",
			2018 => "0010110101101100000100",
			2019 => "0000000001111111011001",
			2020 => "1111111001111111011001",
			2021 => "0011010101011100000100",
			2022 => "0000000001111111011001",
			2023 => "0001000011000100011100",
			2024 => "0001010011000100010000",
			2025 => "0000101111001100001000",
			2026 => "0000111000101000000100",
			2027 => "0000001001111111011001",
			2028 => "0000000001111111011001",
			2029 => "0011011101101000000100",
			2030 => "1111111001111111011001",
			2031 => "0000001001111111011001",
			2032 => "0011000101101100000100",
			2033 => "0000001001111111011001",
			2034 => "0000010111011100000100",
			2035 => "0000001001111111011001",
			2036 => "0000001001111111011001",
			2037 => "0000000001111111011001",
			2038 => "0010101111101000100000",
			2039 => "0010010110000000001100",
			2040 => "0000000000000100001000",
			2041 => "0001100010110000000100",
			2042 => "0000000010000010100101",
			2043 => "0000000010000010100101",
			2044 => "0000000010000010100101",
			2045 => "0001101010011000000100",
			2046 => "0000000010000010100101",
			2047 => "0011010111011100000100",
			2048 => "0000000010000010100101",
			2049 => "0001011011111000001000",
			2050 => "0000101011001100000100",
			2051 => "0000000010000010100101",
			2052 => "0000000010000010100101",
			2053 => "0000000010000010100101",
			2054 => "0001010011000100100000",
			2055 => "0000101100001000010000",
			2056 => "0001101100000100001000",
			2057 => "0001111001010100000100",
			2058 => "0000000010000010100101",
			2059 => "0000000010000010100101",
			2060 => "0001010001010000000100",
			2061 => "0000000010000010100101",
			2062 => "0000000010000010100101",
			2063 => "0010010110101100001100",
			2064 => "0001011011111000001000",
			2065 => "0001010001010000000100",
			2066 => "0000000010000010100101",
			2067 => "0000000010000010100101",
			2068 => "0000000010000010100101",
			2069 => "0000000010000010100101",
			2070 => "0000111011000000010100",
			2071 => "0010010101111000001000",
			2072 => "0011110111000000000100",
			2073 => "0000000010000010100101",
			2074 => "0000000010000010100101",
			2075 => "0000010101010100000100",
			2076 => "0000000010000010100101",
			2077 => "0000001000001100000100",
			2078 => "0000000010000010100101",
			2079 => "0000000010000010100101",
			2080 => "0001101110000100010000",
			2081 => "0000010011010000001000",
			2082 => "0010101000100000000100",
			2083 => "0000000010000010100101",
			2084 => "0000000010000010100101",
			2085 => "0010100000111000000100",
			2086 => "0000000010000010100101",
			2087 => "0000000010000010100101",
			2088 => "0000000010000010100101",
			2089 => "0011010111011100010000",
			2090 => "0001010101111000001000",
			2091 => "0010101000000000000100",
			2092 => "0000000010000101010001",
			2093 => "0000000010000101010001",
			2094 => "0010011111011000000100",
			2095 => "0000000010000101010001",
			2096 => "0000000010000101010001",
			2097 => "0001000110101100101100",
			2098 => "0011011101101000100100",
			2099 => "0011000110000000010100",
			2100 => "0000101111001100010000",
			2101 => "0010001111011000001000",
			2102 => "0011000101011100000100",
			2103 => "0000000010000101010001",
			2104 => "0000000010000101010001",
			2105 => "0011101110100100000100",
			2106 => "0000000010000101010001",
			2107 => "0000000010000101010001",
			2108 => "0000000010000101010001",
			2109 => "0010101101001000001000",
			2110 => "0001111011111000000100",
			2111 => "0000000010000101010001",
			2112 => "0000000010000101010001",
			2113 => "0011111001111000000100",
			2114 => "0000000010000101010001",
			2115 => "0000000010000101010001",
			2116 => "0000000001110100000100",
			2117 => "0000000010000101010001",
			2118 => "0000000010000101010001",
			2119 => "0001001001010000001100",
			2120 => "0000010101011100001000",
			2121 => "0000000110111100000100",
			2122 => "0000000010000101010001",
			2123 => "0000000010000101010001",
			2124 => "0000000010000101010001",
			2125 => "0000110011110100001000",
			2126 => "0000001110110100000100",
			2127 => "0000000010000101010001",
			2128 => "0000000010000101010001",
			2129 => "0000010111011100000100",
			2130 => "0000000010000101010001",
			2131 => "0000000010000101010001",
			2132 => "0011010111011100010100",
			2133 => "0001010011001000001100",
			2134 => "0010011001000100000100",
			2135 => "0000000010000111101101",
			2136 => "0010101000000100000100",
			2137 => "0000000010000111101101",
			2138 => "0000000010000111101101",
			2139 => "0010011111011000000100",
			2140 => "0000000010000111101101",
			2141 => "0000000010000111101101",
			2142 => "0010101100001100110100",
			2143 => "0001011000100000100100",
			2144 => "0001001000111000011100",
			2145 => "0011011101101000010000",
			2146 => "0000100100010100001000",
			2147 => "0011110000000100000100",
			2148 => "0000000010000111101101",
			2149 => "0000000010000111101101",
			2150 => "0001011011111000000100",
			2151 => "0000000010000111101101",
			2152 => "0000000010000111101101",
			2153 => "0010001001010100001000",
			2154 => "0000000001110100000100",
			2155 => "0000000010000111101101",
			2156 => "0000000010000111101101",
			2157 => "0000000010000111101101",
			2158 => "0000010111011100000100",
			2159 => "0000000010000111101101",
			2160 => "0000000010000111101101",
			2161 => "0011110000000100001000",
			2162 => "0011011001001000000100",
			2163 => "0000000010000111101101",
			2164 => "0000000010000111101101",
			2165 => "0001101000001000000100",
			2166 => "0000000010000111101101",
			2167 => "0000000010000111101101",
			2168 => "0001111010011100000100",
			2169 => "0000000010000111101101",
			2170 => "0000000010000111101101",
			2171 => "0001110011110100111000",
			2172 => "0000101111001100101100",
			2173 => "0011110101100100100100",
			2174 => "0000001110110000100000",
			2175 => "0001110001001000010000",
			2176 => "0000100110010100001000",
			2177 => "0011110000000100000100",
			2178 => "0000000010001001111001",
			2179 => "0000000010001001111001",
			2180 => "0010100011000100000100",
			2181 => "0000000010001001111001",
			2182 => "0000000010001001111001",
			2183 => "0000001000010000001000",
			2184 => "0000001100001000000100",
			2185 => "0000000010001001111001",
			2186 => "0000000010001001111001",
			2187 => "0010011100010000000100",
			2188 => "0000000010001001111001",
			2189 => "0000000010001001111001",
			2190 => "0000000010001001111001",
			2191 => "0011000111011100000100",
			2192 => "0000000010001001111001",
			2193 => "0000000010001001111001",
			2194 => "0000111001010000000100",
			2195 => "0000000010001001111001",
			2196 => "0001101110000100000100",
			2197 => "0000000010001001111001",
			2198 => "0000000010001001111001",
			2199 => "0001100101100000000100",
			2200 => "0000000010001001111001",
			2201 => "0000011100101000000100",
			2202 => "0000000010001001111001",
			2203 => "0000010101101100000100",
			2204 => "0000000010001001111001",
			2205 => "0000000010001001111001",
			2206 => "0011010111011100001000",
			2207 => "0010000000110000000100",
			2208 => "1111111010001011110101",
			2209 => "0000000010001011110101",
			2210 => "0010000110101100110000",
			2211 => "0011000011000000011000",
			2212 => "0001111110111000010100",
			2213 => "0000101111001100010000",
			2214 => "0000111011000000001000",
			2215 => "0010100011000100000100",
			2216 => "0000000010001011110101",
			2217 => "0000001010001011110101",
			2218 => "0011011001001000000100",
			2219 => "1111111010001011110101",
			2220 => "0000000010001011110101",
			2221 => "1111111010001011110101",
			2222 => "0000001010001011110101",
			2223 => "0000010111011100010000",
			2224 => "0010111010000100001100",
			2225 => "0001000000111100001000",
			2226 => "0001111001010000000100",
			2227 => "0000000010001011110101",
			2228 => "0000000010001011110101",
			2229 => "0000000010001011110101",
			2230 => "1111111010001011110101",
			2231 => "0011100001100000000100",
			2232 => "0000001010001011110101",
			2233 => "0000000010001011110101",
			2234 => "0000000010100100000100",
			2235 => "0000000010001011110101",
			2236 => "0000001010001011110101",
			2237 => "0010001111011000100000",
			2238 => "0000010011110000000100",
			2239 => "1111111010001110010001",
			2240 => "0011110111000000010100",
			2241 => "0011111001110000000100",
			2242 => "1111111010001110010001",
			2243 => "0000111100101100001000",
			2244 => "0011010111011100000100",
			2245 => "0000000010001110010001",
			2246 => "0000001010001110010001",
			2247 => "0010000000110000000100",
			2248 => "1111111010001110010001",
			2249 => "0000000010001110010001",
			2250 => "0011100100000100000100",
			2251 => "1111111010001110010001",
			2252 => "0000000010001110010001",
			2253 => "0000111100110100101100",
			2254 => "0001010011000100011100",
			2255 => "0011000110000000001000",
			2256 => "0010111100101000000100",
			2257 => "0000000010001110010001",
			2258 => "0000001010001110010001",
			2259 => "0000010111011100001100",
			2260 => "0000010011010000001000",
			2261 => "0000011110011000000100",
			2262 => "1111111010001110010001",
			2263 => "0000001010001110010001",
			2264 => "1111111010001110010001",
			2265 => "0010011100110000000100",
			2266 => "0000000010001110010001",
			2267 => "0000001010001110010001",
			2268 => "0011000101101100000100",
			2269 => "0000000010001110010001",
			2270 => "0000001111010000001000",
			2271 => "0000101010101000000100",
			2272 => "0000000010001110010001",
			2273 => "0000001010001110010001",
			2274 => "0000000010001110010001",
			2275 => "1111111010001110010001",
			2276 => "0010001111001000010000",
			2277 => "0000010011110000000100",
			2278 => "1111111010010000100101",
			2279 => "0000111100010000000100",
			2280 => "1111111010010000100101",
			2281 => "0000111000101000000100",
			2282 => "0000000010010000100101",
			2283 => "0000000010010000100101",
			2284 => "0000111000000000001100",
			2285 => "0001101010011000000100",
			2286 => "0000000010010000100101",
			2287 => "0010101100010000000100",
			2288 => "0000001010010000100101",
			2289 => "0000000010010000100101",
			2290 => "0001011001010100001000",
			2291 => "0010110110000000000100",
			2292 => "1111111010010000100101",
			2293 => "0000000010010000100101",
			2294 => "0010101111101000001000",
			2295 => "0001001111011000000100",
			2296 => "0000001010010000100101",
			2297 => "0000000010010000100101",
			2298 => "0001010011000100010000",
			2299 => "0000111000101000001000",
			2300 => "0011110010101000000100",
			2301 => "0000000010010000100101",
			2302 => "0000000010010000100101",
			2303 => "0000010111011100000100",
			2304 => "1111111010010000100101",
			2305 => "0000001010010000100101",
			2306 => "0010101100001100001000",
			2307 => "0010000011001000000100",
			2308 => "0000000010010000100101",
			2309 => "0000001010010000100101",
			2310 => "0010000011100100000100",
			2311 => "1111111010010000100101",
			2312 => "0000000010010000100101",
			2313 => "0010001010000100010000",
			2314 => "0000010011110000000100",
			2315 => "1111111010010010011001",
			2316 => "0000001011001000001000",
			2317 => "0001100110100000000100",
			2318 => "1111111010010010011001",
			2319 => "0000001010010010011001",
			2320 => "1111111010010010011001",
			2321 => "0011111010011000000100",
			2322 => "1111111010010010011001",
			2323 => "0000011001001000100100",
			2324 => "0000110000111000100000",
			2325 => "0001010011000100010000",
			2326 => "0011111100111100001000",
			2327 => "0000011110011000000100",
			2328 => "0000000010010010011001",
			2329 => "0000001010010010011001",
			2330 => "0011001001000100000100",
			2331 => "0000000010010010011001",
			2332 => "1111111010010010011001",
			2333 => "0001110011000100001000",
			2334 => "0010100000111100000100",
			2335 => "0000000010010010011001",
			2336 => "1111111010010010011001",
			2337 => "0000110000111100000100",
			2338 => "0000001010010010011001",
			2339 => "0000000010010010011001",
			2340 => "1111111010010010011001",
			2341 => "0000001010010010011001",
			2342 => "0000010011110000001000",
			2343 => "0010001111011000000100",
			2344 => "1111111010010100110101",
			2345 => "0000000010010100110101",
			2346 => "0000101111001100110100",
			2347 => "0010100000111100100000",
			2348 => "0010001000000000010100",
			2349 => "0000010101010100010000",
			2350 => "0001111011000000001000",
			2351 => "0011111100111000000100",
			2352 => "0000000010010100110101",
			2353 => "0000000010010100110101",
			2354 => "0010011000000100000100",
			2355 => "0000001010010100110101",
			2356 => "0000000010010100110101",
			2357 => "1111111010010100110101",
			2358 => "0001101101010100001000",
			2359 => "0001101100011000000100",
			2360 => "0000000010010100110101",
			2361 => "0000001010010100110101",
			2362 => "0000000010010100110101",
			2363 => "0001011100011100000100",
			2364 => "1111111010010100110101",
			2365 => "0000111010011100001000",
			2366 => "0001001011000000000100",
			2367 => "0000001010010100110101",
			2368 => "0000000010010100110101",
			2369 => "0000010111011100000100",
			2370 => "1111111010010100110101",
			2371 => "0000000010010100110101",
			2372 => "0011100101100000001100",
			2373 => "0011000101111000001000",
			2374 => "0000111111101000000100",
			2375 => "1111111010010100110101",
			2376 => "0000000010010100110101",
			2377 => "0000001010010100110101",
			2378 => "0000101101011000000100",
			2379 => "0000001010010100110101",
			2380 => "0000000010010100110101",
			2381 => "0011010111011100001000",
			2382 => "0010000000110000000100",
			2383 => "1111111010010111011001",
			2384 => "0000000010010111011001",
			2385 => "0010011000000100101000",
			2386 => "0000111000101000010100",
			2387 => "0000101111001100010000",
			2388 => "0010010110000000000100",
			2389 => "1111111010010111011001",
			2390 => "0011111010011000000100",
			2391 => "1111111010010111011001",
			2392 => "0010010011000000000100",
			2393 => "0000000010010111011001",
			2394 => "0000001010010111011001",
			2395 => "1111111010010111011001",
			2396 => "0001111100101100001100",
			2397 => "0011001001001000000100",
			2398 => "1111111010010111011001",
			2399 => "0011000101101100000100",
			2400 => "0000000010010111011001",
			2401 => "0000000010010111011001",
			2402 => "0000010110001100000100",
			2403 => "0000000010010111011001",
			2404 => "0000000010010111011001",
			2405 => "0001010011000100011000",
			2406 => "0001111110001100010100",
			2407 => "0010101111101000001000",
			2408 => "0001110001001000000100",
			2409 => "1111111010010111011001",
			2410 => "0000000010010111011001",
			2411 => "0011101111010100000100",
			2412 => "0000000010010111011001",
			2413 => "0000010111011100000100",
			2414 => "1111111010010111011001",
			2415 => "0000000010010111011001",
			2416 => "0000001010010111011001",
			2417 => "0000110000111000001000",
			2418 => "0010000011001000000100",
			2419 => "0000000010010111011001",
			2420 => "0000001010010111011001",
			2421 => "1111111010010111011001",
			2422 => "0001110011110101010000",
			2423 => "0011110000001100011100",
			2424 => "0001100010110000010000",
			2425 => "0011010111011100000100",
			2426 => "1111111010011010011101",
			2427 => "0011000101011100000100",
			2428 => "0000000010011010011101",
			2429 => "0011111101100000000100",
			2430 => "0000000010011010011101",
			2431 => "0000000010011010011101",
			2432 => "0000011001100000000100",
			2433 => "0000000010011010011101",
			2434 => "0001000110011100000100",
			2435 => "0000001010011010011101",
			2436 => "0000000010011010011101",
			2437 => "0001010001001000100100",
			2438 => "0010000011100100011100",
			2439 => "0001001010000100001100",
			2440 => "0000001011010000000100",
			2441 => "1111111010011010011101",
			2442 => "0011110101100100000100",
			2443 => "0000000010011010011101",
			2444 => "1111111010011010011101",
			2445 => "0010110101010100001000",
			2446 => "0001111100101100000100",
			2447 => "0000000010011010011101",
			2448 => "0000000010011010011101",
			2449 => "0001011011111000000100",
			2450 => "0000000010011010011101",
			2451 => "1111111010011010011101",
			2452 => "0011111001111000000100",
			2453 => "0000000010011010011101",
			2454 => "0000000010011010011101",
			2455 => "0000111011000000001000",
			2456 => "0011011100101000000100",
			2457 => "0000000010011010011101",
			2458 => "0000001010011010011101",
			2459 => "0011001101101000000100",
			2460 => "0000000010011010011101",
			2461 => "0000000010011010011101",
			2462 => "0011000011000000000100",
			2463 => "0000001010011010011101",
			2464 => "0011010011000000001000",
			2465 => "0000111011111000000100",
			2466 => "0000000010011010011101",
			2467 => "0000000010011010011101",
			2468 => "0000000010101100000100",
			2469 => "0000000010011010011101",
			2470 => "0000000010011010011101",
			2471 => "0011011001001000110100",
			2472 => "0011001100101000100100",
			2473 => "0010010011000000011100",
			2474 => "0000100000100100010100",
			2475 => "0001000011000000001100",
			2476 => "0010011001000100000100",
			2477 => "0000000010011110000001",
			2478 => "0000000110000100000100",
			2479 => "0000000010011110000001",
			2480 => "0000000010011110000001",
			2481 => "0000000000100100000100",
			2482 => "0000000010011110000001",
			2483 => "0000000010011110000001",
			2484 => "0001010001001000000100",
			2485 => "0000000010011110000001",
			2486 => "0000000010011110000001",
			2487 => "0001111101001000000100",
			2488 => "0000000010011110000001",
			2489 => "0000000010011110000001",
			2490 => "0001010001001000000100",
			2491 => "0000000010011110000001",
			2492 => "0010100000111100000100",
			2493 => "0000000010011110000001",
			2494 => "0001111000100000000100",
			2495 => "0000000010011110000001",
			2496 => "0000000010011110000001",
			2497 => "0001000011000000011100",
			2498 => "0010000011001000001000",
			2499 => "0001110100101100000100",
			2500 => "0000000010011110000001",
			2501 => "0000000010011110000001",
			2502 => "0010001100110000010000",
			2503 => "0001001100101000001000",
			2504 => "0001000101010100000100",
			2505 => "0000000010011110000001",
			2506 => "0000000010011110000001",
			2507 => "0011101111010100000100",
			2508 => "0000000010011110000001",
			2509 => "0000000010011110000001",
			2510 => "0000000010011110000001",
			2511 => "0010101100001100011100",
			2512 => "0011011010000100001100",
			2513 => "0000001000001100001000",
			2514 => "0001111001011000000100",
			2515 => "0000000010011110000001",
			2516 => "0000000010011110000001",
			2517 => "0000000010011110000001",
			2518 => "0010010110101100001000",
			2519 => "0001010011000100000100",
			2520 => "0000000010011110000001",
			2521 => "0000000010011110000001",
			2522 => "0000001100100100000100",
			2523 => "0000000010011110000001",
			2524 => "0000000010011110000001",
			2525 => "0000111100110100000100",
			2526 => "0000000010011110000001",
			2527 => "0000000010011110000001",
			2528 => "0010000011100101000000",
			2529 => "0000100110010100110000",
			2530 => "0001111100010000000100",
			2531 => "1111111010100001001101",
			2532 => "0010011000000100011000",
			2533 => "0000010011110000001100",
			2534 => "0010101001010100001000",
			2535 => "0000111000000000000100",
			2536 => "0000000010100001001101",
			2537 => "0000000010100001001101",
			2538 => "0000000010100001001101",
			2539 => "0010010011000000001000",
			2540 => "0010101001010100000100",
			2541 => "0000000010100001001101",
			2542 => "0000000010100001001101",
			2543 => "0000001010100001001101",
			2544 => "0010101111101000001000",
			2545 => "0000111100101000000100",
			2546 => "0000000010100001001101",
			2547 => "0000000010100001001101",
			2548 => "0010011000000000000100",
			2549 => "1111111010100001001101",
			2550 => "0010011100010000000100",
			2551 => "0000000010100001001101",
			2552 => "0000000010100001001101",
			2553 => "0010111001001000001100",
			2554 => "0001011000100000000100",
			2555 => "1111111010100001001101",
			2556 => "0010100000111100000100",
			2557 => "0000000010100001001101",
			2558 => "0000000010100001001101",
			2559 => "0000000010100001001101",
			2560 => "0000101111001100011100",
			2561 => "0011000101111000001100",
			2562 => "0001100001100000000100",
			2563 => "0000000010100001001101",
			2564 => "0011100001100000000100",
			2565 => "0000001010100001001101",
			2566 => "0000000010100001001101",
			2567 => "0000010111011100001000",
			2568 => "0001110011110100000100",
			2569 => "1111111010100001001101",
			2570 => "0000000010100001001101",
			2571 => "0000001010101000000100",
			2572 => "0000000010100001001101",
			2573 => "0000000010100001001101",
			2574 => "0000111001010000000100",
			2575 => "0000000010100001001101",
			2576 => "0010101001000000000100",
			2577 => "0000001010100001001101",
			2578 => "0000000010100001001101",
			2579 => "0000010011110000001000",
			2580 => "0010001111011000000100",
			2581 => "1111111010100011011001",
			2582 => "0000000010100011011001",
			2583 => "0001111110001100111000",
			2584 => "0000101111001100101000",
			2585 => "0011000101111000010100",
			2586 => "0010001000000000001100",
			2587 => "0000010101010100001000",
			2588 => "0001010011001000000100",
			2589 => "0000001010100011011001",
			2590 => "0000000010100011011001",
			2591 => "1111111010100011011001",
			2592 => "0011101000101100000100",
			2593 => "0000001010100011011001",
			2594 => "0000000010100011011001",
			2595 => "0000010111011100001100",
			2596 => "0001110011110100001000",
			2597 => "0010011100110000000100",
			2598 => "0000000010100011011001",
			2599 => "1111111010100011011001",
			2600 => "0000000010100011011001",
			2601 => "0011001000000000000100",
			2602 => "0000000010100011011001",
			2603 => "0000000010100011011001",
			2604 => "0011100101100000001100",
			2605 => "0000101001101000001000",
			2606 => "0010101011000000000100",
			2607 => "1111111010100011011001",
			2608 => "0000000010100011011001",
			2609 => "0000000010100011011001",
			2610 => "0000000010100011011001",
			2611 => "0000000011001100000100",
			2612 => "0000000010100011011001",
			2613 => "0000001010100011011001",
			2614 => "0001110011110101000000",
			2615 => "0000010011110000001000",
			2616 => "0010001111011000000100",
			2617 => "1111111010100101111101",
			2618 => "0000000010100101111101",
			2619 => "0001100101100000011000",
			2620 => "0011111011011100010100",
			2621 => "0011110000001100010000",
			2622 => "0011111101100000001000",
			2623 => "0011010101011100000100",
			2624 => "0000000010100101111101",
			2625 => "0000000010100101111101",
			2626 => "0001100010110000000100",
			2627 => "0000000010100101111101",
			2628 => "0000000010100101111101",
			2629 => "0000000010100101111101",
			2630 => "0000000010100101111101",
			2631 => "0001111001011000001000",
			2632 => "0011010101010100000100",
			2633 => "0000000010100101111101",
			2634 => "1111111010100101111101",
			2635 => "0011011001000100001100",
			2636 => "0000001110101000001000",
			2637 => "0011111011110100000100",
			2638 => "0000000010100101111101",
			2639 => "0000001010100101111101",
			2640 => "0000000010100101111101",
			2641 => "0011110101100100001000",
			2642 => "0011111001111000000100",
			2643 => "0000000010100101111101",
			2644 => "1111111010100101111101",
			2645 => "0000000010100101111101",
			2646 => "0011000011000000000100",
			2647 => "0000001010100101111101",
			2648 => "0011010011000000001000",
			2649 => "0000111011111000000100",
			2650 => "0000000010100101111101",
			2651 => "0000000010100101111101",
			2652 => "0000101011111100000100",
			2653 => "0000000010100101111101",
			2654 => "0000000010100101111101",
			2655 => "0010001111001000010000",
			2656 => "0000010011110000000100",
			2657 => "1111111010101000011001",
			2658 => "0010010110000000000100",
			2659 => "0000000010101000011001",
			2660 => "0010011010000100000100",
			2661 => "0000000010101000011001",
			2662 => "0000000010101000011001",
			2663 => "0010101100010000001000",
			2664 => "0001101010011000000100",
			2665 => "0000000010101000011001",
			2666 => "0000001010101000011001",
			2667 => "0010010011000000001100",
			2668 => "0000011101000000001000",
			2669 => "0011010111011100000100",
			2670 => "0000000010101000011001",
			2671 => "0000000010101000011001",
			2672 => "1111111010101000011001",
			2673 => "0001000011000000010000",
			2674 => "0001001101101000001100",
			2675 => "0010101111101000001000",
			2676 => "0001001100101000000100",
			2677 => "0000000010101000011001",
			2678 => "0000001010101000011001",
			2679 => "0000000010101000011001",
			2680 => "1111111010101000011001",
			2681 => "0010100000111100010000",
			2682 => "0011000110000000001000",
			2683 => "0000100101101000000100",
			2684 => "0000001010101000011001",
			2685 => "0000000010101000011001",
			2686 => "0010011000111000000100",
			2687 => "1111111010101000011001",
			2688 => "0000000010101000011001",
			2689 => "0011101110010000001000",
			2690 => "0000010111011100000100",
			2691 => "0000000010101000011001",
			2692 => "0000000010101000011001",
			2693 => "0000001010101000011001",
			2694 => "0011010111011100010100",
			2695 => "0010001111001000000100",
			2696 => "1111111010101010101101",
			2697 => "0001010011001000001000",
			2698 => "0000011001100000000100",
			2699 => "1111111010101010101101",
			2700 => "0000001010101010101101",
			2701 => "0001001000111000000100",
			2702 => "1111111010101010101101",
			2703 => "0000000010101010101101",
			2704 => "0011111010011000000100",
			2705 => "1111111010101010101101",
			2706 => "0000111010011100101100",
			2707 => "0001011000100000011100",
			2708 => "0010101111101000001100",
			2709 => "0010010110000000000100",
			2710 => "1111111010101010101101",
			2711 => "0001100100011100000100",
			2712 => "0000001010101010101101",
			2713 => "0000000010101010101101",
			2714 => "0010000011100100001000",
			2715 => "0000001000010000000100",
			2716 => "0000000010101010101101",
			2717 => "1111111010101010101101",
			2718 => "0000001110101000000100",
			2719 => "0000001010101010101101",
			2720 => "0000000010101010101101",
			2721 => "0010001010000100000100",
			2722 => "1111111010101010101101",
			2723 => "0001110000111100001000",
			2724 => "0000111100101100000100",
			2725 => "0000001010101010101101",
			2726 => "0000000010101010101101",
			2727 => "0000001010101010101101",
			2728 => "0011010011000000000100",
			2729 => "1111111010101010101101",
			2730 => "0000000010101010101101",
			2731 => "0010001111011000100000",
			2732 => "0000010011110000000100",
			2733 => "1111111010101101000001",
			2734 => "0011111001110000000100",
			2735 => "1111111010101101000001",
			2736 => "0011110111010000010000",
			2737 => "0011000111011100000100",
			2738 => "0000000010101101000001",
			2739 => "0000111100101100000100",
			2740 => "0000001010101101000001",
			2741 => "0010000000110000000100",
			2742 => "1111111010101101000001",
			2743 => "0000000010101101000001",
			2744 => "0001101011110100000100",
			2745 => "1111111010101101000001",
			2746 => "0000000010101101000001",
			2747 => "0011110000110100000100",
			2748 => "1111111010101101000001",
			2749 => "0000110000111000100100",
			2750 => "0001010011000100010100",
			2751 => "0000111000000000000100",
			2752 => "0000001010101101000001",
			2753 => "0000100100010100001000",
			2754 => "0010001000000000000100",
			2755 => "0000000010101101000001",
			2756 => "0000001010101101000001",
			2757 => "0000111001010000000100",
			2758 => "1111111010101101000001",
			2759 => "0000000010101101000001",
			2760 => "0001110000111100001000",
			2761 => "0010011100000000000100",
			2762 => "0000000010101101000001",
			2763 => "0000001010101101000001",
			2764 => "0011000110000000000100",
			2765 => "0000001010101101000001",
			2766 => "0000001010101101000001",
			2767 => "1111111010101101000001",
			2768 => "0011100010110101001000",
			2769 => "0000001010010100111100",
			2770 => "0011100110111000110100",
			2771 => "0000011110011000100000",
			2772 => "0001000011000000010000",
			2773 => "0001001001000100001000",
			2774 => "0000011101000000000100",
			2775 => "0000000010110000011101",
			2776 => "0000000010110000011101",
			2777 => "0000010011110000000100",
			2778 => "0000000010110000011101",
			2779 => "0000000010110000011101",
			2780 => "0000111001010100001000",
			2781 => "0001011011111000000100",
			2782 => "0000000010110000011101",
			2783 => "0000000010110000011101",
			2784 => "0010001111011000000100",
			2785 => "0000000010110000011101",
			2786 => "0000000010110000011101",
			2787 => "0000101100010100010000",
			2788 => "0010101011111000001000",
			2789 => "0011011101101000000100",
			2790 => "0000000010110000011101",
			2791 => "0000000010110000011101",
			2792 => "0011111010011000000100",
			2793 => "0000000010110000011101",
			2794 => "0000000010110000011101",
			2795 => "0000001010110000011101",
			2796 => "0001010011000100000100",
			2797 => "0000000010110000011101",
			2798 => "0000000010110000011101",
			2799 => "0010011100000000001000",
			2800 => "0001001100010000000100",
			2801 => "1111111010110000011101",
			2802 => "0000000010110000011101",
			2803 => "0000000010110000011101",
			2804 => "0000111001010000011000",
			2805 => "0010101000101000001000",
			2806 => "0001000101010100000100",
			2807 => "0000000010110000011101",
			2808 => "0000000010110000011101",
			2809 => "0000101101111000001000",
			2810 => "0000010110001100000100",
			2811 => "0000000010110000011101",
			2812 => "0000000010110000011101",
			2813 => "0011111110011100000100",
			2814 => "1111111010110000011101",
			2815 => "0000000010110000011101",
			2816 => "0010100000111100001000",
			2817 => "0010110101010100000100",
			2818 => "0000000010110000011101",
			2819 => "0000001010110000011101",
			2820 => "0001001101001000000100",
			2821 => "0000000010110000011101",
			2822 => "0000000010110000011101",
			2823 => "0011010101011100100000",
			2824 => "0001111100110000000100",
			2825 => "0000000010110011001001",
			2826 => "0000100101011000010000",
			2827 => "0010111110011000000100",
			2828 => "0000000010110011001001",
			2829 => "0001011000100000001000",
			2830 => "0000011001100000000100",
			2831 => "0000000010110011001001",
			2832 => "0000000010110011001001",
			2833 => "0000000010110011001001",
			2834 => "0000111011111000000100",
			2835 => "0000000010110011001001",
			2836 => "0011001100101000000100",
			2837 => "0000000010110011001001",
			2838 => "0000000010110011001001",
			2839 => "0000111100110100110100",
			2840 => "0001011000100000101100",
			2841 => "0000011110011000010000",
			2842 => "0010101011111000001100",
			2843 => "0010110101101100001000",
			2844 => "0010001010000100000100",
			2845 => "0000000010110011001001",
			2846 => "0000000010110011001001",
			2847 => "0000000010110011001001",
			2848 => "0000000010110011001001",
			2849 => "0001000011000000010000",
			2850 => "0001001001000100001000",
			2851 => "0011001100000000000100",
			2852 => "0000000010110011001001",
			2853 => "0000000010110011001001",
			2854 => "0011100011101000000100",
			2855 => "0000000010110011001001",
			2856 => "0000000010110011001001",
			2857 => "0000101111001100001000",
			2858 => "0010100100101100000100",
			2859 => "0000000010110011001001",
			2860 => "0000001010110011001001",
			2861 => "0000000010110011001001",
			2862 => "0000010110001100000100",
			2863 => "0000000010110011001001",
			2864 => "0000001010110011001001",
			2865 => "0000000010110011001001",
			2866 => "0011011101101001100100",
			2867 => "0001011100101100111000",
			2868 => "0000001101001100010100",
			2869 => "0000100100001000001100",
			2870 => "0011010111011100000100",
			2871 => "0000000010110111010101",
			2872 => "0011101100001100000100",
			2873 => "0000000010110111010101",
			2874 => "0000000010110111010101",
			2875 => "0010110111011100000100",
			2876 => "0000001010110111010101",
			2877 => "0000000010110111010101",
			2878 => "0011100010110100010000",
			2879 => "0000101111101100001100",
			2880 => "0000001100100100001000",
			2881 => "0000111100010000000100",
			2882 => "0000000010110111010101",
			2883 => "0000000010110111010101",
			2884 => "0000000010110111010101",
			2885 => "1111111010110111010101",
			2886 => "0010101000101000001000",
			2887 => "0011110111001100000100",
			2888 => "0000000010110111010101",
			2889 => "0000000010110111010101",
			2890 => "0000101101111000001000",
			2891 => "0000001100100100000100",
			2892 => "0000000010110111010101",
			2893 => "0000000010110111010101",
			2894 => "1111111010110111010101",
			2895 => "0011011001001000011100",
			2896 => "0011001001001000010000",
			2897 => "0001111011111000001100",
			2898 => "0000111001010000001000",
			2899 => "0001111100110000000100",
			2900 => "0000000010110111010101",
			2901 => "0000000010110111010101",
			2902 => "0000000010110111010101",
			2903 => "0000000010110111010101",
			2904 => "0011001001000100000100",
			2905 => "1111111010110111010101",
			2906 => "0011000110000000000100",
			2907 => "0000000010110111010101",
			2908 => "0000000010110111010101",
			2909 => "0000001110101000001100",
			2910 => "0000111110001100001000",
			2911 => "0001110110011100000100",
			2912 => "0000000010110111010101",
			2913 => "0000001010110111010101",
			2914 => "0000000010110111010101",
			2915 => "0000000010110111010101",
			2916 => "0001000110101100010000",
			2917 => "0010001001010100001000",
			2918 => "0000000001110100000100",
			2919 => "0000000010110111010101",
			2920 => "0000001010110111010101",
			2921 => "0001010110011100000100",
			2922 => "0000000010110111010101",
			2923 => "0000000010110111010101",
			2924 => "0011011010000100000100",
			2925 => "0000000010110111010101",
			2926 => "0000010111011100001000",
			2927 => "0010001000000000000100",
			2928 => "0000000010110111010101",
			2929 => "1111111010110111010101",
			2930 => "0000000010100100000100",
			2931 => "0000000010110111010101",
			2932 => "0000000010110111010101",
			2933 => "0010001000000001010000",
			2934 => "0011111100111100111000",
			2935 => "0001101010101100110100",
			2936 => "0000111001010100011100",
			2937 => "0010010110000000001100",
			2938 => "0001010101111000001000",
			2939 => "0010101000000000000100",
			2940 => "0000000010111010111001",
			2941 => "0000000010111010111001",
			2942 => "0000000010111010111001",
			2943 => "0010011000000100001000",
			2944 => "0001101010011000000100",
			2945 => "0000000010111010111001",
			2946 => "0000000010111010111001",
			2947 => "0011011001000100000100",
			2948 => "0000000010111010111001",
			2949 => "0000000010111010111001",
			2950 => "0001001100000000001100",
			2951 => "0011110010111100001000",
			2952 => "0011011100101000000100",
			2953 => "0000000010111010111001",
			2954 => "0000000010111010111001",
			2955 => "0000000010111010111001",
			2956 => "0010000011100100001000",
			2957 => "0001110001001000000100",
			2958 => "0000000010111010111001",
			2959 => "0000000010111010111001",
			2960 => "0000000010111010111001",
			2961 => "0000000010111010111001",
			2962 => "0010101011000000001100",
			2963 => "0001001001001000001000",
			2964 => "0001001100101000000100",
			2965 => "0000000010111010111001",
			2966 => "0000000010111010111001",
			2967 => "0000000010111010111001",
			2968 => "0001110000111100001000",
			2969 => "0000111111101000000100",
			2970 => "0000000010111010111001",
			2971 => "0000000010111010111001",
			2972 => "0000000010111010111001",
			2973 => "0011100110110000001100",
			2974 => "0010101111101000000100",
			2975 => "0000000010111010111001",
			2976 => "0001101010001000000100",
			2977 => "0000000010111010111001",
			2978 => "0000000010111010111001",
			2979 => "0000101111001100001000",
			2980 => "0001101101010100000100",
			2981 => "0000000010111010111001",
			2982 => "0000000010111010111001",
			2983 => "0000101110110000000100",
			2984 => "0000000010111010111001",
			2985 => "0001100110011000000100",
			2986 => "0000000010111010111001",
			2987 => "0011110011100000000100",
			2988 => "0000000010111010111001",
			2989 => "0000000010111010111001",
			2990 => "0001110011110101011100",
			2991 => "0001010001001001000000",
			2992 => "0010101111101000100000",
			2993 => "0001001010000100010000",
			2994 => "0010010110000000000100",
			2995 => "0000000010111101111101",
			2996 => "0001000101010100000100",
			2997 => "0000000010111101111101",
			2998 => "0001101111000100000100",
			2999 => "0000000010111101111101",
			3000 => "0000000010111101111101",
			3001 => "0001111101001000001000",
			3002 => "0010011001000100000100",
			3003 => "0000000010111101111101",
			3004 => "0000000010111101111101",
			3005 => "0001001111011000000100",
			3006 => "0000000010111101111101",
			3007 => "0000000010111101111101",
			3008 => "0000101100001000010000",
			3009 => "0001010100101100000100",
			3010 => "0000000010111101111101",
			3011 => "0000111000101000000100",
			3012 => "0000000010111101111101",
			3013 => "0011010101011100000100",
			3014 => "0000000010111101111101",
			3015 => "0000000010111101111101",
			3016 => "0010000011100100001100",
			3017 => "0010110101010100001000",
			3018 => "0001010110011100000100",
			3019 => "0000000010111101111101",
			3020 => "0000000010111101111101",
			3021 => "0000000010111101111101",
			3022 => "0000000010111101111101",
			3023 => "0000111011000000001000",
			3024 => "0010001010000100000100",
			3025 => "0000000010111101111101",
			3026 => "0000000010111101111101",
			3027 => "0000010011010000001100",
			3028 => "0001111110111000001000",
			3029 => "0010101000100000000100",
			3030 => "0000000010111101111101",
			3031 => "0000000010111101111101",
			3032 => "0000000010111101111101",
			3033 => "0000110001001000000100",
			3034 => "0000000010111101111101",
			3035 => "0000000010111101111101",
			3036 => "0001100101100000000100",
			3037 => "0000000010111101111101",
			3038 => "0000000010111101111101",
			3039 => "0001110011110101001100",
			3040 => "0011110000001100100000",
			3041 => "0001111100010000000100",
			3042 => "0000000011000000111001",
			3043 => "0011011010100100000100",
			3044 => "0000000011000000111001",
			3045 => "0001000110011100010000",
			3046 => "0001000110000000001000",
			3047 => "0000001101001100000100",
			3048 => "0000000011000000111001",
			3049 => "0000000011000000111001",
			3050 => "0001101010001100000100",
			3051 => "0000000011000000111001",
			3052 => "0000001011000000111001",
			3053 => "0001101101100100000100",
			3054 => "0000000011000000111001",
			3055 => "0000000011000000111001",
			3056 => "0001111011111000000100",
			3057 => "1111111011000000111001",
			3058 => "0001000011000000010000",
			3059 => "0001001010000100001100",
			3060 => "0010101111101000001000",
			3061 => "0001000101010100000100",
			3062 => "0000000011000000111001",
			3063 => "0000001011000000111001",
			3064 => "0000000011000000111001",
			3065 => "1111111011000000111001",
			3066 => "0001001100000000001000",
			3067 => "0000101111001100000100",
			3068 => "0000001011000000111001",
			3069 => "0000000011000000111001",
			3070 => "0010000011100100001000",
			3071 => "0001011000100000000100",
			3072 => "1111111011000000111001",
			3073 => "0000000011000000111001",
			3074 => "0011011010000100000100",
			3075 => "0000001011000000111001",
			3076 => "0000000011000000111001",
			3077 => "0011000011000000000100",
			3078 => "0000001011000000111001",
			3079 => "0011010011000000001000",
			3080 => "0001011010011100000100",
			3081 => "0000000011000000111001",
			3082 => "0000000011000000111001",
			3083 => "0000101011111100000100",
			3084 => "0000000011000000111001",
			3085 => "0000000011000000111001",
			3086 => "0010001111011000101000",
			3087 => "0000111011111000100000",
			3088 => "0001100001000000011100",
			3089 => "0001100010110000010100",
			3090 => "0001010110011100001100",
			3091 => "0000100001000000001000",
			3092 => "0000000111100000000100",
			3093 => "0000000011000100011101",
			3094 => "0000000011000100011101",
			3095 => "0000000011000100011101",
			3096 => "0000001100111000000100",
			3097 => "0000000011000100011101",
			3098 => "0000000011000100011101",
			3099 => "0000110011001000000100",
			3100 => "0000000011000100011101",
			3101 => "0000000011000100011101",
			3102 => "0000000011000100011101",
			3103 => "0010101001011000000100",
			3104 => "0000000011000100011101",
			3105 => "0000000011000100011101",
			3106 => "0000101111001100111100",
			3107 => "0000111111101000100100",
			3108 => "0000000100010100010100",
			3109 => "0010011000000100001000",
			3110 => "0011111010011000000100",
			3111 => "0000000011000100011101",
			3112 => "0000000011000100011101",
			3113 => "0010001000000000000100",
			3114 => "0000000011000100011101",
			3115 => "0011100001001100000100",
			3116 => "0000000011000100011101",
			3117 => "0000000011000100011101",
			3118 => "0011000110000000000100",
			3119 => "0000000011000100011101",
			3120 => "0001101010110000000100",
			3121 => "0000000011000100011101",
			3122 => "0001100101111100000100",
			3123 => "0000000011000100011101",
			3124 => "0000000011000100011101",
			3125 => "0001010011000100000100",
			3126 => "0000000011000100011101",
			3127 => "0001101010111100001100",
			3128 => "0001111011000000000100",
			3129 => "0000000011000100011101",
			3130 => "0000011010100100000100",
			3131 => "0000000011000100011101",
			3132 => "0000000011000100011101",
			3133 => "0001001011000000000100",
			3134 => "0000000011000100011101",
			3135 => "0000000011000100011101",
			3136 => "0010110011000000001100",
			3137 => "0000111001010000000100",
			3138 => "0000000011000100011101",
			3139 => "0001100101111100000100",
			3140 => "0000000011000100011101",
			3141 => "0000000011000100011101",
			3142 => "0000000011000100011101",
			3143 => "0001110011110101010000",
			3144 => "0000010011110000001000",
			3145 => "0010001111011000000100",
			3146 => "1111111011000111100001",
			3147 => "0000000011000111100001",
			3148 => "0011110000001100100000",
			3149 => "0001100010110000011100",
			3150 => "0011010101011100010000",
			3151 => "0010001001000100001000",
			3152 => "0010000101101100000100",
			3153 => "0000000011000111100001",
			3154 => "0000000011000111100001",
			3155 => "0000111101101000000100",
			3156 => "0000000011000111100001",
			3157 => "1111111011000111100001",
			3158 => "0001101010001100000100",
			3159 => "0000000011000111100001",
			3160 => "0000100101100100000100",
			3161 => "0000001011000111100001",
			3162 => "0000000011000111100001",
			3163 => "0000001011000111100001",
			3164 => "0001010011000100011000",
			3165 => "0001001010000100001100",
			3166 => "0010101111101000001000",
			3167 => "0001011000111000000100",
			3168 => "0000000011000111100001",
			3169 => "0000001011000111100001",
			3170 => "0000000011000111100001",
			3171 => "0010000011100100001000",
			3172 => "0010110101010100000100",
			3173 => "0000000011000111100001",
			3174 => "1111111011000111100001",
			3175 => "0000000011000111100001",
			3176 => "0000111011000000001000",
			3177 => "0010000011001000000100",
			3178 => "0000000011000111100001",
			3179 => "0000001011000111100001",
			3180 => "0011100111100000000100",
			3181 => "0000000011000111100001",
			3182 => "0000000011000111100001",
			3183 => "0011000011000000000100",
			3184 => "0000001011000111100001",
			3185 => "0011010011000000001000",
			3186 => "0000111011111000000100",
			3187 => "0000000011000111100001",
			3188 => "0000000011000111100001",
			3189 => "0000000010101100000100",
			3190 => "0000000011000111100001",
			3191 => "0000000011000111100001",
			3192 => "0011010111011100001000",
			3193 => "0010000000110000000100",
			3194 => "1111111011001001111101",
			3195 => "0000000011001001111101",
			3196 => "0000111100110101000100",
			3197 => "0001011000100000101100",
			3198 => "0000101111101100010000",
			3199 => "0011111010011000000100",
			3200 => "1111111011001001111101",
			3201 => "0011100110111000001000",
			3202 => "0011010101101100000100",
			3203 => "0000000011001001111101",
			3204 => "0000001011001001111101",
			3205 => "0000000011001001111101",
			3206 => "0010000011100100010000",
			3207 => "0000001001101000001000",
			3208 => "0000111001010100000100",
			3209 => "1111111011001001111101",
			3210 => "1111111011001001111101",
			3211 => "0000010110001100000100",
			3212 => "1111111011001001111101",
			3213 => "0000000011001001111101",
			3214 => "0001011011111000000100",
			3215 => "0000001011001001111101",
			3216 => "0000111001010000000100",
			3217 => "1111111011001001111101",
			3218 => "0000000011001001111101",
			3219 => "0011110000000100001100",
			3220 => "0010000011001000001000",
			3221 => "0000110011000100000100",
			3222 => "0000000011001001111101",
			3223 => "1111111011001001111101",
			3224 => "0000001011001001111101",
			3225 => "0000000101010000000100",
			3226 => "0000001011001001111101",
			3227 => "0011110100110100000100",
			3228 => "0000000011001001111101",
			3229 => "0000001011001001111101",
			3230 => "1111111011001001111101",
			3231 => "0001111100011101010100",
			3232 => "0000101111001101001100",
			3233 => "0000111000101000101000",
			3234 => "0000111100110000010100",
			3235 => "0000010011010000010000",
			3236 => "0011000111011100001000",
			3237 => "0001010011001000000100",
			3238 => "0000000011001101001001",
			3239 => "0000000011001101001001",
			3240 => "0001101010011000000100",
			3241 => "0000000011001101001001",
			3242 => "0000000011001101001001",
			3243 => "0000000011001101001001",
			3244 => "0001111011000000010000",
			3245 => "0001100100010000001000",
			3246 => "0000100111100000000100",
			3247 => "0000000011001101001001",
			3248 => "0000000011001101001001",
			3249 => "0001001010000100000100",
			3250 => "0000000011001101001001",
			3251 => "0000000011001101001001",
			3252 => "0000000011001101001001",
			3253 => "0010000011001000010100",
			3254 => "0010110111011100001000",
			3255 => "0000100010100100000100",
			3256 => "0000000011001101001001",
			3257 => "0000000011001101001001",
			3258 => "0011010101101100000100",
			3259 => "0000000011001101001001",
			3260 => "0011011001000100000100",
			3261 => "0000000011001101001001",
			3262 => "0000000011001101001001",
			3263 => "0001111001000000001100",
			3264 => "0000111100110100001000",
			3265 => "0011100011011000000100",
			3266 => "0000000011001101001001",
			3267 => "0000000011001101001001",
			3268 => "0000000011001101001001",
			3269 => "0000000011001101001001",
			3270 => "0000000010100000000100",
			3271 => "0000000011001101001001",
			3272 => "0000000011001101001001",
			3273 => "0000111010100000010000",
			3274 => "0000011100101000000100",
			3275 => "0000000011001101001001",
			3276 => "0011101000110100001000",
			3277 => "0000011001000100000100",
			3278 => "0000000011001101001001",
			3279 => "0000000011001101001001",
			3280 => "0000000011001101001001",
			3281 => "0000000011001101001001",
			3282 => "0000010011110000001000",
			3283 => "0010001111011000000100",
			3284 => "1111111011001111100111",
			3285 => "0000000011001111100111",
			3286 => "0010010110000000000100",
			3287 => "1111111011001111100111",
			3288 => "0000101000010000100100",
			3289 => "0011111010011000000100",
			3290 => "1111111011001111100111",
			3291 => "0010101001011000010000",
			3292 => "0010011000000100001000",
			3293 => "0001001111011000000100",
			3294 => "0000001011001111100111",
			3295 => "0000001011001111100111",
			3296 => "0000000100010100000100",
			3297 => "0000000011001111100111",
			3298 => "0000001011001111100111",
			3299 => "0010000011001000001000",
			3300 => "0001110001011000000100",
			3301 => "1111111011001111100111",
			3302 => "0000000011001111100111",
			3303 => "0011100011011000000100",
			3304 => "0000000011001111100111",
			3305 => "0000001011001111100111",
			3306 => "0001111100011100010100",
			3307 => "0010000011100100001100",
			3308 => "0000111001010100000100",
			3309 => "1111111011001111100111",
			3310 => "0011011001001000000100",
			3311 => "1111111011001111100111",
			3312 => "0000000011001111100111",
			3313 => "0010101000100000000100",
			3314 => "0000000011001111100111",
			3315 => "0000000011001111100111",
			3316 => "0000111001010000001000",
			3317 => "0001111100110100000100",
			3318 => "0000000011001111100111",
			3319 => "0000001011001111100111",
			3320 => "0000001011001111100111",
			3321 => "0000010110001100011100",
			3322 => "0010000000110000010000",
			3323 => "0000010011110000000100",
			3324 => "1111111011010001011001",
			3325 => "0010110111011100001000",
			3326 => "0010011001000100000100",
			3327 => "1111111011010001011001",
			3328 => "0000001011010001011001",
			3329 => "1111111011010001011001",
			3330 => "0010111001001000001000",
			3331 => "0011111101010100000100",
			3332 => "0000001011010001011001",
			3333 => "0000000011010001011001",
			3334 => "1111111011010001011001",
			3335 => "0011111010011000000100",
			3336 => "1111111011010001011001",
			3337 => "0010101110010100011000",
			3338 => "0011010101011100000100",
			3339 => "0000000011010001011001",
			3340 => "0001011000100000001100",
			3341 => "0000000110101000000100",
			3342 => "0000001011010001011001",
			3343 => "0001110011110100000100",
			3344 => "0000000011010001011001",
			3345 => "0000001011010001011001",
			3346 => "0011000101101100000100",
			3347 => "0000001011010001011001",
			3348 => "0000001011010001011001",
			3349 => "1111111011010001011001",
			3350 => "0010000011001000101000",
			3351 => "0010101001010100010000",
			3352 => "0010011001000100000100",
			3353 => "0000000011010100010101",
			3354 => "0011111100111000001000",
			3355 => "0001101010011000000100",
			3356 => "0000000011010100010101",
			3357 => "0000000011010100010101",
			3358 => "0000000011010100010101",
			3359 => "0011100110000100001100",
			3360 => "0010111010100100001000",
			3361 => "0000111100110000000100",
			3362 => "0000000011010100010101",
			3363 => "0000000011010100010101",
			3364 => "0000000011010100010101",
			3365 => "0000101010010100000100",
			3366 => "0000000011010100010101",
			3367 => "0011010101010100000100",
			3368 => "0000000011010100010101",
			3369 => "0000000011010100010101",
			3370 => "0000111001010000010100",
			3371 => "0000111000000000001000",
			3372 => "0000001110111100000100",
			3373 => "0000000011010100010101",
			3374 => "0000000011010100010101",
			3375 => "0000100110010100000100",
			3376 => "0000000011010100010101",
			3377 => "0001111110001100000100",
			3378 => "0000000011010100010101",
			3379 => "0000000011010100010101",
			3380 => "0010101110111000010100",
			3381 => "0000001000010000001000",
			3382 => "0000000110101000000100",
			3383 => "0000000011010100010101",
			3384 => "0000000011010100010101",
			3385 => "0011000101111000000100",
			3386 => "0000000011010100010101",
			3387 => "0011010101111000000100",
			3388 => "0000000011010100010101",
			3389 => "0000000011010100010101",
			3390 => "0000010111011100001000",
			3391 => "0001110011110100000100",
			3392 => "0000000011010100010101",
			3393 => "0000000011010100010101",
			3394 => "0000000010100100000100",
			3395 => "0000000011010100010101",
			3396 => "0000000011010100010101",
			3397 => "0000011110011000110100",
			3398 => "0000010110001100100100",
			3399 => "0000010011110000001000",
			3400 => "0010001111011000000100",
			3401 => "1111111011010110111001",
			3402 => "1111111011010110111001",
			3403 => "0011110100010000001100",
			3404 => "0011000101011100001000",
			3405 => "0001011100110000000100",
			3406 => "1111111011010110111001",
			3407 => "0000000011010110111001",
			3408 => "1111111011010110111001",
			3409 => "0010000000110000001000",
			3410 => "0000001011111100000100",
			3411 => "0000000011010110111001",
			3412 => "1111111011010110111001",
			3413 => "0011110110011000000100",
			3414 => "0000010011010110111001",
			3415 => "0000000011010110111001",
			3416 => "0011111101100000001000",
			3417 => "0001101010011000000100",
			3418 => "1111111011010110111001",
			3419 => "0000000011010110111001",
			3420 => "0001010011000100000100",
			3421 => "0000000011010110111001",
			3422 => "0000010011010110111001",
			3423 => "0011110011101000001000",
			3424 => "0011000011001000000100",
			3425 => "0000000011010110111001",
			3426 => "1111111011010110111001",
			3427 => "0010010011001000000100",
			3428 => "0000001011010110111001",
			3429 => "0000111100110000001000",
			3430 => "0001111110111000000100",
			3431 => "0000001011010110111001",
			3432 => "0000010011010110111001",
			3433 => "0011110110011000000100",
			3434 => "0000010011010110111001",
			3435 => "0011111011110100000100",
			3436 => "0000010011010110111001",
			3437 => "0000010011010110111001",
			3438 => "0011010101011100010000",
			3439 => "0001010101111000001000",
			3440 => "0010101000000000000100",
			3441 => "0000000011011001011101",
			3442 => "0000000011011001011101",
			3443 => "0011100101001100000100",
			3444 => "0000000011011001011101",
			3445 => "0000000011011001011101",
			3446 => "0010011000000100011100",
			3447 => "0001001010000100001100",
			3448 => "0010110101101100001000",
			3449 => "0001000101010100000100",
			3450 => "0000000011011001011101",
			3451 => "0000000011011001011101",
			3452 => "0000000011011001011101",
			3453 => "0001001000000100001000",
			3454 => "0011110110011000000100",
			3455 => "0000000011011001011101",
			3456 => "0000000011011001011101",
			3457 => "0001101110001000000100",
			3458 => "0000000011011001011101",
			3459 => "0000000011011001011101",
			3460 => "0001010011000100011100",
			3461 => "0010010110101100010100",
			3462 => "0001011011111000001100",
			3463 => "0000111100010000001000",
			3464 => "0001001100101000000100",
			3465 => "0000000011011001011101",
			3466 => "0000000011011001011101",
			3467 => "0000000011011001011101",
			3468 => "0000010101011100000100",
			3469 => "0000000011011001011101",
			3470 => "0000000011011001011101",
			3471 => "0000001100100100000100",
			3472 => "0000000011011001011101",
			3473 => "0000000011011001011101",
			3474 => "0000110000111000001000",
			3475 => "0001011000100000000100",
			3476 => "0000000011011001011101",
			3477 => "0000000011011001011101",
			3478 => "0000000011011001011101",
			3479 => "0011110000001000100100",
			3480 => "0011111001110000001100",
			3481 => "0000000111101000000100",
			3482 => "0000000011011100100001",
			3483 => "0000000001111000000100",
			3484 => "0000000011011100100001",
			3485 => "0000000011011100100001",
			3486 => "0010010110000000001000",
			3487 => "0000000000000100000100",
			3488 => "0000000011011100100001",
			3489 => "0000000011011100100001",
			3490 => "0011010111011100001000",
			3491 => "0010011111011000000100",
			3492 => "0000000011011100100001",
			3493 => "0000000011011100100001",
			3494 => "0001011010100000000100",
			3495 => "0000000011011100100001",
			3496 => "0000000011011100100001",
			3497 => "0011100010110100010100",
			3498 => "0001110001001000001100",
			3499 => "0010110101010100001000",
			3500 => "0010110111011100000100",
			3501 => "0000000011011100100001",
			3502 => "0000000011011100100001",
			3503 => "0000000011011100100001",
			3504 => "0001011000100000000100",
			3505 => "0000000011011100100001",
			3506 => "0000000011011100100001",
			3507 => "0000111001010000010100",
			3508 => "0010101000101000001000",
			3509 => "0001000101010100000100",
			3510 => "0000000011011100100001",
			3511 => "0000000011011100100001",
			3512 => "0000101101111000001000",
			3513 => "0000010110001100000100",
			3514 => "0000000011011100100001",
			3515 => "0000000011011100100001",
			3516 => "0000000011011100100001",
			3517 => "0010100000111100001100",
			3518 => "0011011001001000001000",
			3519 => "0000000101101000000100",
			3520 => "0000000011011100100001",
			3521 => "0000000011011100100001",
			3522 => "0000000011011100100001",
			3523 => "0001001101001000000100",
			3524 => "0000000011011100100001",
			3525 => "0000001010010000000100",
			3526 => "0000000011011100100001",
			3527 => "0000000011011100100001",
			3528 => "0000010110001100100100",
			3529 => "0010000000110000010100",
			3530 => "0000010011110000000100",
			3531 => "1111111011011110101101",
			3532 => "0010111010100100001000",
			3533 => "0011011010100100000100",
			3534 => "1111111011011110101101",
			3535 => "0000001011011110101101",
			3536 => "0010110111011100000100",
			3537 => "0000000011011110101101",
			3538 => "1111111011011110101101",
			3539 => "0011001001000100001100",
			3540 => "0001111101001000000100",
			3541 => "1111111011011110101101",
			3542 => "0011110100011000000100",
			3543 => "0000001011011110101101",
			3544 => "0000000011011110101101",
			3545 => "1111111011011110101101",
			3546 => "0001101010001100000100",
			3547 => "1111111011011110101101",
			3548 => "0000110000111000011100",
			3549 => "0011010101011100000100",
			3550 => "0000000011011110101101",
			3551 => "0000101111001100001100",
			3552 => "0011100100001100000100",
			3553 => "0000001011011110101101",
			3554 => "0001111001011000000100",
			3555 => "0000000011011110101101",
			3556 => "0000001011011110101101",
			3557 => "0011101110010000000100",
			3558 => "1111111011011110101101",
			3559 => "0000111001010000000100",
			3560 => "0000000011011110101101",
			3561 => "0000001011011110101101",
			3562 => "1111111011011110101101",
			3563 => "0010010011000000011100",
			3564 => "0000100000100100010000",
			3565 => "0000100000001100000100",
			3566 => "0000000011100001011001",
			3567 => "0011101111111000000100",
			3568 => "0000000011100001011001",
			3569 => "0000110011001000000100",
			3570 => "0000000011100001011001",
			3571 => "0000000011100001011001",
			3572 => "0001010001001000000100",
			3573 => "0000000011100001011001",
			3574 => "0001011110111000000100",
			3575 => "0000000011100001011001",
			3576 => "0000000011100001011001",
			3577 => "0001000011000000010000",
			3578 => "0001001010000100001100",
			3579 => "0010101111101000001000",
			3580 => "0001011000111000000100",
			3581 => "0000000011100001011001",
			3582 => "0000000011100001011001",
			3583 => "0000000011100001011001",
			3584 => "0000000011100001011001",
			3585 => "0010100000111100011000",
			3586 => "0000101111001100010000",
			3587 => "0010001111011000000100",
			3588 => "0000000011100001011001",
			3589 => "0011010110000000000100",
			3590 => "0000000011100001011001",
			3591 => "0010111101101000000100",
			3592 => "0000000011100001011001",
			3593 => "0000000011100001011001",
			3594 => "0000111001010000000100",
			3595 => "0000000011100001011001",
			3596 => "0000000011100001011001",
			3597 => "0001101110000100010000",
			3598 => "0000000101101000001100",
			3599 => "0011011001001000000100",
			3600 => "0000000011100001011001",
			3601 => "0001001110111000000100",
			3602 => "0000000011100001011001",
			3603 => "0000000011100001011001",
			3604 => "0000000011100001011001",
			3605 => "0000000011100001011001",
			3606 => "0011010111011100010100",
			3607 => "0010001111001000000100",
			3608 => "1111111011100011100101",
			3609 => "0001010011001000001000",
			3610 => "0011101000101000000100",
			3611 => "0000000011100011100101",
			3612 => "0000001011100011100101",
			3613 => "0001001000111000000100",
			3614 => "1111111011100011100101",
			3615 => "0000000011100011100101",
			3616 => "0000111100110100110000",
			3617 => "0001011000100000010100",
			3618 => "0001001100010000010000",
			3619 => "0001111010011100001100",
			3620 => "0011100101000000001000",
			3621 => "0011100010110100000100",
			3622 => "0000000011100011100101",
			3623 => "0000001011100011100101",
			3624 => "1111111011100011100101",
			3625 => "0000001011100011100101",
			3626 => "1111111011100011100101",
			3627 => "0011110000000100001100",
			3628 => "0010000011001000001000",
			3629 => "0010111100101000000100",
			3630 => "0000000011100011100101",
			3631 => "1111111011100011100101",
			3632 => "0000001011100011100101",
			3633 => "0000100101101000001000",
			3634 => "0000001110110000000100",
			3635 => "0000001011100011100101",
			3636 => "0000001011100011100101",
			3637 => "0011100101100000000100",
			3638 => "0000000011100011100101",
			3639 => "0000001011100011100101",
			3640 => "1111111011100011100101",
			3641 => "0011010111011100010100",
			3642 => "0010001111001000000100",
			3643 => "1111111011100101111001",
			3644 => "0001010011001000001000",
			3645 => "0001111000111000000100",
			3646 => "0000000011100101111001",
			3647 => "0000001011100101111001",
			3648 => "0011000101011100000100",
			3649 => "1111111011100101111001",
			3650 => "0000000011100101111001",
			3651 => "0001111100011100101000",
			3652 => "0011111010011000000100",
			3653 => "1111111011100101111001",
			3654 => "0000000100110100001000",
			3655 => "0001000001011000000100",
			3656 => "0000001011100101111001",
			3657 => "1111111011100101111001",
			3658 => "0010000011100100010000",
			3659 => "0001001010000100001000",
			3660 => "0000111100010000000100",
			3661 => "0000000011100101111001",
			3662 => "0000001011100101111001",
			3663 => "0001101101010000000100",
			3664 => "0000000011100101111001",
			3665 => "1111111011100101111001",
			3666 => "0001000011000000000100",
			3667 => "0000000011100101111001",
			3668 => "0010001100110000000100",
			3669 => "0000001011100101111001",
			3670 => "0000000011100101111001",
			3671 => "0001011011000000001000",
			3672 => "0001111110001100000100",
			3673 => "0000000011100101111001",
			3674 => "0000001011100101111001",
			3675 => "0000111010100000000100",
			3676 => "0000001011100101111001",
			3677 => "1111111011100101111001",
			3678 => "0010001000000001000100",
			3679 => "0011011001001000101100",
			3680 => "0011001100101000100000",
			3681 => "0010010011000000011000",
			3682 => "0000100000100100001100",
			3683 => "0001111100010000000100",
			3684 => "0000000011101000111101",
			3685 => "0010111110011000000100",
			3686 => "0000000011101000111101",
			3687 => "0000000011101000111101",
			3688 => "0001010001001000000100",
			3689 => "1111111011101000111101",
			3690 => "0001011110111000000100",
			3691 => "0000000011101000111101",
			3692 => "0000000011101000111101",
			3693 => "0010101001011000000100",
			3694 => "0000000011101000111101",
			3695 => "0000000011101000111101",
			3696 => "0001110001001000001000",
			3697 => "0010011111011000000100",
			3698 => "1111111011101000111101",
			3699 => "0000000011101000111101",
			3700 => "0000000011101000111101",
			3701 => "0000000100010100001100",
			3702 => "0011110100001000001000",
			3703 => "0001101111110100000100",
			3704 => "0000000011101000111101",
			3705 => "0000000011101000111101",
			3706 => "0000000011101000111101",
			3707 => "0000100101101000001000",
			3708 => "0000001111001100000100",
			3709 => "0000001011101000111101",
			3710 => "0000000011101000111101",
			3711 => "0000000011101000111101",
			3712 => "0000101111001100011000",
			3713 => "0010100000111100001100",
			3714 => "0001101100011000000100",
			3715 => "0000000011101000111101",
			3716 => "0001100101111100000100",
			3717 => "0000001011101000111101",
			3718 => "0000000011101000111101",
			3719 => "0000100110100100001000",
			3720 => "0001100110000100000100",
			3721 => "0000000011101000111101",
			3722 => "0000000011101000111101",
			3723 => "0000000011101000111101",
			3724 => "0000111001010000000100",
			3725 => "0000000011101000111101",
			3726 => "0000000011101000111101",
			3727 => "0011010111011100010000",
			3728 => "0010011111011000001000",
			3729 => "0010000000110000000100",
			3730 => "1111111011101011100001",
			3731 => "0000000011101011100001",
			3732 => "0010001001000100000100",
			3733 => "0000000011101011100001",
			3734 => "0000000011101011100001",
			3735 => "0010001000000000101000",
			3736 => "0001111110111000100000",
			3737 => "0011100001000000011000",
			3738 => "0001110001001000010000",
			3739 => "0000100110010100001000",
			3740 => "0010011000000100000100",
			3741 => "0000000011101011100001",
			3742 => "1111111011101011100001",
			3743 => "0011011100101000000100",
			3744 => "1111111011101011100001",
			3745 => "0000000011101011100001",
			3746 => "0000010110001100000100",
			3747 => "0000000011101011100001",
			3748 => "0000001011101011100001",
			3749 => "0001010011000100000100",
			3750 => "1111111011101011100001",
			3751 => "0000000011101011100001",
			3752 => "0000111010100000000100",
			3753 => "0000001011101011100001",
			3754 => "0000000011101011100001",
			3755 => "0000111001010000010100",
			3756 => "0000101111001100010000",
			3757 => "0011100110110000001000",
			3758 => "0010001000111000000100",
			3759 => "0000000011101011100001",
			3760 => "0000000011101011100001",
			3761 => "0001100111010000000100",
			3762 => "0000001011101011100001",
			3763 => "0000000011101011100001",
			3764 => "0000000011101011100001",
			3765 => "0000111100110100000100",
			3766 => "0000001011101011100001",
			3767 => "1111111011101011100001",
			3768 => "0010001111011000100000",
			3769 => "0000010011110000000100",
			3770 => "1111111011101101101101",
			3771 => "0011110111010000010100",
			3772 => "0011111101100000001100",
			3773 => "0011111001110000000100",
			3774 => "1111111011101101101101",
			3775 => "0011111111110000000100",
			3776 => "0000001011101101101101",
			3777 => "1111111011101101101101",
			3778 => "0011111010101100000100",
			3779 => "0000001011101101101101",
			3780 => "0000000011101101101101",
			3781 => "0000001000001100000100",
			3782 => "1111111011101101101101",
			3783 => "0000000011101101101101",
			3784 => "0011111010011000000100",
			3785 => "1111111011101101101101",
			3786 => "0000110000111000100000",
			3787 => "0001010011000100010000",
			3788 => "0001001010000100000100",
			3789 => "0000001011101101101101",
			3790 => "0011011001001000000100",
			3791 => "1111111011101101101101",
			3792 => "0011110110011000000100",
			3793 => "0000001011101101101101",
			3794 => "0000000011101101101101",
			3795 => "0001110000111100001000",
			3796 => "0000111011111000000100",
			3797 => "0000001011101101101101",
			3798 => "0000000011101101101101",
			3799 => "0010000011100100000100",
			3800 => "0000001011101101101101",
			3801 => "0000001011101101101101",
			3802 => "1111111011101101101101",
			3803 => "0011011101101001001000",
			3804 => "0000100100010100101100",
			3805 => "0011110000000100100000",
			3806 => "0011111100111000011100",
			3807 => "0011010101010100010000",
			3808 => "0001010011001000001000",
			3809 => "0010001111001000000100",
			3810 => "0000000011110000111001",
			3811 => "0000000011110000111001",
			3812 => "0011100010001000000100",
			3813 => "0000000011110000111001",
			3814 => "0000000011110000111001",
			3815 => "0011111010011000000100",
			3816 => "0000000011110000111001",
			3817 => "0011000110000000000100",
			3818 => "0000000011110000111001",
			3819 => "0000000011110000111001",
			3820 => "0000000011110000111001",
			3821 => "0001011001010000000100",
			3822 => "0000000011110000111001",
			3823 => "0001001000000000000100",
			3824 => "0000000011110000111001",
			3825 => "0000000011110000111001",
			3826 => "0001001000000000010000",
			3827 => "0010101101001000001000",
			3828 => "0001011000111000000100",
			3829 => "0000000011110000111001",
			3830 => "0000000011110000111001",
			3831 => "0001010011000100000100",
			3832 => "0000000011110000111001",
			3833 => "0000000011110000111001",
			3834 => "0000111011000000001000",
			3835 => "0011010101010100000100",
			3836 => "0000000011110000111001",
			3837 => "0000000011110000111001",
			3838 => "0000000011110000111001",
			3839 => "0001000110101100010000",
			3840 => "0010001001010100001000",
			3841 => "0000000001110100000100",
			3842 => "0000000011110000111001",
			3843 => "0000000011110000111001",
			3844 => "0001100101111100000100",
			3845 => "0000000011110000111001",
			3846 => "0000000011110000111001",
			3847 => "0011011010000100000100",
			3848 => "0000000011110000111001",
			3849 => "0000010111011100000100",
			3850 => "0000000011110000111001",
			3851 => "0000000010100100000100",
			3852 => "0000000011110000111001",
			3853 => "0000000011110000111001",
			3854 => "0011100010110100111100",
			3855 => "0000101000010000110000",
			3856 => "0011100110111000101100",
			3857 => "0011110000000100011100",
			3858 => "0010101001010100001100",
			3859 => "0011100010011100000100",
			3860 => "0000000011110011100101",
			3861 => "0011000111011100000100",
			3862 => "0000000011110011100101",
			3863 => "0000000011110011100101",
			3864 => "0011010101101100001000",
			3865 => "0001110000111100000100",
			3866 => "0000000011110011100101",
			3867 => "0000000011110011100101",
			3868 => "0010110101111000000100",
			3869 => "0000000011110011100101",
			3870 => "0000000011110011100101",
			3871 => "0001001100000000001000",
			3872 => "0010010011000000000100",
			3873 => "0000000011110011100101",
			3874 => "0000000011110011100101",
			3875 => "0000111011111000000100",
			3876 => "0000000011110011100101",
			3877 => "0000000011110011100101",
			3878 => "0000000011110011100101",
			3879 => "0010110101010100001000",
			3880 => "0010110111011100000100",
			3881 => "0000000011110011100101",
			3882 => "0000000011110011100101",
			3883 => "0000000011110011100101",
			3884 => "0000010111011100010000",
			3885 => "0001010011000100001000",
			3886 => "0001101110000100000100",
			3887 => "0000000011110011100101",
			3888 => "0000000011110011100101",
			3889 => "0001101110000100000100",
			3890 => "0000000011110011100101",
			3891 => "0000000011110011100101",
			3892 => "0000011100101000000100",
			3893 => "0000000011110011100101",
			3894 => "0010010110101100000100",
			3895 => "0000000011110011100101",
			3896 => "0000000011110011100101",
			3897 => "0000011001100000000100",
			3898 => "1111111011110101001001",
			3899 => "0010101000111000001000",
			3900 => "0001101100100000000100",
			3901 => "1111111011110101001001",
			3902 => "0000001011110101001001",
			3903 => "0010010110000000000100",
			3904 => "1111111011110101001001",
			3905 => "0011110000001100010000",
			3906 => "0011111010011000000100",
			3907 => "1111111011110101001001",
			3908 => "0001000110011100001000",
			3909 => "0011001101101000000100",
			3910 => "0000001011110101001001",
			3911 => "0000000011110101001001",
			3912 => "0000000011110101001001",
			3913 => "0001111011111000001000",
			3914 => "0001010001010000000100",
			3915 => "0000000011110101001001",
			3916 => "1111111011110101001001",
			3917 => "0000111100010000000100",
			3918 => "0000000011110101001001",
			3919 => "0011011001001000000100",
			3920 => "0000000011110101001001",
			3921 => "0000000011110101001001",
			3922 => "0011010111011100010100",
			3923 => "0010001111001000000100",
			3924 => "1111111011110111110101",
			3925 => "0001010011001000001000",
			3926 => "0000000000100000000100",
			3927 => "0000000011110111110101",
			3928 => "0000001011110111110101",
			3929 => "0001001000111000000100",
			3930 => "1111111011110111110101",
			3931 => "0000000011110111110101",
			3932 => "0001111100011100110100",
			3933 => "0000101111001100101100",
			3934 => "0011000101111000011000",
			3935 => "0010001000000000010000",
			3936 => "0000111000101000001000",
			3937 => "0001011001010000000100",
			3938 => "0000000011110111110101",
			3939 => "0000001011110111110101",
			3940 => "0010000011001000000100",
			3941 => "1111111011110111110101",
			3942 => "0000000011110111110101",
			3943 => "0001001100000000000100",
			3944 => "0000000011110111110101",
			3945 => "0000001011110111110101",
			3946 => "0010100000111100001000",
			3947 => "0001001001001000000100",
			3948 => "1111111011110111110101",
			3949 => "0000000011110111110101",
			3950 => "0001110001011000001000",
			3951 => "0001110001001000000100",
			3952 => "1111111011110111110101",
			3953 => "0000000011110111110101",
			3954 => "1111111011110111110101",
			3955 => "0001101110000100000100",
			3956 => "1111111011110111110101",
			3957 => "0000000011110111110101",
			3958 => "0001011011000000001000",
			3959 => "0010101111101000000100",
			3960 => "0000001011110111110101",
			3961 => "0000000011110111110101",
			3962 => "0000111010100000000100",
			3963 => "0000001011110111110101",
			3964 => "1111111011110111110101",
			3965 => "0000010110001100100000",
			3966 => "0010000000110000010000",
			3967 => "0000010011110000000100",
			3968 => "1111111011111010010001",
			3969 => "0011000101010100001000",
			3970 => "0010011001000100000100",
			3971 => "1111111011111010010001",
			3972 => "0000000011111010010001",
			3973 => "1111111011111010010001",
			3974 => "0011001001000100001100",
			3975 => "0001111101001000000100",
			3976 => "1111111011111010010001",
			3977 => "0001011100101100000100",
			3978 => "0000000011111010010001",
			3979 => "0000001011111010010001",
			3980 => "1111111011111010010001",
			3981 => "0011111010011000000100",
			3982 => "1111111011111010010001",
			3983 => "0010101110010100101000",
			3984 => "0011011101101000010100",
			3985 => "0011111100111000000100",
			3986 => "0000001011111010010001",
			3987 => "0001111001011000001000",
			3988 => "0011110000001000000100",
			3989 => "0000000011111010010001",
			3990 => "1111111011111010010001",
			3991 => "0000111100110000000100",
			3992 => "0000000011111010010001",
			3993 => "0000001011111010010001",
			3994 => "0000010111011100001000",
			3995 => "0001011000100000000100",
			3996 => "0000000011111010010001",
			3997 => "0000001011111010010001",
			3998 => "0000111001010000001000",
			3999 => "0011000101111000000100",
			4000 => "0000001011111010010001",
			4001 => "0000001011111010010001",
			4002 => "0000001011111010010001",
			4003 => "1111111011111010010001",
			4004 => "0010001111011000100000",
			4005 => "0000010011110000000100",
			4006 => "1111111011111100100101",
			4007 => "0011110111010000010100",
			4008 => "0011111101100000001100",
			4009 => "0000010110001100000100",
			4010 => "1111111011111100100101",
			4011 => "0001110110101100000100",
			4012 => "0000000011111100100101",
			4013 => "1111111011111100100101",
			4014 => "0000001011001000000100",
			4015 => "0000001011111100100101",
			4016 => "0000000011111100100101",
			4017 => "0011100100000100000100",
			4018 => "1111111011111100100101",
			4019 => "0000000011111100100101",
			4020 => "0011111010011000000100",
			4021 => "1111111011111100100101",
			4022 => "0000110000111000100100",
			4023 => "0001111100011100010100",
			4024 => "0000101111001100010000",
			4025 => "0011111101010000001000",
			4026 => "0010110110000000000100",
			4027 => "0000001011111100100101",
			4028 => "0000001011111100100101",
			4029 => "0001111001011000000100",
			4030 => "0000000011111100100101",
			4031 => "0000001011111100100101",
			4032 => "1111111011111100100101",
			4033 => "0001011011000000001000",
			4034 => "0000001001101000000100",
			4035 => "0000001011111100100101",
			4036 => "0000000011111100100101",
			4037 => "0011001101101000000100",
			4038 => "0000001011111100100101",
			4039 => "0000001011111100100101",
			4040 => "1111111011111100100101",
			4041 => "0010001111011000100100",
			4042 => "0011111010111100011100",
			4043 => "0001100010110000010100",
			4044 => "0000011101000000000100",
			4045 => "0000000011111111001001",
			4046 => "0001111100110000001000",
			4047 => "0000110011001000000100",
			4048 => "0000000011111111001001",
			4049 => "0000000011111111001001",
			4050 => "0001100110100000000100",
			4051 => "0000000011111111001001",
			4052 => "0000000011111111001001",
			4053 => "0000011001100000000100",
			4054 => "0000000011111111001001",
			4055 => "0000000011111111001001",
			4056 => "0001001100110000000100",
			4057 => "1111111011111111001001",
			4058 => "0000000011111111001001",
			4059 => "0000111100110100101100",
			4060 => "0001011000100000100000",
			4061 => "0010101001011000011100",
			4062 => "0010111101101000010000",
			4063 => "0011111100111100001000",
			4064 => "0000101100010100000100",
			4065 => "0000000011111111001001",
			4066 => "0000000011111111001001",
			4067 => "0011001001000100000100",
			4068 => "0000000011111111001001",
			4069 => "0000000011111111001001",
			4070 => "0000000001110100000100",
			4071 => "0000000011111111001001",
			4072 => "0011100111101000000100",
			4073 => "0000001011111111001001",
			4074 => "0000000011111111001001",
			4075 => "0000000011111111001001",
			4076 => "0011000101101100000100",
			4077 => "0000000011111111001001",
			4078 => "0011100001000100000100",
			4079 => "0000000011111111001001",
			4080 => "0000001011111111001001",
			4081 => "0000000011111111001001",
			4082 => "0010000000110000100100",
			4083 => "0010111010100100001100",
			4084 => "0001000110000000000100",
			4085 => "0000000100000010001101",
			4086 => "0000010011110000000100",
			4087 => "0000000100000010001101",
			4088 => "0000000100000010001101",
			4089 => "0000100001000000001000",
			4090 => "0000100100010000000100",
			4091 => "0000000100000010001101",
			4092 => "0000000100000010001101",
			4093 => "0001110001011000001100",
			4094 => "0001000101011100001000",
			4095 => "0001000101010100000100",
			4096 => "0000000100000010001101",
			4097 => "0000000100000010001101",
			4098 => "0000000100000010001101",
			4099 => "0000000100000010001101",
			4100 => "0010101100001100110100",
			4101 => "0001011000100000101000",
			4102 => "0000101111001100100000",
			4103 => "0010000011100100010000",
			4104 => "0010101001010100001000",
			4105 => "0001111101001000000100",
			4106 => "0000000100000010001101",
			4107 => "0000000100000010001101",
			4108 => "0010010101111000000100",
			4109 => "0000000100000010001101",
			4110 => "0000000100000010001101",
			4111 => "0011000101111000001000",
			4112 => "0000000100010100000100",
			4113 => "0000000100000010001101",
			4114 => "0000000100000010001101",
			4115 => "0001101010110000000100",
			4116 => "0000000100000010001101",
			4117 => "0000000100000010001101",
			4118 => "0001110011110100000100",
			4119 => "0000000100000010001101",
			4120 => "0000000100000010001101",
			4121 => "0011110000000100001000",
			4122 => "0000001100001000000100",
			4123 => "0000000100000010001101",
			4124 => "0000000100000010001101",
			4125 => "0000000100000010001101",
			4126 => "0000010101010100001000",
			4127 => "0001111010011100000100",
			4128 => "0000000100000010001101",
			4129 => "0000000100000010001101",
			4130 => "0000000100000010001101",
			4131 => "0010000011100101001000",
			4132 => "0010101001010100010000",
			4133 => "0010011001000100000100",
			4134 => "0000000100000101101001",
			4135 => "0001101010011000000100",
			4136 => "0000000100000101101001",
			4137 => "0010001111001000000100",
			4138 => "0000000100000101101001",
			4139 => "0000000100000101101001",
			4140 => "0001010001001000011100",
			4141 => "0000000100111100001000",
			4142 => "0000001000110100000100",
			4143 => "0000000100000101101001",
			4144 => "0000000100000101101001",
			4145 => "0000101001101000010000",
			4146 => "0001001001001000001000",
			4147 => "0000000100010100000100",
			4148 => "0000000100000101101001",
			4149 => "0000000100000101101001",
			4150 => "0000001001101000000100",
			4151 => "0000000100000101101001",
			4152 => "0000000100000101101001",
			4153 => "0000000100000101101001",
			4154 => "0010100011110100010100",
			4155 => "0011110000000100001100",
			4156 => "0010101001000000001000",
			4157 => "0001011110111000000100",
			4158 => "0000000100000101101001",
			4159 => "0000000100000101101001",
			4160 => "0000000100000101101001",
			4161 => "0011010101011100000100",
			4162 => "0000000100000101101001",
			4163 => "0000000100000101101001",
			4164 => "0001111100011100000100",
			4165 => "0000000100000101101001",
			4166 => "0000000100000101101001",
			4167 => "0001000011000000010000",
			4168 => "0000111000000000001100",
			4169 => "0010001000000000000100",
			4170 => "0000000100000101101001",
			4171 => "0010111000000100000100",
			4172 => "0000000100000101101001",
			4173 => "0000000100000101101001",
			4174 => "0000000100000101101001",
			4175 => "0000011110011000001000",
			4176 => "0000100011100000000100",
			4177 => "0000000100000101101001",
			4178 => "0000000100000101101001",
			4179 => "0010001001010100001000",
			4180 => "0000111110001100000100",
			4181 => "0000000100000101101001",
			4182 => "0000000100000101101001",
			4183 => "0011101010001000000100",
			4184 => "0000000100000101101001",
			4185 => "0000000100000101101001",
			4186 => "0001111100011101000000",
			4187 => "0000101111001100110100",
			4188 => "0000011001100000000100",
			4189 => "1111111100001000010101",
			4190 => "0010011000000100011000",
			4191 => "0010010011001000010000",
			4192 => "0000100110010100001000",
			4193 => "0001111100010000000100",
			4194 => "1111111100001000010101",
			4195 => "0000000100001000010101",
			4196 => "0001100100100000000100",
			4197 => "1111111100001000010101",
			4198 => "0000000100001000010101",
			4199 => "0011110011101000000100",
			4200 => "0000000100001000010101",
			4201 => "0000001100001000010101",
			4202 => "0000111100110000001100",
			4203 => "0000010011010000001000",
			4204 => "0011001010000100000100",
			4205 => "0000001100001000010101",
			4206 => "0000000100001000010101",
			4207 => "1111111100001000010101",
			4208 => "0001011011111000000100",
			4209 => "0000001100001000010101",
			4210 => "0000010111011100000100",
			4211 => "0000000100001000010101",
			4212 => "0000001100001000010101",
			4213 => "0011101110010000000100",
			4214 => "1111111100001000010101",
			4215 => "0000111101001000000100",
			4216 => "0000000100001000010101",
			4217 => "0000000100001000010101",
			4218 => "0011000011000000001000",
			4219 => "0000100101010000000100",
			4220 => "0000001100001000010101",
			4221 => "0000000100001000010101",
			4222 => "0011010011000000001000",
			4223 => "0001011010011100000100",
			4224 => "0000000100001000010101",
			4225 => "0000000100001000010101",
			4226 => "0000101011111100000100",
			4227 => "0000000100001000010101",
			4228 => "0000001100001000010101",
			4229 => "0001110011110101001100",
			4230 => "0011000110000000111000",
			4231 => "0001111001011000101000",
			4232 => "0000100010100100010100",
			4233 => "0001111100010000000100",
			4234 => "0000000100001011011001",
			4235 => "0010101001011000001000",
			4236 => "0010010011000000000100",
			4237 => "0000000100001011011001",
			4238 => "0000001100001011011001",
			4239 => "0010010011001000000100",
			4240 => "0000000100001011011001",
			4241 => "0000000100001011011001",
			4242 => "0001100111101000001000",
			4243 => "0001100100000100000100",
			4244 => "0000000100001011011001",
			4245 => "0000000100001011011001",
			4246 => "0000011101000000001000",
			4247 => "0001010110011100000100",
			4248 => "0000000100001011011001",
			4249 => "0000000100001011011001",
			4250 => "1111111100001011011001",
			4251 => "0001010001010000000100",
			4252 => "0000000100001011011001",
			4253 => "0000001110101000001000",
			4254 => "0001101100111000000100",
			4255 => "0000000100001011011001",
			4256 => "0000001100001011011001",
			4257 => "0000000100001011011001",
			4258 => "0011111001111000001100",
			4259 => "0001101010001000000100",
			4260 => "0000000100001011011001",
			4261 => "0001111001000000000100",
			4262 => "0000000100001011011001",
			4263 => "0000000100001011011001",
			4264 => "0001010011000100000100",
			4265 => "0000000100001011011001",
			4266 => "0000000100001011011001",
			4267 => "0011000011000000000100",
			4268 => "0000001100001011011001",
			4269 => "0010000110101100001100",
			4270 => "0000111111101000000100",
			4271 => "0000000100001011011001",
			4272 => "0000111111110000000100",
			4273 => "0000000100001011011001",
			4274 => "0000000100001011011001",
			4275 => "0000000010100100000100",
			4276 => "0000000100001011011001",
			4277 => "0000000100001011011001",
			4278 => "0010000000110000100100",
			4279 => "0010111010100100001100",
			4280 => "0001000110000000000100",
			4281 => "0000000100001110110101",
			4282 => "0011011010100100000100",
			4283 => "0000000100001110110101",
			4284 => "0000000100001110110101",
			4285 => "0000100001000000001000",
			4286 => "0000100100010000000100",
			4287 => "0000000100001110110101",
			4288 => "0000000100001110110101",
			4289 => "0001110001011000001100",
			4290 => "0001000101011100001000",
			4291 => "0001000101010100000100",
			4292 => "0000000100001110110101",
			4293 => "0000000100001110110101",
			4294 => "0000000100001110110101",
			4295 => "0000000100001110110101",
			4296 => "0010100000111100111000",
			4297 => "0000101111001100101100",
			4298 => "0010000011100100011000",
			4299 => "0011000110000000001100",
			4300 => "0011101110100100001000",
			4301 => "0001001111011000000100",
			4302 => "0000000100001110110101",
			4303 => "0000000100001110110101",
			4304 => "0000000100001110110101",
			4305 => "0010011000111000000100",
			4306 => "0000000100001110110101",
			4307 => "0010011100010000000100",
			4308 => "0000000100001110110101",
			4309 => "0000000100001110110101",
			4310 => "0000011100101000001100",
			4311 => "0011100001100000001000",
			4312 => "0001100000110100000100",
			4313 => "0000000100001110110101",
			4314 => "0000001100001110110101",
			4315 => "0000000100001110110101",
			4316 => "0000000110111100000100",
			4317 => "0000000100001110110101",
			4318 => "0000000100001110110101",
			4319 => "0001110011110100000100",
			4320 => "0000000100001110110101",
			4321 => "0000011100101000000100",
			4322 => "0000000100001110110101",
			4323 => "0000000100001110110101",
			4324 => "0001001001010000001100",
			4325 => "0001011100011100000100",
			4326 => "0000000100001110110101",
			4327 => "0011101000101100000100",
			4328 => "0000000100001110110101",
			4329 => "0000000100001110110101",
			4330 => "0000110000111000000100",
			4331 => "0000000100001110110101",
			4332 => "0000000100001110110101",
			4333 => "0010001111011000111000",
			4334 => "0011101110100000110000",
			4335 => "0001111000101000100000",
			4336 => "0010101100010000010100",
			4337 => "0001001010000100001100",
			4338 => "0011000111011100000100",
			4339 => "0000000100010010011001",
			4340 => "0011000101011100000100",
			4341 => "0000000100010010011001",
			4342 => "0000000100010010011001",
			4343 => "0001011001010100000100",
			4344 => "0000000100010010011001",
			4345 => "0000000100010010011001",
			4346 => "0010111010100100001000",
			4347 => "0010111110011000000100",
			4348 => "0000000100010010011001",
			4349 => "0000000100010010011001",
			4350 => "0000000100010010011001",
			4351 => "0001000110011100001100",
			4352 => "0000001000010000001000",
			4353 => "0000010011110000000100",
			4354 => "0000000100010010011001",
			4355 => "0000000100010010011001",
			4356 => "0000000100010010011001",
			4357 => "0000000100010010011001",
			4358 => "0011100101001100000100",
			4359 => "1111111100010010011001",
			4360 => "0000000100010010011001",
			4361 => "0010100000111100100100",
			4362 => "0000001010111000011000",
			4363 => "0011100110110000001100",
			4364 => "0011110100001000001000",
			4365 => "0011111010011000000100",
			4366 => "0000000100010010011001",
			4367 => "0000000100010010011001",
			4368 => "0000000100010010011001",
			4369 => "0011000110000000000100",
			4370 => "0000001100010010011001",
			4371 => "0010001000111000000100",
			4372 => "0000000100010010011001",
			4373 => "0000000100010010011001",
			4374 => "0011011101101000000100",
			4375 => "0000000100010010011001",
			4376 => "0001001000000000000100",
			4377 => "0000000100010010011001",
			4378 => "0000000100010010011001",
			4379 => "0001101110000100010100",
			4380 => "0000010111011100001100",
			4381 => "0000000110111100001000",
			4382 => "0000001101110100000100",
			4383 => "0000000100010010011001",
			4384 => "0000000100010010011001",
			4385 => "0000000100010010011001",
			4386 => "0000000010100100000100",
			4387 => "0000000100010010011001",
			4388 => "0000000100010010011001",
			4389 => "0000000100010010011001",
			4390 => "0010001111011000100100",
			4391 => "0011111010111100011100",
			4392 => "0001100010110000010100",
			4393 => "0000011101000000000100",
			4394 => "0000000100010101010101",
			4395 => "0001111100110000001000",
			4396 => "0000110011001000000100",
			4397 => "0000000100010101010101",
			4398 => "0000000100010101010101",
			4399 => "0001100110100000000100",
			4400 => "0000000100010101010101",
			4401 => "0000000100010101010101",
			4402 => "0000011001100000000100",
			4403 => "0000000100010101010101",
			4404 => "0000000100010101010101",
			4405 => "0001001100110000000100",
			4406 => "1111111100010101010101",
			4407 => "0000000100010101010101",
			4408 => "0000111100110100111000",
			4409 => "0001011000100000011100",
			4410 => "0000111111101000010100",
			4411 => "0000111001010000001100",
			4412 => "0011001001001000000100",
			4413 => "0000000100010101010101",
			4414 => "0011011101101000000100",
			4415 => "0000000100010101010101",
			4416 => "0000000100010101010101",
			4417 => "0000100011001100000100",
			4418 => "0000000100010101010101",
			4419 => "0000001100010101010101",
			4420 => "0010101011000000000100",
			4421 => "0000000100010101010101",
			4422 => "0000000100010101010101",
			4423 => "0000111011000000010000",
			4424 => "0010100011000100001100",
			4425 => "0010101011000000000100",
			4426 => "0000000100010101010101",
			4427 => "0001100100100000000100",
			4428 => "0000000100010101010101",
			4429 => "0000000100010101010101",
			4430 => "0000001100010101010101",
			4431 => "0001011010011100000100",
			4432 => "0000000100010101010101",
			4433 => "0001100001111000000100",
			4434 => "0000000100010101010101",
			4435 => "0000000100010101010101",
			4436 => "0000000100010101010101",
			4437 => "0010001111011000101000",
			4438 => "0000111011111000100000",
			4439 => "0001100001000000011100",
			4440 => "0001100010110000010100",
			4441 => "0001010110011100001100",
			4442 => "0000100001000000001000",
			4443 => "0000000111100000000100",
			4444 => "0000000100011000101001",
			4445 => "0000000100011000101001",
			4446 => "0000000100011000101001",
			4447 => "0000001100111000000100",
			4448 => "0000000100011000101001",
			4449 => "0000000100011000101001",
			4450 => "0000110011001000000100",
			4451 => "0000000100011000101001",
			4452 => "0000000100011000101001",
			4453 => "0000000100011000101001",
			4454 => "0010101001011000000100",
			4455 => "0000000100011000101001",
			4456 => "0000000100011000101001",
			4457 => "0000101111001100110100",
			4458 => "0000111111101000011100",
			4459 => "0010011000000100001000",
			4460 => "0011111010011000000100",
			4461 => "0000000100011000101001",
			4462 => "0000000100011000101001",
			4463 => "0001000011000000001100",
			4464 => "0010001100110000001000",
			4465 => "0001001100101000000100",
			4466 => "0000000100011000101001",
			4467 => "0000000100011000101001",
			4468 => "0000000100011000101001",
			4469 => "0011001101101000000100",
			4470 => "0000000100011000101001",
			4471 => "0000000100011000101001",
			4472 => "0001010011000100000100",
			4473 => "0000000100011000101001",
			4474 => "0000110011000100001000",
			4475 => "0010100011000100000100",
			4476 => "0000000100011000101001",
			4477 => "0000000100011000101001",
			4478 => "0001111000100000000100",
			4479 => "0000000100011000101001",
			4480 => "0000110000111000000100",
			4481 => "0000000100011000101001",
			4482 => "0000000100011000101001",
			4483 => "0010110011000000001100",
			4484 => "0000111001010000000100",
			4485 => "0000000100011000101001",
			4486 => "0001100101111100000100",
			4487 => "0000000100011000101001",
			4488 => "0000000100011000101001",
			4489 => "0000000100011000101001",
			4490 => "0011100010110101001000",
			4491 => "0000001010010100111100",
			4492 => "0011100110111000110100",
			4493 => "0000011110011000100000",
			4494 => "0001000011000000010000",
			4495 => "0001001001000100001000",
			4496 => "0000010110001100000100",
			4497 => "0000000100011100000101",
			4498 => "0000000100011100000101",
			4499 => "0000010011110000000100",
			4500 => "0000000100011100000101",
			4501 => "0000000100011100000101",
			4502 => "0000111001010100001000",
			4503 => "0001011011111000000100",
			4504 => "0000000100011100000101",
			4505 => "0000000100011100000101",
			4506 => "0010001111011000000100",
			4507 => "0000000100011100000101",
			4508 => "0000000100011100000101",
			4509 => "0000101100010100010000",
			4510 => "0000011010100100001000",
			4511 => "0001111100101100000100",
			4512 => "0000000100011100000101",
			4513 => "0000000100011100000101",
			4514 => "0000111000000000000100",
			4515 => "0000000100011100000101",
			4516 => "0000000100011100000101",
			4517 => "0000001100011100000101",
			4518 => "0001010011000100000100",
			4519 => "0000000100011100000101",
			4520 => "0000000100011100000101",
			4521 => "0010110101101100001000",
			4522 => "0001001100010000000100",
			4523 => "1111111100011100000101",
			4524 => "0000000100011100000101",
			4525 => "0000000100011100000101",
			4526 => "0000111001010000011000",
			4527 => "0010101000101000001000",
			4528 => "0001000101010100000100",
			4529 => "0000000100011100000101",
			4530 => "0000000100011100000101",
			4531 => "0000101101111000001000",
			4532 => "0000010110001100000100",
			4533 => "0000000100011100000101",
			4534 => "0000000100011100000101",
			4535 => "0011111110011100000100",
			4536 => "1111111100011100000101",
			4537 => "0000000100011100000101",
			4538 => "0010100000111100001000",
			4539 => "0010110101010100000100",
			4540 => "0000000100011100000101",
			4541 => "0000001100011100000101",
			4542 => "0011101110010000000100",
			4543 => "0000000100011100000101",
			4544 => "0000000100011100000101",
			4545 => "0010001000000001100000",
			4546 => "0011011001001000111000",
			4547 => "0011001100101000100000",
			4548 => "0010010011000000011000",
			4549 => "0000100000100100001100",
			4550 => "0001111100010000000100",
			4551 => "0000000100100000011001",
			4552 => "0010111110011000000100",
			4553 => "0000000100100000011001",
			4554 => "0000000100100000011001",
			4555 => "0001010001001000000100",
			4556 => "1111111100100000011001",
			4557 => "0001011110111000000100",
			4558 => "0000000100100000011001",
			4559 => "0000000100100000011001",
			4560 => "0010101001011000000100",
			4561 => "0000000100100000011001",
			4562 => "0000000100100000011001",
			4563 => "0001010001001000001100",
			4564 => "0001100110000100001000",
			4565 => "0000000110011000000100",
			4566 => "0000000100100000011001",
			4567 => "0000000100100000011001",
			4568 => "1111111100100000011001",
			4569 => "0010100000111100000100",
			4570 => "0000000100100000011001",
			4571 => "0001111000100000000100",
			4572 => "0000000100100000011001",
			4573 => "0000000100100000011001",
			4574 => "0000000100010100011100",
			4575 => "0010011000000100001000",
			4576 => "0000000100001000000100",
			4577 => "0000000100100000011001",
			4578 => "0000000100100000011001",
			4579 => "0001010011000100001100",
			4580 => "0010011000111000000100",
			4581 => "1111111100100000011001",
			4582 => "0011000011000000000100",
			4583 => "0000000100100000011001",
			4584 => "0000000100100000011001",
			4585 => "0000001110110100000100",
			4586 => "0000000100100000011001",
			4587 => "0000000100100000011001",
			4588 => "0000100111111000000100",
			4589 => "0000001100100000011001",
			4590 => "0011001001000100000100",
			4591 => "0000000100100000011001",
			4592 => "0000000100100000011001",
			4593 => "0001111110111000010000",
			4594 => "0000111100110000001000",
			4595 => "0010110011001000000100",
			4596 => "0000000100100000011001",
			4597 => "0000000100100000011001",
			4598 => "0000110001001000000100",
			4599 => "0000001100100000011001",
			4600 => "0000000100100000011001",
			4601 => "0001101010110000001100",
			4602 => "0000001111001100001000",
			4603 => "0001101100000100000100",
			4604 => "0000000100100000011001",
			4605 => "0000000100100000011001",
			4606 => "0000000100100000011001",
			4607 => "0000010101010100000100",
			4608 => "0000000100100000011001",
			4609 => "0000011100101000000100",
			4610 => "0000000100100000011001",
			4611 => "0000011001000100000100",
			4612 => "0000000100100000011001",
			4613 => "0000000100100000011001",
			4614 => "0010001111001000000100",
			4615 => "1111111100100010111101",
			4616 => "0000001101011100101000",
			4617 => "0001100010110000011100",
			4618 => "0011010101011100010100",
			4619 => "0000010011110000001100",
			4620 => "0001001010000100001000",
			4621 => "0001111100010000000100",
			4622 => "0000000100100010111101",
			4623 => "0000000100100010111101",
			4624 => "0000000100100010111101",
			4625 => "0001011000000000000100",
			4626 => "0000000100100010111101",
			4627 => "1111111100100010111101",
			4628 => "0010111001001000000100",
			4629 => "0000000100100010111101",
			4630 => "0000000100100010111101",
			4631 => "0010101001011000000100",
			4632 => "0000001100100010111101",
			4633 => "0001011100110100000100",
			4634 => "0000000100100010111101",
			4635 => "0000000100100010111101",
			4636 => "0010010110101100100000",
			4637 => "0010001111011000001000",
			4638 => "0000001000001100000100",
			4639 => "1111111100100010111101",
			4640 => "0000000100100010111101",
			4641 => "0001010011000100001100",
			4642 => "0001010110011100001000",
			4643 => "0000101011001100000100",
			4644 => "0000000100100010111101",
			4645 => "0000000100100010111101",
			4646 => "1111111100100010111101",
			4647 => "0001110000111100001000",
			4648 => "0001010001011000000100",
			4649 => "0000000100100010111101",
			4650 => "0000000100100010111101",
			4651 => "0000001100100010111101",
			4652 => "0011110000001000000100",
			4653 => "0000000100100010111101",
			4654 => "0000001100100010111101",
			4655 => "0010001111001000001100",
			4656 => "0000010011110000000100",
			4657 => "1111111100100101101001",
			4658 => "0001011001010000000100",
			4659 => "0000000100100101101001",
			4660 => "0000000100100101101001",
			4661 => "0010100000111100110100",
			4662 => "0001010001001000110000",
			4663 => "0011111100111100011000",
			4664 => "0001101100000100010000",
			4665 => "0010101001010100001000",
			4666 => "0001101010011000000100",
			4667 => "0000000100100101101001",
			4668 => "0000001100100101101001",
			4669 => "0001100100011100000100",
			4670 => "0000000100100101101001",
			4671 => "1111111100100101101001",
			4672 => "0010010011000000000100",
			4673 => "0000000100100101101001",
			4674 => "0000001100100101101001",
			4675 => "0011100010110100001100",
			4676 => "0001010001010000000100",
			4677 => "1111111100100101101001",
			4678 => "0000111000101000000100",
			4679 => "0000000100100101101001",
			4680 => "1111111100100101101001",
			4681 => "0010101111101000000100",
			4682 => "0000001100100101101001",
			4683 => "0001001000000000000100",
			4684 => "0000000100100101101001",
			4685 => "0000000100100101101001",
			4686 => "0000001100100101101001",
			4687 => "0011101110010000010100",
			4688 => "0000010111011100001100",
			4689 => "0001001001010000000100",
			4690 => "1111111100100101101001",
			4691 => "0001011001101100000100",
			4692 => "0000000100100101101001",
			4693 => "0000000100100101101001",
			4694 => "0010101110010100000100",
			4695 => "0000000100100101101001",
			4696 => "0000000100100101101001",
			4697 => "0000001100100101101001",
			4698 => "0000011001100000000100",
			4699 => "1111111100100111101101",
			4700 => "0010101111101000011000",
			4701 => "0001101010011000000100",
			4702 => "1111111100100111101101",
			4703 => "0010011001000100000100",
			4704 => "1111111100100111101101",
			4705 => "0011111100111000000100",
			4706 => "0000001100100111101101",
			4707 => "0010010011000000000100",
			4708 => "1111111100100111101101",
			4709 => "0011001101101000000100",
			4710 => "0000001100100111101101",
			4711 => "0000000100100111101101",
			4712 => "0001010001010000000100",
			4713 => "1111111100100111101101",
			4714 => "0010000000110000001000",
			4715 => "0001110000111100000100",
			4716 => "1111111100100111101101",
			4717 => "0000000100100111101101",
			4718 => "0000101100001000010000",
			4719 => "0010101001011000001000",
			4720 => "0000001010101000000100",
			4721 => "0000000100100111101101",
			4722 => "0000001100100111101101",
			4723 => "0001001100010000000100",
			4724 => "1111111100100111101101",
			4725 => "0000000100100111101101",
			4726 => "0001111001011000000100",
			4727 => "0000000100100111101101",
			4728 => "0001101101010000000100",
			4729 => "0000001100100111101101",
			4730 => "0000000100100111101101",
			4731 => "0011010101011100100000",
			4732 => "0001111100110000000100",
			4733 => "0000000100101010011001",
			4734 => "0000100110010100010100",
			4735 => "0010101001011000010000",
			4736 => "0010011001000100000100",
			4737 => "0000000100101010011001",
			4738 => "0011011010100100000100",
			4739 => "0000000100101010011001",
			4740 => "0000011001100000000100",
			4741 => "0000000100101010011001",
			4742 => "0000000100101010011001",
			4743 => "0000000100101010011001",
			4744 => "0011100101100000000100",
			4745 => "0000000100101010011001",
			4746 => "0000000100101010011001",
			4747 => "0000111100110100110100",
			4748 => "0001011000100000101100",
			4749 => "0000011110011000010000",
			4750 => "0010101011111000001100",
			4751 => "0010110101101100001000",
			4752 => "0010001010000100000100",
			4753 => "0000000100101010011001",
			4754 => "0000000100101010011001",
			4755 => "0000000100101010011001",
			4756 => "0000000100101010011001",
			4757 => "0001000011000000010000",
			4758 => "0001001001000100001000",
			4759 => "0011001100000000000100",
			4760 => "0000000100101010011001",
			4761 => "0000000100101010011001",
			4762 => "0011100011101000000100",
			4763 => "0000000100101010011001",
			4764 => "0000000100101010011001",
			4765 => "0000101111001100001000",
			4766 => "0010100100101100000100",
			4767 => "0000000100101010011001",
			4768 => "0000001100101010011001",
			4769 => "0000000100101010011001",
			4770 => "0000010110001100000100",
			4771 => "0000000100101010011001",
			4772 => "0000001100101010011001",
			4773 => "0000000100101010011001",
			4774 => "0010011001000100000100",
			4775 => "1111111100101100101101",
			4776 => "0010111010100100001000",
			4777 => "0000001110000100000100",
			4778 => "0000000100101100101101",
			4779 => "0000001100101100101101",
			4780 => "0001111100011100101000",
			4781 => "0010000000110000010100",
			4782 => "0010101101001000001100",
			4783 => "0011010111011100000100",
			4784 => "0000000100101100101101",
			4785 => "0001111001010000000100",
			4786 => "0000000100101100101101",
			4787 => "0000000100101100101101",
			4788 => "0001001001001000000100",
			4789 => "0000000100101100101101",
			4790 => "1111111100101100101101",
			4791 => "0000101111001100010000",
			4792 => "0010011000000100001000",
			4793 => "0001111001011000000100",
			4794 => "0000000100101100101101",
			4795 => "0000001100101100101101",
			4796 => "0000111100110000000100",
			4797 => "0000000100101100101101",
			4798 => "0000000100101100101101",
			4799 => "1111111100101100101101",
			4800 => "0011000011000000001000",
			4801 => "0000100101010000000100",
			4802 => "0000001100101100101101",
			4803 => "0000000100101100101101",
			4804 => "0011010011000000001000",
			4805 => "0001011010011100000100",
			4806 => "0000000100101100101101",
			4807 => "0000000100101100101101",
			4808 => "0000101011111100000100",
			4809 => "0000000100101100101101",
			4810 => "0000001100101100101101",
			4811 => "0001110011110101011100",
			4812 => "0011111100111100111100",
			4813 => "0000011110011000110000",
			4814 => "0001000011000000010100",
			4815 => "0000010011110000001000",
			4816 => "0010001111011000000100",
			4817 => "0000000100110000010001",
			4818 => "0000000100110000010001",
			4819 => "0001100011101100001000",
			4820 => "0010010110000000000100",
			4821 => "0000000100110000010001",
			4822 => "0000000100110000010001",
			4823 => "0000000100110000010001",
			4824 => "0001111011000000010000",
			4825 => "0010111010100100001000",
			4826 => "0000111100010000000100",
			4827 => "0000000100110000010001",
			4828 => "0000000100110000010001",
			4829 => "0010010011001000000100",
			4830 => "1111111100110000010001",
			4831 => "0000000100110000010001",
			4832 => "0001110110011100000100",
			4833 => "0000000100110000010001",
			4834 => "0011010101101100000100",
			4835 => "0000000100110000010001",
			4836 => "0000000100110000010001",
			4837 => "0010111100101000000100",
			4838 => "0000000100110000010001",
			4839 => "0010011101001000000100",
			4840 => "0000001100110000010001",
			4841 => "0000000100110000010001",
			4842 => "0001010011000100011000",
			4843 => "0000111000101000010100",
			4844 => "0000111001010000010000",
			4845 => "0001001001001000001000",
			4846 => "0001101110000100000100",
			4847 => "0000000100110000010001",
			4848 => "0000000100110000010001",
			4849 => "0001001111011000000100",
			4850 => "1111111100110000010001",
			4851 => "0000000100110000010001",
			4852 => "0000000100110000010001",
			4853 => "1111111100110000010001",
			4854 => "0001111000100000000100",
			4855 => "0000000100110000010001",
			4856 => "0000000100110000010001",
			4857 => "0011000011000000000100",
			4858 => "0000000100110000010001",
			4859 => "0010000110101100001100",
			4860 => "0000111111101000000100",
			4861 => "0000000100110000010001",
			4862 => "0000111111110000000100",
			4863 => "0000000100110000010001",
			4864 => "0000000100110000010001",
			4865 => "0000000010100100000100",
			4866 => "0000000100110000010001",
			4867 => "0000000100110000010001",
			4868 => "0000011001100000000100",
			4869 => "1111111100110010100101",
			4870 => "0010101111101000011000",
			4871 => "0001101010011000000100",
			4872 => "1111111100110010100101",
			4873 => "0010011001000100000100",
			4874 => "1111111100110010100101",
			4875 => "0001011000101000001100",
			4876 => "0010101001010100001000",
			4877 => "0001100101000000000100",
			4878 => "0000001100110010100101",
			4879 => "0000000100110010100101",
			4880 => "0000000100110010100101",
			4881 => "0000000100110010100101",
			4882 => "0001010001010000000100",
			4883 => "1111111100110010100101",
			4884 => "0010011111011000010000",
			4885 => "0010110101010100001000",
			4886 => "0001100111101000000100",
			4887 => "1111111100110010100101",
			4888 => "0000001100110010100101",
			4889 => "0001001001010100000100",
			4890 => "1111111100110010100101",
			4891 => "0000000100110010100101",
			4892 => "0000000101010000001100",
			4893 => "0000111000101000000100",
			4894 => "0000001100110010100101",
			4895 => "0000100011001100000100",
			4896 => "0000000100110010100101",
			4897 => "0000000100110010100101",
			4898 => "0001001000000000001000",
			4899 => "0001111100001100000100",
			4900 => "1111111100110010100101",
			4901 => "0000001100110010100101",
			4902 => "0001000110101100000100",
			4903 => "0000001100110010100101",
			4904 => "0000000100110010100101",
			4905 => "0011011101101001111000",
			4906 => "0001011100101101000100",
			4907 => "0011111100111000100000",
			4908 => "0001110110101100001100",
			4909 => "0011010101011100000100",
			4910 => "0000000100110111011001",
			4911 => "0011000101101100000100",
			4912 => "0000000100110111011001",
			4913 => "0000000100110111011001",
			4914 => "0000001110000100001100",
			4915 => "0010001111011000000100",
			4916 => "0000000100110111011001",
			4917 => "0011100011000000000100",
			4918 => "0000000100110111011001",
			4919 => "0000000100110111011001",
			4920 => "0000011001100000000100",
			4921 => "0000000100110111011001",
			4922 => "0000001100110111011001",
			4923 => "0011100110110000010000",
			4924 => "0001000110000000001000",
			4925 => "0001001001000100000100",
			4926 => "0000000100110111011001",
			4927 => "0000000100110111011001",
			4928 => "0001011100110000000100",
			4929 => "0000000100110111011001",
			4930 => "1111111100110111011001",
			4931 => "0011111011110100001000",
			4932 => "0001111100101100000100",
			4933 => "0000000100110111011001",
			4934 => "0000001100110111011001",
			4935 => "0011100010110100000100",
			4936 => "1111111100110111011001",
			4937 => "0010101000101000000100",
			4938 => "0000000100110111011001",
			4939 => "0000000100110111011001",
			4940 => "0011011001001000100100",
			4941 => "0011001001001000010000",
			4942 => "0001111011111000001100",
			4943 => "0000111001010000001000",
			4944 => "0001111100110000000100",
			4945 => "0000000100110111011001",
			4946 => "0000000100110111011001",
			4947 => "0000000100110111011001",
			4948 => "0000000100110111011001",
			4949 => "0011001001000100001100",
			4950 => "0001111011111000001000",
			4951 => "0001111001010000000100",
			4952 => "0000000100110111011001",
			4953 => "0000000100110111011001",
			4954 => "1111111100110111011001",
			4955 => "0011000110000000000100",
			4956 => "0000000100110111011001",
			4957 => "0000000100110111011001",
			4958 => "0000001110101000001100",
			4959 => "0000111110001100001000",
			4960 => "0001110110011100000100",
			4961 => "0000000100110111011001",
			4962 => "0000001100110111011001",
			4963 => "0000000100110111011001",
			4964 => "0000000100110111011001",
			4965 => "0001000110101100010000",
			4966 => "0010001001010100001000",
			4967 => "0000000001110100000100",
			4968 => "0000000100110111011001",
			4969 => "0000001100110111011001",
			4970 => "0011110100110100000100",
			4971 => "0000000100110111011001",
			4972 => "0000000100110111011001",
			4973 => "0011011010000100000100",
			4974 => "0000000100110111011001",
			4975 => "0000010111011100001000",
			4976 => "0010001000000000000100",
			4977 => "0000000100110111011001",
			4978 => "1111111100110111011001",
			4979 => "0000000010100100000100",
			4980 => "0000000100110111011001",
			4981 => "0000000100110111011001",
			4982 => "0001111100011101110000",
			4983 => "0010000011100101010000",
			4984 => "0010101111101000101100",
			4985 => "0010010110000000001100",
			4986 => "0001010101111000001000",
			4987 => "0010101000000000000100",
			4988 => "0000000100111011011111",
			4989 => "0000000100111011011111",
			4990 => "0000000100111011011111",
			4991 => "0000111000000000010000",
			4992 => "0010101000000000001000",
			4993 => "0000001110101100000100",
			4994 => "0000000100111011011111",
			4995 => "0000000100111011011111",
			4996 => "0000001010101100000100",
			4997 => "0000000100111011011111",
			4998 => "0000000100111011011111",
			4999 => "0001001010000100001000",
			5000 => "0001011100110000000100",
			5001 => "0000000100111011011111",
			5002 => "0000000100111011011111",
			5003 => "0000111101001000000100",
			5004 => "0000000100111011011111",
			5005 => "0000000100111011011111",
			5006 => "0000101100001000010100",
			5007 => "0001011100101100001000",
			5008 => "0011111100111100000100",
			5009 => "0000000100111011011111",
			5010 => "0000000100111011011111",
			5011 => "0001011001011000000100",
			5012 => "0000000100111011011111",
			5013 => "0010011111011000000100",
			5014 => "0000000100111011011111",
			5015 => "0000000100111011011111",
			5016 => "0001010001001000001100",
			5017 => "0001011011111000001000",
			5018 => "0001011111101000000100",
			5019 => "0000000100111011011111",
			5020 => "0000000100111011011111",
			5021 => "1111111100111011011111",
			5022 => "0000000100111011011111",
			5023 => "0000111100110000001100",
			5024 => "0000010011010000001000",
			5025 => "0001000101010100000100",
			5026 => "0000000100111011011111",
			5027 => "0000000100111011011111",
			5028 => "0000000100111011011111",
			5029 => "0010001100110000001100",
			5030 => "0000011110011000000100",
			5031 => "0000000100111011011111",
			5032 => "0000101010101000000100",
			5033 => "0000000100111011011111",
			5034 => "0000000100111011011111",
			5035 => "0010111101101000000100",
			5036 => "0000000100111011011111",
			5037 => "0000000100111011011111",
			5038 => "0000111010100000010000",
			5039 => "0000011100101000000100",
			5040 => "0000000100111011011111",
			5041 => "0011101000110100001000",
			5042 => "0000011001000100000100",
			5043 => "0000000100111011011111",
			5044 => "0000000100111011011111",
			5045 => "0000000100111011011111",
			5046 => "0000000100111011011111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1715, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3321, initial_addr_3'length));
	end generate gen_rom_0;

	gen_rom_1: if SELECT_ROM = 1 generate
		bank <= (
			0 => "0011101100011000010100",
			1 => "0000010111110000010000",
			2 => "0001111100010000000100",
			3 => "0000000000000001001101",
			4 => "0000001011011000001000",
			5 => "0001001010000100000100",
			6 => "0000000000000001001101",
			7 => "0000000000000001001101",
			8 => "0000000000000001001101",
			9 => "0000000000000001001101",
			10 => "0000100010101100001000",
			11 => "0000010110001100000100",
			12 => "0000000000000001001101",
			13 => "0000000000000001001101",
			14 => "0001101011010100000100",
			15 => "0000000000000001001101",
			16 => "0000111001010100000100",
			17 => "0000000000000001001101",
			18 => "0000000000000001001101",
			19 => "0011100010110100100100",
			20 => "0000001011001000010000",
			21 => "0011111111110000000100",
			22 => "0000000000000010110001",
			23 => "0001011100110000001000",
			24 => "0000011000011000000100",
			25 => "0000000000000010110001",
			26 => "0000000000000010110001",
			27 => "0000000000000010110001",
			28 => "0001001000000100001100",
			29 => "0001110110011100000100",
			30 => "0000000000000010110001",
			31 => "0001110001001000000100",
			32 => "0000000000000010110001",
			33 => "0000000000000010110001",
			34 => "0001100000010000000100",
			35 => "0000000000000010110001",
			36 => "0000000000000010110001",
			37 => "0000001101111000001100",
			38 => "0010001111001000001000",
			39 => "0000111100110000000100",
			40 => "0000000000000010110001",
			41 => "0000000000000010110001",
			42 => "0000000000000010110001",
			43 => "0000000000000010110001",
			44 => "0000111100110000100100",
			45 => "0001111001010000010100",
			46 => "0000001110000100001100",
			47 => "0001101101000100000100",
			48 => "0000000000000100011101",
			49 => "0001000111011100000100",
			50 => "0000000000000100011101",
			51 => "0000000000000100011101",
			52 => "0010110011010000000100",
			53 => "0000000000000100011101",
			54 => "0000000000000100011101",
			55 => "0000001011001100001100",
			56 => "0010011101101000001000",
			57 => "0010011100101000000100",
			58 => "0000000000000100011101",
			59 => "0000000000000100011101",
			60 => "0000000000000100011101",
			61 => "0000000000000100011101",
			62 => "0000100011011100001000",
			63 => "0011100011010100000100",
			64 => "0000000000000100011101",
			65 => "0000000000000100011101",
			66 => "0001001111011000000100",
			67 => "0000000000000100011101",
			68 => "0010011010000100000100",
			69 => "0000000000000100011101",
			70 => "0000000000000100011101",
			71 => "0000100011011100100000",
			72 => "0011101001011100010100",
			73 => "0010010101010100001000",
			74 => "0000001110100000000100",
			75 => "0000000000000110011001",
			76 => "0000000000000110011001",
			77 => "0011100010010100000100",
			78 => "0000000000000110011001",
			79 => "0010001001000100000100",
			80 => "0000000000000110011001",
			81 => "0000000000000110011001",
			82 => "0001011100110000000100",
			83 => "0000000000000110011001",
			84 => "0000010110010000000100",
			85 => "0000000000000110011001",
			86 => "0000000000000110011001",
			87 => "0001101101010100010000",
			88 => "0011000111011100000100",
			89 => "0000000000000110011001",
			90 => "0011100110111000000100",
			91 => "0000000000000110011001",
			92 => "0010010011000000000100",
			93 => "0000000000000110011001",
			94 => "0000000000000110011001",
			95 => "0000111100110000001000",
			96 => "0000001001101000000100",
			97 => "0000000000000110011001",
			98 => "0000000000000110011001",
			99 => "0001001111011000000100",
			100 => "0000000000000110011001",
			101 => "0000000000000110011001",
			102 => "0000001110110100100000",
			103 => "0011100101110100011000",
			104 => "0001000101011100001100",
			105 => "0001101101000100000100",
			106 => "0000000000001000001101",
			107 => "0000001011011100000100",
			108 => "0000000000001000001101",
			109 => "0000000000001000001101",
			110 => "0000110011000000001000",
			111 => "0000111101101000000100",
			112 => "0000000000001000001101",
			113 => "0000000000001000001101",
			114 => "0000000000001000001101",
			115 => "0000010110010000000100",
			116 => "0000000000001000001101",
			117 => "0000000000001000001101",
			118 => "0011100101001100010100",
			119 => "0000111000101000001100",
			120 => "0001001000000100001000",
			121 => "0001111000100000000100",
			122 => "0000000000001000001101",
			123 => "0000000000001000001101",
			124 => "0000000000001000001101",
			125 => "0010011010000100000100",
			126 => "0000000000001000001101",
			127 => "0000000000001000001101",
			128 => "0000111001010100000100",
			129 => "0000000000001000001101",
			130 => "0000000000001000001101",
			131 => "0011100010110100100000",
			132 => "0000000011011100010000",
			133 => "0011101101000100000100",
			134 => "0000000000001001111001",
			135 => "0001011001010100001000",
			136 => "0000011000011000000100",
			137 => "0000000000001001111001",
			138 => "0000000000001001111001",
			139 => "0000000000001001111001",
			140 => "0000010000011000001100",
			141 => "0001001001000100000100",
			142 => "0000000000001001111001",
			143 => "0000011001100100000100",
			144 => "0000000000001001111001",
			145 => "0000000000001001111001",
			146 => "0000000000001001111001",
			147 => "0000000011001100000100",
			148 => "0000000000001001111001",
			149 => "0001100000100100001100",
			150 => "0011111011000100000100",
			151 => "0000000000001001111001",
			152 => "0010101001010100000100",
			153 => "0000000000001001111001",
			154 => "0000000000001001111001",
			155 => "0001100101100100000100",
			156 => "0000000000001001111001",
			157 => "0000000000001001111001",
			158 => "0010011101101000101000",
			159 => "0001111001010000010000",
			160 => "0000001110000100001100",
			161 => "0001101101000100000100",
			162 => "1111111000001011100101",
			163 => "0011110110110000000100",
			164 => "0000000000001011100101",
			165 => "0000001000001011100101",
			166 => "1111111000001011100101",
			167 => "0000000011001100010000",
			168 => "0001000101010100000100",
			169 => "0000001000001011100101",
			170 => "0011011010100100001000",
			171 => "0000010111100100000100",
			172 => "0000001000001011100101",
			173 => "0000000000001011100101",
			174 => "0000001000001011100101",
			175 => "0001101011010100000100",
			176 => "1111111000001011100101",
			177 => "0000000000001011100101",
			178 => "0000010000011000001100",
			179 => "0001001100000000001000",
			180 => "0000001011101100000100",
			181 => "0000000000001011100101",
			182 => "0000001000001011100101",
			183 => "1111111000001011100101",
			184 => "1111111000001011100101",
			185 => "0011101100011000101000",
			186 => "0001000101011100010000",
			187 => "0001101111000100000100",
			188 => "0000000000001101101001",
			189 => "0000000101011000001000",
			190 => "0010011100101000000100",
			191 => "0000000000001101101001",
			192 => "0000000000001101101001",
			193 => "0000000000001101101001",
			194 => "0001110001010000010000",
			195 => "0000110011000000001100",
			196 => "0001011111011000001000",
			197 => "0000111100101000000100",
			198 => "0000000000001101101001",
			199 => "0000000000001101101001",
			200 => "0000000000001101101001",
			201 => "1111111000001101101001",
			202 => "0001011100010000000100",
			203 => "0000000000001101101001",
			204 => "0000000000001101101001",
			205 => "0000100010101100001100",
			206 => "0010101011111000001000",
			207 => "0001011000000000000100",
			208 => "0000001000001101101001",
			209 => "0000000000001101101001",
			210 => "0000000000001101101001",
			211 => "0011110011100000001000",
			212 => "0011010110110100000100",
			213 => "0000000000001101101001",
			214 => "1111111000001101101001",
			215 => "0000111001010100000100",
			216 => "0000001000001101101001",
			217 => "0000000000001101101001",
			218 => "0011101001011100010100",
			219 => "0010111011101100001000",
			220 => "0001110011000000000100",
			221 => "1111111000001111001101",
			222 => "0000001000001111001101",
			223 => "0011101001110000000100",
			224 => "1111111000001111001101",
			225 => "0000011000011000000100",
			226 => "0000000000001111001101",
			227 => "1111111000001111001101",
			228 => "0000001101111000011100",
			229 => "0010010101111000011000",
			230 => "0000100011011100001100",
			231 => "0011100001101100001000",
			232 => "0001000101011100000100",
			233 => "0000001000001111001101",
			234 => "0000000000001111001101",
			235 => "0000001000001111001101",
			236 => "0011100110111000000100",
			237 => "1111111000001111001101",
			238 => "0000111100110000000100",
			239 => "0000001000001111001101",
			240 => "0000000000001111001101",
			241 => "1111111000001111001101",
			242 => "1111111000001111001101",
			243 => "0001100100001000101100",
			244 => "0001011010000100001100",
			245 => "0001101101000100000100",
			246 => "0000000000010001001001",
			247 => "0000001100010100000100",
			248 => "0000000000010001001001",
			249 => "0000000000010001001001",
			250 => "0010001111111100010000",
			251 => "0001110001010000001100",
			252 => "0000101011011100001000",
			253 => "0001111100110000000100",
			254 => "0000000000010001001001",
			255 => "0000000000010001001001",
			256 => "0000000000010001001001",
			257 => "0000000000010001001001",
			258 => "0000010111110000001000",
			259 => "0001000110000000000100",
			260 => "0000000000010001001001",
			261 => "0000000000010001001001",
			262 => "0001000011010000000100",
			263 => "0000000000010001001001",
			264 => "0000000000010001001001",
			265 => "0000000011001100000100",
			266 => "0000000000010001001001",
			267 => "0001000111011100001000",
			268 => "0000111000000000000100",
			269 => "0000000000010001001001",
			270 => "0000000000010001001001",
			271 => "0001001001001000000100",
			272 => "0000000000010001001001",
			273 => "0000000000010001001001",
			274 => "0011101100011000101000",
			275 => "0001000101011100010000",
			276 => "0001101101000100000100",
			277 => "0000000000010011001101",
			278 => "0000001110000100000100",
			279 => "0000001000010011001101",
			280 => "0001111101001000000100",
			281 => "0000000000010011001101",
			282 => "0000000000010011001101",
			283 => "0000110011000000001100",
			284 => "0001110110101100000100",
			285 => "0000000000010011001101",
			286 => "0001010101101100000100",
			287 => "0000000000010011001101",
			288 => "0000000000010011001101",
			289 => "0001110001010000000100",
			290 => "1111111000010011001101",
			291 => "0011100010110000000100",
			292 => "0000000000010011001101",
			293 => "0000000000010011001101",
			294 => "0000001101111000011000",
			295 => "0000111100110000001100",
			296 => "0011011110011000001000",
			297 => "0011100111100000000100",
			298 => "0000000000010011001101",
			299 => "0000000000010011001101",
			300 => "0000001000010011001101",
			301 => "0001011001010100000100",
			302 => "0000000000010011001101",
			303 => "0000011101000000000100",
			304 => "0000001000010011001101",
			305 => "0000000000010011001101",
			306 => "1111111000010011001101",
			307 => "0011101100011000100100",
			308 => "0001000101011100011000",
			309 => "0001111100010000001100",
			310 => "0010010111011100001000",
			311 => "0000011001100100000100",
			312 => "0000000000010101100001",
			313 => "0000000000010101100001",
			314 => "0000000000010101100001",
			315 => "0000001110110100001000",
			316 => "0010011101101000000100",
			317 => "0000000000010101100001",
			318 => "0000000000010101100001",
			319 => "0000000000010101100001",
			320 => "0000110011000000001000",
			321 => "0000111101101000000100",
			322 => "0000000000010101100001",
			323 => "0000000000010101100001",
			324 => "0000000000010101100001",
			325 => "0000100010101100010100",
			326 => "0010101011111000010000",
			327 => "0001011000000000001000",
			328 => "0001010011001000000100",
			329 => "0000000000010101100001",
			330 => "0000000000010101100001",
			331 => "0001011100110000000100",
			332 => "0000000000010101100001",
			333 => "0000000000010101100001",
			334 => "0000000000010101100001",
			335 => "0001100000100100001100",
			336 => "0011010110110100000100",
			337 => "0000000000010101100001",
			338 => "0000110011001000000100",
			339 => "0000000000010101100001",
			340 => "0000000000010101100001",
			341 => "0000111001010100000100",
			342 => "0000000000010101100001",
			343 => "0000000000010101100001",
			344 => "0011100011101000101000",
			345 => "0001000011010000001100",
			346 => "0001101101000100000100",
			347 => "0000000000010111001101",
			348 => "0000001100010100000100",
			349 => "0000000000010111001101",
			350 => "0000000000010111001101",
			351 => "0010001001000100011000",
			352 => "0001110001010000010000",
			353 => "0000111001000100000100",
			354 => "0000000000010111001101",
			355 => "0001010101111000000100",
			356 => "0000000000010111001101",
			357 => "0001100100100000000100",
			358 => "0000000000010111001101",
			359 => "0000000000010111001101",
			360 => "0001011000101000000100",
			361 => "0000000000010111001101",
			362 => "0000000000010111001101",
			363 => "0000000000010111001101",
			364 => "0000001101111000001100",
			365 => "0000011101000000001000",
			366 => "0001001100101000000100",
			367 => "0000000000010111001101",
			368 => "0000000000010111001101",
			369 => "0000000000010111001101",
			370 => "0000000000010111001101",
			371 => "0001000101011100100000",
			372 => "0000101001110100010000",
			373 => "0001101101000100000100",
			374 => "0000000000011001100001",
			375 => "0001000111011100000100",
			376 => "0000001000011001100001",
			377 => "0001010011001000000100",
			378 => "0000000000011001100001",
			379 => "0000000000011001100001",
			380 => "0001100000100100001100",
			381 => "0010001001001100000100",
			382 => "0000000000011001100001",
			383 => "0001011111011000000100",
			384 => "0000000000011001100001",
			385 => "1111111000011001100001",
			386 => "0000000000011001100001",
			387 => "0011101100011000011000",
			388 => "0001111100101100010000",
			389 => "0000110011000000001100",
			390 => "0000111101101000001000",
			391 => "0001010101111000000100",
			392 => "0000000000011001100001",
			393 => "0000000000011001100001",
			394 => "0000000000011001100001",
			395 => "0000000000011001100001",
			396 => "0001011100010000000100",
			397 => "0000000000011001100001",
			398 => "0000000000011001100001",
			399 => "0011111011110100001000",
			400 => "0000000010101100000100",
			401 => "0000000000011001100001",
			402 => "0000000000011001100001",
			403 => "0011011010100100000100",
			404 => "1111111000011001100001",
			405 => "0000001011100100000100",
			406 => "0000000000011001100001",
			407 => "0000000000011001100001",
			408 => "0001110001010000101000",
			409 => "0010011001001000011000",
			410 => "0000001110110100010100",
			411 => "0001111100010000001100",
			412 => "0001011100101000001000",
			413 => "0000101101000100000100",
			414 => "0000000000011011101101",
			415 => "0000001000011011101101",
			416 => "1111111000011011101101",
			417 => "0001111101001000000100",
			418 => "0000000000011011101101",
			419 => "0000001000011011101101",
			420 => "1111111000011011101101",
			421 => "0001010101111000001100",
			422 => "0001010110000000000100",
			423 => "0000000000011011101101",
			424 => "0001011101101000000100",
			425 => "0000000000011011101101",
			426 => "0000000000011011101101",
			427 => "1111111000011011101101",
			428 => "0000100011011100001000",
			429 => "0010010101111000000100",
			430 => "0000001000011011101101",
			431 => "0000000000011011101101",
			432 => "0010001111001000010000",
			433 => "0000011001100000001000",
			434 => "0000010111100100000100",
			435 => "0000000000011011101101",
			436 => "1111111000011011101101",
			437 => "0011101100000100000100",
			438 => "0000000000011011101101",
			439 => "0000001000011011101101",
			440 => "0000000011111000000100",
			441 => "0000000000011011101101",
			442 => "1111111000011011101101",
			443 => "0001101101010100111000",
			444 => "0000101011101000010100",
			445 => "0011100010010100001100",
			446 => "0010010101010100001000",
			447 => "0011011101000000000100",
			448 => "0000000000011101110001",
			449 => "0000000000011101110001",
			450 => "0000000000011101110001",
			451 => "0001011001010100000100",
			452 => "0000000000011101110001",
			453 => "0000000000011101110001",
			454 => "0011000111011100010100",
			455 => "0001001001000100001100",
			456 => "0000110011100100001000",
			457 => "0000111111011000000100",
			458 => "0000000000011101110001",
			459 => "0000000000011101110001",
			460 => "0000000000011101110001",
			461 => "0000010111100100000100",
			462 => "0000000000011101110001",
			463 => "0000000000011101110001",
			464 => "0000011000011000001000",
			465 => "0011101100011000000100",
			466 => "0000000000011101110001",
			467 => "0000000000011101110001",
			468 => "0001000110000000000100",
			469 => "0000000000011101110001",
			470 => "0000000000011101110001",
			471 => "0010111011101100000100",
			472 => "0000000000011101110001",
			473 => "0000011101000000000100",
			474 => "0000000000011101110001",
			475 => "0000000000011101110001",
			476 => "0010000101101100100000",
			477 => "0001110110101100010000",
			478 => "0000000001111000001100",
			479 => "0001111000000100000100",
			480 => "0000000000100000000101",
			481 => "0000111101101000000100",
			482 => "0000000000100000000101",
			483 => "0000000000100000000101",
			484 => "0000000000100000000101",
			485 => "0000001101111000001100",
			486 => "0010111011101100000100",
			487 => "0000000000100000000101",
			488 => "0001010011110100000100",
			489 => "0000000000100000000101",
			490 => "0000000000100000000101",
			491 => "0000000000100000000101",
			492 => "0011101100000100100000",
			493 => "0010111011101100001000",
			494 => "0001010011001000000100",
			495 => "0000000000100000000101",
			496 => "0000000000100000000101",
			497 => "0000101011101000001100",
			498 => "0001110001010000000100",
			499 => "0000000000100000000101",
			500 => "0001011100110000000100",
			501 => "0000000000100000000101",
			502 => "0000000000100000000101",
			503 => "0000111100101100000100",
			504 => "0000000000100000000101",
			505 => "0001010000111100000100",
			506 => "0000000000100000000101",
			507 => "0000000000100000000101",
			508 => "0010101111101000000100",
			509 => "0000000000100000000101",
			510 => "0011010101010100000100",
			511 => "0000000000100000000101",
			512 => "0000000000100000000101",
			513 => "0001100100001000110000",
			514 => "0000000011011100100100",
			515 => "0011101110111100010100",
			516 => "0010010101010100001000",
			517 => "0010100101101100000100",
			518 => "0000000000100010010001",
			519 => "0000000000100010010001",
			520 => "0011100010010100000100",
			521 => "0000000000100010010001",
			522 => "0000010111110000000100",
			523 => "0000000000100010010001",
			524 => "0000000000100010010001",
			525 => "0010000000110000001100",
			526 => "0001011100110000001000",
			527 => "0000000101111100000100",
			528 => "0000000000100010010001",
			529 => "0000000000100010010001",
			530 => "0000000000100010010001",
			531 => "0000000000100010010001",
			532 => "0001111011000000000100",
			533 => "0000000000100010010001",
			534 => "0010001010000100000100",
			535 => "0000000000100010010001",
			536 => "0000000000100010010001",
			537 => "0000000011001100000100",
			538 => "0000000000100010010001",
			539 => "0001100000100100001100",
			540 => "0011111011000100000100",
			541 => "0000000000100010010001",
			542 => "0000110011001000000100",
			543 => "0000000000100010010001",
			544 => "0000000000100010010001",
			545 => "0000111001010100000100",
			546 => "0000000000100010010001",
			547 => "0000000000100010010001",
			548 => "0001101101010100110000",
			549 => "0000100011011100100000",
			550 => "0011100101110100011000",
			551 => "0000010111110000010100",
			552 => "0000001110000100001100",
			553 => "0000001110100000000100",
			554 => "0000000000100011111101",
			555 => "0010111010100100000100",
			556 => "0000000000100011111101",
			557 => "0000000000100011111101",
			558 => "0000011001100100000100",
			559 => "0000000000100011111101",
			560 => "0000000000100011111101",
			561 => "0000000000100011111101",
			562 => "0001111011111000000100",
			563 => "0000000000100011111101",
			564 => "0000000000100011111101",
			565 => "0011000111011100000100",
			566 => "0000000000100011111101",
			567 => "0011100110111000000100",
			568 => "0000000000100011111101",
			569 => "0010110101011100000100",
			570 => "0000000000100011111101",
			571 => "0000000000100011111101",
			572 => "0000001101111000000100",
			573 => "0000000000100011111101",
			574 => "0000000000100011111101",
			575 => "0011101100011000100100",
			576 => "0010010101010100001100",
			577 => "0001111000000100000100",
			578 => "0000000000100110001001",
			579 => "0000001100010100000100",
			580 => "0000000000100110001001",
			581 => "0000000000100110001001",
			582 => "0001110001010000001100",
			583 => "0010001010100100000100",
			584 => "0000000000100110001001",
			585 => "0000011000111100000100",
			586 => "0000000000100110001001",
			587 => "0000000000100110001001",
			588 => "0010001001000100001000",
			589 => "0001111011111000000100",
			590 => "0000000000100110001001",
			591 => "0000000000100110001001",
			592 => "0000000000100110001001",
			593 => "0000001101111000100000",
			594 => "0000111100110000001100",
			595 => "0000011001100000001000",
			596 => "0000101000011100000100",
			597 => "0000000000100110001001",
			598 => "0000000000100110001001",
			599 => "0000000000100110001001",
			600 => "0011111011000100010000",
			601 => "0011111001111000001100",
			602 => "0011110000001000001000",
			603 => "0010101011000000000100",
			604 => "0000000000100110001001",
			605 => "0000000000100110001001",
			606 => "0000000000100110001001",
			607 => "0000000000100110001001",
			608 => "0000000000100110001001",
			609 => "0000000000100110001001",
			610 => "0001111001010000011100",
			611 => "0001011101101000010000",
			612 => "0010100101101100000100",
			613 => "0000000000101000101101",
			614 => "0000001110000100001000",
			615 => "0000001110100000000100",
			616 => "0000000000101000101101",
			617 => "0000000000101000101101",
			618 => "0000000000101000101101",
			619 => "0000111001000100000100",
			620 => "0000000000101000101101",
			621 => "0001001010100100000100",
			622 => "0000000000101000101101",
			623 => "0000000000101000101101",
			624 => "0010101111101000011100",
			625 => "0001011100010000010000",
			626 => "0011010101010100001100",
			627 => "0011011110011000001000",
			628 => "0001100100001000000100",
			629 => "0000000000101000101101",
			630 => "0000000000101000101101",
			631 => "0000000000101000101101",
			632 => "0000000000101000101101",
			633 => "0011111000001000001000",
			634 => "0001101000110100000100",
			635 => "0000000000101000101101",
			636 => "0000000000101000101101",
			637 => "0000000000101000101101",
			638 => "0000010111100100001000",
			639 => "0001011010011100000100",
			640 => "0000000000101000101101",
			641 => "0000000000101000101101",
			642 => "0011110111101100010000",
			643 => "0011010101010100001000",
			644 => "0000001011001000000100",
			645 => "0000000000101000101101",
			646 => "0000000000101000101101",
			647 => "0001100110011000000100",
			648 => "0000000000101000101101",
			649 => "0000000000101000101101",
			650 => "0000000000101000101101",
			651 => "0011101100011000101000",
			652 => "0001000101011100010100",
			653 => "0001101101000100000100",
			654 => "1111111000101010111001",
			655 => "0000000001110100001100",
			656 => "0000000000001100000100",
			657 => "0000001000101010111001",
			658 => "0000110011000000000100",
			659 => "0000000000101010111001",
			660 => "0000001000101010111001",
			661 => "1111111000101010111001",
			662 => "0001110001010000001100",
			663 => "0000110011000000001000",
			664 => "0010100011000000000100",
			665 => "0000000000101010111001",
			666 => "0000000000101010111001",
			667 => "1111111000101010111001",
			668 => "0001011001010100000100",
			669 => "0000000000101010111001",
			670 => "1111111000101010111001",
			671 => "0000001101111000011100",
			672 => "0000000011011100000100",
			673 => "0000001000101010111001",
			674 => "0001100100001000001100",
			675 => "0011111101010100001000",
			676 => "0010101011000000000100",
			677 => "0000001000101010111001",
			678 => "1111111000101010111001",
			679 => "1111111000101010111001",
			680 => "0001011001010000001000",
			681 => "0011001010100100000100",
			682 => "0000000000101010111001",
			683 => "0000000000101010111001",
			684 => "0000001000101010111001",
			685 => "1111111000101010111001",
			686 => "0011101010001000111000",
			687 => "0000000011011100011100",
			688 => "0011100101110100011000",
			689 => "0000010111110000010000",
			690 => "0011111111110000000100",
			691 => "0000000000101101001101",
			692 => "0000001110000100000100",
			693 => "0000000000101101001101",
			694 => "0010110101010100000100",
			695 => "0000000000101101001101",
			696 => "0000000000101101001101",
			697 => "0010001001001100000100",
			698 => "0000000000101101001101",
			699 => "1111111000101101001101",
			700 => "0000001000101101001101",
			701 => "0001111100101100010100",
			702 => "0000110011001000001000",
			703 => "0010000101101100000100",
			704 => "0000000000101101001101",
			705 => "0000000000101101001101",
			706 => "0010001001001100001000",
			707 => "0001001000000100000100",
			708 => "0000000000101101001101",
			709 => "0000000000101101001101",
			710 => "1111111000101101001101",
			711 => "0000011000011000000100",
			712 => "0000000000101101001101",
			713 => "0000000000101101001101",
			714 => "0010001111001000001100",
			715 => "0000000000101000000100",
			716 => "0000000000101101001101",
			717 => "0011110111101100000100",
			718 => "0000000000101101001101",
			719 => "0000000000101101001101",
			720 => "0011111011110100000100",
			721 => "0000000000101101001101",
			722 => "0000000000101101001101",
			723 => "0000111100110000110000",
			724 => "0011100011101000100100",
			725 => "0000001011111100100000",
			726 => "0010000101101100010000",
			727 => "0001111000000100000100",
			728 => "0000000000101111101001",
			729 => "0011010011010000001000",
			730 => "0001111100010000000100",
			731 => "0000000000101111101001",
			732 => "0000000000101111101001",
			733 => "0000000000101111101001",
			734 => "0010111110011000001000",
			735 => "0011001011101100000100",
			736 => "0000000000101111101001",
			737 => "0000000000101111101001",
			738 => "0011101001011100000100",
			739 => "0000000000101111101001",
			740 => "0000000000101111101001",
			741 => "0000000000101111101001",
			742 => "0010001111001000001000",
			743 => "0000001011001100000100",
			744 => "0000000000101111101001",
			745 => "0000000000101111101001",
			746 => "0000000000101111101001",
			747 => "0010010101101100010000",
			748 => "0000001010010100001000",
			749 => "0000000111101100000100",
			750 => "0000000000101111101001",
			751 => "1111111000101111101001",
			752 => "0000000101101000000100",
			753 => "0000000000101111101001",
			754 => "0000000000101111101001",
			755 => "0011100011101000001000",
			756 => "0001011001010000000100",
			757 => "0000000000101111101001",
			758 => "0000000000101111101001",
			759 => "0000000110111100000100",
			760 => "0000000000101111101001",
			761 => "0000000000101111101001",
			762 => "0011101100011000101100",
			763 => "0001000101011100010100",
			764 => "0000010111100100010000",
			765 => "0001101101000100000100",
			766 => "0000000000110001110101",
			767 => "0000001110000100000100",
			768 => "0000001000110001110101",
			769 => "0001111101001000000100",
			770 => "0000000000110001110101",
			771 => "0000000000110001110101",
			772 => "0000000000110001110101",
			773 => "0000110011000000001100",
			774 => "0001110110101100000100",
			775 => "0000000000110001110101",
			776 => "0001010101101100000100",
			777 => "0000000000110001110101",
			778 => "0000000000110001110101",
			779 => "0001110001010000000100",
			780 => "1111111000110001110101",
			781 => "0011100010110000000100",
			782 => "0000000000110001110101",
			783 => "0000000000110001110101",
			784 => "0000001101111000011000",
			785 => "0001011111011000000100",
			786 => "0000001000110001110101",
			787 => "0001011000000100000100",
			788 => "0000000000110001110101",
			789 => "0000100011011100000100",
			790 => "0000001000110001110101",
			791 => "0001101100111100001000",
			792 => "0011000111011100000100",
			793 => "1111111000110001110101",
			794 => "0000000000110001110101",
			795 => "0000000000110001110101",
			796 => "1111111000110001110101",
			797 => "0001100010001000001100",
			798 => "0010010111011100001000",
			799 => "0011011101000000000100",
			800 => "0000000000110011100001",
			801 => "0000000000110011100001",
			802 => "1111111000110011100001",
			803 => "0011000110001100000100",
			804 => "0000001000110011100001",
			805 => "0001010011000000001000",
			806 => "0010111011101100000100",
			807 => "0000000000110011100001",
			808 => "0000001000110011100001",
			809 => "0001110001010000001100",
			810 => "0000000111000100001000",
			811 => "0010011001001000000100",
			812 => "0000000000110011100001",
			813 => "1111111000110011100001",
			814 => "1111111000110011100001",
			815 => "0000101011100000001000",
			816 => "0001011001010000000100",
			817 => "0000001000110011100001",
			818 => "0000000000110011100001",
			819 => "0000010111100100000100",
			820 => "0000000000110011100001",
			821 => "0010101001010100000100",
			822 => "0000001000110011100001",
			823 => "0000000000110011100001",
			824 => "0001101101010101000000",
			825 => "0000001110110100101000",
			826 => "0011101110111100011100",
			827 => "0010010101010100001100",
			828 => "0010110110110100000100",
			829 => "0000000000110101110101",
			830 => "0011100010111000000100",
			831 => "0000000000110101110101",
			832 => "0000000000110101110101",
			833 => "0011010110110100001000",
			834 => "0010001001001100000100",
			835 => "0000000000110101110101",
			836 => "0000000000110101110101",
			837 => "0010000011010000000100",
			838 => "0000000000110101110101",
			839 => "1111111000110101110101",
			840 => "0010111110011000000100",
			841 => "0000000000110101110101",
			842 => "0001011001010000000100",
			843 => "0000001000110101110101",
			844 => "0000000000110101110101",
			845 => "0000110011000100010000",
			846 => "0011101100000100001100",
			847 => "0000010000011000001000",
			848 => "0001000101111000000100",
			849 => "0000000000110101110101",
			850 => "0000000000110101110101",
			851 => "1111111000110101110101",
			852 => "0000000000110101110101",
			853 => "0000110001001000000100",
			854 => "0000000000110101110101",
			855 => "0000000000110101110101",
			856 => "0010111011101100000100",
			857 => "0000000000110101110101",
			858 => "0000011101000000000100",
			859 => "0000001000110101110101",
			860 => "0000000000110101110101",
			861 => "0001100100001000111100",
			862 => "0000000011011100101000",
			863 => "0011101110111100011000",
			864 => "0010010101010100001000",
			865 => "0010100101101100000100",
			866 => "0000000000111000011001",
			867 => "0000000000111000011001",
			868 => "0011101001011100001100",
			869 => "0000011000111100000100",
			870 => "0000000000111000011001",
			871 => "0010000011010000000100",
			872 => "0000000000111000011001",
			873 => "0000000000111000011001",
			874 => "0000000000111000011001",
			875 => "0010000000110000001100",
			876 => "0001011100110000001000",
			877 => "0000000101111100000100",
			878 => "0000000000111000011001",
			879 => "0000000000111000011001",
			880 => "0000000000111000011001",
			881 => "0000000000111000011001",
			882 => "0000010000011000001000",
			883 => "0011101100011000000100",
			884 => "0000000000111000011001",
			885 => "0000000000111000011001",
			886 => "0010001111111100001000",
			887 => "0001111101001000000100",
			888 => "0000000000111000011001",
			889 => "0000000000111000011001",
			890 => "1111111000111000011001",
			891 => "0000000011001100000100",
			892 => "0000000000111000011001",
			893 => "0001100000100100001100",
			894 => "0011111011000100000100",
			895 => "0000000000111000011001",
			896 => "0000110011001000000100",
			897 => "0000000000111000011001",
			898 => "1111111000111000011001",
			899 => "0000111001010100000100",
			900 => "0000000000111000011001",
			901 => "0000000000111000011001",
			902 => "0001100010001000001100",
			903 => "0010010101010100001000",
			904 => "0001101110010100000100",
			905 => "1111111000111010011101",
			906 => "0000001000111010011101",
			907 => "1111111000111010011101",
			908 => "0000000011001100100100",
			909 => "0010010101111000100000",
			910 => "0011100010110000010000",
			911 => "0000011000011000001100",
			912 => "0000000110001000001000",
			913 => "0000001011000100000100",
			914 => "0000001000111010011101",
			915 => "0000001000111010011101",
			916 => "1111111000111010011101",
			917 => "1111111000111010011101",
			918 => "0011000111011100001100",
			919 => "0000100011011100001000",
			920 => "0001110100101100000100",
			921 => "0000001000111010011101",
			922 => "0000001000111010011101",
			923 => "0000000000111010011101",
			924 => "0000001000111010011101",
			925 => "1111111000111010011101",
			926 => "0001101011010100001100",
			927 => "0011010110110100001000",
			928 => "0000111001010100000100",
			929 => "1111111000111010011101",
			930 => "0000001000111010011101",
			931 => "1111111000111010011101",
			932 => "0010011001001000000100",
			933 => "0000001000111010011101",
			934 => "1111111000111010011101",
			935 => "0011101010001001000000",
			936 => "0000100101011000100100",
			937 => "0011101110111100011000",
			938 => "0010010101010100001100",
			939 => "0011011101000000000100",
			940 => "0000000000111101000001",
			941 => "0000111110011000000100",
			942 => "0000000000111101000001",
			943 => "0000000000111101000001",
			944 => "0011010110110100000100",
			945 => "0000000000111101000001",
			946 => "0010000011010000000100",
			947 => "0000000000111101000001",
			948 => "0000000000111101000001",
			949 => "0001011001010000001000",
			950 => "0001101111010100000100",
			951 => "0000000000111101000001",
			952 => "0000000000111101000001",
			953 => "0000000000111101000001",
			954 => "0001001001000100000100",
			955 => "0000000000111101000001",
			956 => "0001100000010000010000",
			957 => "0010000101101100001100",
			958 => "0001000101111000001000",
			959 => "0010001001001100000100",
			960 => "0000000000111101000001",
			961 => "0000000000111101000001",
			962 => "0000000000111101000001",
			963 => "0000000000111101000001",
			964 => "0010011101101000000100",
			965 => "0000000000111101000001",
			966 => "0000000000111101000001",
			967 => "0010001111001000001100",
			968 => "0000000110101000000100",
			969 => "0000000000111101000001",
			970 => "0011110011100000000100",
			971 => "0000000000111101000001",
			972 => "0000000000111101000001",
			973 => "0011111011110100000100",
			974 => "0000000000111101000001",
			975 => "0000000000111101000001",
			976 => "0011101101100100110000",
			977 => "0001011100101000001000",
			978 => "0000001110100000000100",
			979 => "0000000000111111100101",
			980 => "0000000000111111100101",
			981 => "0001111111101000100000",
			982 => "0011101111010100011000",
			983 => "0001011101101000010000",
			984 => "0001010101101100001000",
			985 => "0001001011101100000100",
			986 => "0000000000111111100101",
			987 => "0000000000111111100101",
			988 => "0001001011101100000100",
			989 => "0000000000111111100101",
			990 => "0000000000111111100101",
			991 => "0001000011010000000100",
			992 => "0000000000111111100101",
			993 => "0000000000111111100101",
			994 => "0001001010000100000100",
			995 => "0000000000111111100101",
			996 => "0000000000111111100101",
			997 => "0001000110000000000100",
			998 => "0000000000111111100101",
			999 => "0000000000111111100101",
			1000 => "0000000011001100001100",
			1001 => "0001011000000000000100",
			1002 => "0000000000111111100101",
			1003 => "0001011101001000000100",
			1004 => "0000000000111111100101",
			1005 => "0000000000111111100101",
			1006 => "0001100000100100010000",
			1007 => "0000111111101000001000",
			1008 => "0000110011001000000100",
			1009 => "0000000000111111100101",
			1010 => "0000000000111111100101",
			1011 => "0010101001011000000100",
			1012 => "0000000000111111100101",
			1013 => "0000000000111111100101",
			1014 => "0000111001010100000100",
			1015 => "0000000000111111100101",
			1016 => "0000000000111111100101",
			1017 => "0011101100011000100000",
			1018 => "0000011000011000011100",
			1019 => "0001011100010000011000",
			1020 => "0001111100010000001100",
			1021 => "0001011100101000001000",
			1022 => "0010101111111100000100",
			1023 => "0000000001000001100001",
			1024 => "0000000001000001100001",
			1025 => "0000000001000001100001",
			1026 => "0000001110110100001000",
			1027 => "0001100010001000000100",
			1028 => "0000000001000001100001",
			1029 => "0000001001000001100001",
			1030 => "0000000001000001100001",
			1031 => "0000000001000001100001",
			1032 => "1111111001000001100001",
			1033 => "0000001101111000011100",
			1034 => "0000110011100100000100",
			1035 => "0000001001000001100001",
			1036 => "0010000101101100001000",
			1037 => "0011110000100100000100",
			1038 => "0000001001000001100001",
			1039 => "0000000001000001100001",
			1040 => "0011011010100100000100",
			1041 => "0000000001000001100001",
			1042 => "0000100010101100001000",
			1043 => "0010100100101100000100",
			1044 => "0000001001000001100001",
			1045 => "0000000001000001100001",
			1046 => "0000000001000001100001",
			1047 => "0000000001000001100001",
			1048 => "0010011101101000111100",
			1049 => "0001111100010000001100",
			1050 => "0010010101010100001000",
			1051 => "0001111000000100000100",
			1052 => "1111111001000011101101",
			1053 => "0000001001000011101101",
			1054 => "1111111001000011101101",
			1055 => "0000100011011100010000",
			1056 => "0011100010010100000100",
			1057 => "0000000001000011101101",
			1058 => "0010001001000100001000",
			1059 => "0010001111111100000100",
			1060 => "0000001001000011101101",
			1061 => "0000001001000011101101",
			1062 => "0000001001000011101101",
			1063 => "0001101101010100011000",
			1064 => "0010011001000100010000",
			1065 => "0000110011001000001000",
			1066 => "0011001010100100000100",
			1067 => "0000000001000011101101",
			1068 => "1111111001000011101101",
			1069 => "0001100000001100000100",
			1070 => "1111111001000011101101",
			1071 => "1111111001000011101101",
			1072 => "0001100001111000000100",
			1073 => "1111111001000011101101",
			1074 => "0000001001000011101101",
			1075 => "0001111011111000000100",
			1076 => "0000010001000011101101",
			1077 => "0000001001000011101101",
			1078 => "0010001001000100001000",
			1079 => "0011100011010100000100",
			1080 => "1111111001000011101101",
			1081 => "0000001001000011101101",
			1082 => "1111111001000011101101",
			1083 => "0010000101101100100100",
			1084 => "0001101101000100000100",
			1085 => "0000000001000110000001",
			1086 => "0000001101111000011100",
			1087 => "0000010111100100010000",
			1088 => "0001010011110100001100",
			1089 => "0010000011010000001000",
			1090 => "0011010110110100000100",
			1091 => "0000000001000110000001",
			1092 => "0000000001000110000001",
			1093 => "0000000001000110000001",
			1094 => "0000000001000110000001",
			1095 => "0010000101011100000100",
			1096 => "0000000001000110000001",
			1097 => "0001011000000000000100",
			1098 => "0000000001000110000001",
			1099 => "0000000001000110000001",
			1100 => "0000000001000110000001",
			1101 => "0000110011100100001000",
			1102 => "0011101111010100000100",
			1103 => "0000000001000110000001",
			1104 => "0000000001000110000001",
			1105 => "0000000011011100001000",
			1106 => "0001011100110000000100",
			1107 => "0000000001000110000001",
			1108 => "0000000001000110000001",
			1109 => "0001001111011000001100",
			1110 => "0001110011000100001000",
			1111 => "0011010101010100000100",
			1112 => "0000000001000110000001",
			1113 => "0000000001000110000001",
			1114 => "0000000001000110000001",
			1115 => "0011010101011100001000",
			1116 => "0001001100010000000100",
			1117 => "0000000001000110000001",
			1118 => "0000000001000110000001",
			1119 => "0000000001000110000001",
			1120 => "0011101111010100101000",
			1121 => "0000011000011000100100",
			1122 => "0001001101101000011100",
			1123 => "0001111100010000010000",
			1124 => "0001011100101000001100",
			1125 => "0001111000000100000100",
			1126 => "0000000001001000010101",
			1127 => "0001011011101100000100",
			1128 => "0000000001001000010101",
			1129 => "0000000001001000010101",
			1130 => "0000000001001000010101",
			1131 => "0000001010101000001000",
			1132 => "0001100010001000000100",
			1133 => "0000000001001000010101",
			1134 => "0000000001001000010101",
			1135 => "0000000001001000010101",
			1136 => "0001010110101100000100",
			1137 => "0000000001001000010101",
			1138 => "0000000001001000010101",
			1139 => "0000000001001000010101",
			1140 => "0000001101111000100000",
			1141 => "0010101111101000010000",
			1142 => "0001011100010000001100",
			1143 => "0001011000000100001000",
			1144 => "0000101011100000000100",
			1145 => "0000000001001000010101",
			1146 => "0000000001001000010101",
			1147 => "0000001001001000010101",
			1148 => "0000000001001000010101",
			1149 => "0001011001010000000100",
			1150 => "0000000001001000010101",
			1151 => "0011100110111000000100",
			1152 => "0000000001001000010101",
			1153 => "0001110011110100000100",
			1154 => "0000000001001000010101",
			1155 => "0000000001001000010101",
			1156 => "0000000001001000010101",
			1157 => "0011100011101000111000",
			1158 => "0011111101010100110000",
			1159 => "0011101100011000101000",
			1160 => "0001000101011100010000",
			1161 => "0001101101000100000100",
			1162 => "1111111001001010110001",
			1163 => "0000000000001100000100",
			1164 => "0000001001001010110001",
			1165 => "0001111100110000000100",
			1166 => "1111111001001010110001",
			1167 => "0000000001001010110001",
			1168 => "0001111111101000010000",
			1169 => "0001010101111000001000",
			1170 => "0000111100101000000100",
			1171 => "0000000001001010110001",
			1172 => "0000000001001010110001",
			1173 => "0000110110000000000100",
			1174 => "0000000001001010110001",
			1175 => "1111111001001010110001",
			1176 => "0001011001010000000100",
			1177 => "0000000001001010110001",
			1178 => "0000000001001010110001",
			1179 => "0001011000101000000100",
			1180 => "0000001001001010110001",
			1181 => "0000000001001010110001",
			1182 => "0001010101111000000100",
			1183 => "0000000001001010110001",
			1184 => "1111111001001010110001",
			1185 => "0000011101000000010000",
			1186 => "0011110011100000001100",
			1187 => "0000000110101000000100",
			1188 => "0000000001001010110001",
			1189 => "0011101110010000000100",
			1190 => "0000000001001010110001",
			1191 => "1111111001001010110001",
			1192 => "0000001001001010110001",
			1193 => "0000111100010000000100",
			1194 => "0000000001001010110001",
			1195 => "1111111001001010110001",
			1196 => "0001100100001001000100",
			1197 => "0000000011011100101100",
			1198 => "0011101110111100100000",
			1199 => "0010010101010100001000",
			1200 => "0010100101101100000100",
			1201 => "0000000001001101110101",
			1202 => "0000000001001101110101",
			1203 => "0001111111101000010000",
			1204 => "0010000011010000001000",
			1205 => "0000011000111100000100",
			1206 => "0000000001001101110101",
			1207 => "0000000001001101110101",
			1208 => "0011010110110100000100",
			1209 => "0000000001001101110101",
			1210 => "0000000001001101110101",
			1211 => "0011101001011100000100",
			1212 => "0000000001001101110101",
			1213 => "0000000001001101110101",
			1214 => "0010010110000000000100",
			1215 => "0000000001001101110101",
			1216 => "0010000000110000000100",
			1217 => "0000000001001101110101",
			1218 => "0000000001001101110101",
			1219 => "0000010000011000001000",
			1220 => "0011101100011000000100",
			1221 => "0000000001001101110101",
			1222 => "0000000001001101110101",
			1223 => "0011100010110100001100",
			1224 => "0010000101011100001000",
			1225 => "0010001001001100000100",
			1226 => "0000000001001101110101",
			1227 => "0000000001001101110101",
			1228 => "0000000001001101110101",
			1229 => "0000000001001101110101",
			1230 => "0011111011000100000100",
			1231 => "0000000001001101110101",
			1232 => "0001101101010100001100",
			1233 => "0001110011000100000100",
			1234 => "0000000001001101110101",
			1235 => "0011100100110000000100",
			1236 => "0000000001001101110101",
			1237 => "0000000001001101110101",
			1238 => "0001111100101100001000",
			1239 => "0000001011001100000100",
			1240 => "0000000001001101110101",
			1241 => "0000000001001101110101",
			1242 => "0000111100110000000100",
			1243 => "0000000001001101110101",
			1244 => "0000000001001101110101",
			1245 => "0011100011101000111100",
			1246 => "0000001011111100111000",
			1247 => "0010001001000100011100",
			1248 => "0011101101000100010000",
			1249 => "0010010101010100001000",
			1250 => "0000001111010100000100",
			1251 => "0000000001010001000001",
			1252 => "0000000001010001000001",
			1253 => "0011010110110100000100",
			1254 => "0000000001010001000001",
			1255 => "1111111001010001000001",
			1256 => "0000111111101000001000",
			1257 => "0001111101001000000100",
			1258 => "0000000001010001000001",
			1259 => "0000001001010001000001",
			1260 => "0000000001010001000001",
			1261 => "0001000011010000001000",
			1262 => "0000101000010100000100",
			1263 => "0000000001010001000001",
			1264 => "0000000001010001000001",
			1265 => "0001001010000100001100",
			1266 => "0001010011000000001000",
			1267 => "0001011001000100000100",
			1268 => "0000000001010001000001",
			1269 => "0000000001010001000001",
			1270 => "1111111001010001000001",
			1271 => "0001001111011000000100",
			1272 => "0000000001010001000001",
			1273 => "0000000001010001000001",
			1274 => "1111111001010001000001",
			1275 => "0000111100110000010000",
			1276 => "0010001111001000001000",
			1277 => "0000001011001100000100",
			1278 => "0000001001010001000001",
			1279 => "0000000001010001000001",
			1280 => "0011100101000000000100",
			1281 => "0000000001010001000001",
			1282 => "0000000001010001000001",
			1283 => "0011100001111000011000",
			1284 => "0000111000101000001100",
			1285 => "0000111001010100001000",
			1286 => "0011100101000000000100",
			1287 => "0000000001010001000001",
			1288 => "0000000001010001000001",
			1289 => "1111111001010001000001",
			1290 => "0011100100000100001000",
			1291 => "0000100110101000000100",
			1292 => "0000001001010001000001",
			1293 => "0000000001010001000001",
			1294 => "0000000001010001000001",
			1295 => "1111111001010001000001",
			1296 => "0001101101010101000000",
			1297 => "0011111011000100110100",
			1298 => "0001100100001000110000",
			1299 => "0000000011011100011100",
			1300 => "0011101001011100010000",
			1301 => "0010010101010100001000",
			1302 => "0010100101101100000100",
			1303 => "0000000001010011001111",
			1304 => "0000000001010011001111",
			1305 => "0000011000111100000100",
			1306 => "0000000001010011001111",
			1307 => "0000000001010011001111",
			1308 => "0001011100110000000100",
			1309 => "0000000001010011001111",
			1310 => "0010001010000100000100",
			1311 => "0000000001010011001111",
			1312 => "0000000001010011001111",
			1313 => "0000010000011000001000",
			1314 => "0011100111001000000100",
			1315 => "0000000001010011001111",
			1316 => "0000000001010011001111",
			1317 => "0010001111111100001000",
			1318 => "0011100111001000000100",
			1319 => "0000000001010011001111",
			1320 => "0000000001010011001111",
			1321 => "0000000001010011001111",
			1322 => "0000000001010011001111",
			1323 => "0001110011000100000100",
			1324 => "0000000001010011001111",
			1325 => "0011100100110000000100",
			1326 => "0000000001010011001111",
			1327 => "0000000001010011001111",
			1328 => "0000001101111000000100",
			1329 => "0000000001010011001111",
			1330 => "0000000001010011001111",
			1331 => "0011101100011000010100",
			1332 => "0001000101011100010000",
			1333 => "0001111100010000000100",
			1334 => "0000000001010100011001",
			1335 => "0000001110110100001000",
			1336 => "0000010111100100000100",
			1337 => "0000000001010100011001",
			1338 => "0000000001010100011001",
			1339 => "0000000001010100011001",
			1340 => "0000000001010100011001",
			1341 => "0000100010101100001000",
			1342 => "0000010110001100000100",
			1343 => "0000000001010100011001",
			1344 => "0000000001010100011001",
			1345 => "0001101011010100000100",
			1346 => "0000000001010100011001",
			1347 => "0000111001010100000100",
			1348 => "0000000001010100011001",
			1349 => "0000000001010100011001",
			1350 => "0011100010110100011100",
			1351 => "0000000011011100010000",
			1352 => "0001100010001000000100",
			1353 => "0000000001010101111101",
			1354 => "0001011001010100001000",
			1355 => "0000011000011000000100",
			1356 => "0000000001010101111101",
			1357 => "0000000001010101111101",
			1358 => "0000000001010101111101",
			1359 => "0011110100100000001000",
			1360 => "0001111011000000000100",
			1361 => "0000000001010101111101",
			1362 => "0000000001010101111101",
			1363 => "0000000001010101111101",
			1364 => "0000000011001100000100",
			1365 => "0000000001010101111101",
			1366 => "0001100000100100001100",
			1367 => "0011111011000100000100",
			1368 => "0000000001010101111101",
			1369 => "0010101001010100000100",
			1370 => "0000000001010101111101",
			1371 => "0000000001010101111101",
			1372 => "0001100101100100000100",
			1373 => "0000000001010101111101",
			1374 => "0000000001010101111101",
			1375 => "0011101100011000100000",
			1376 => "0001000101011100010000",
			1377 => "0001101111000100000100",
			1378 => "0000000001010111110001",
			1379 => "0000000101011000001000",
			1380 => "0010000101011100000100",
			1381 => "0000000001010111110001",
			1382 => "0000000001010111110001",
			1383 => "0000000001010111110001",
			1384 => "0001110001010000001000",
			1385 => "0001011010000100000100",
			1386 => "0000000001010111110001",
			1387 => "1111111001010111110001",
			1388 => "0001011100010000000100",
			1389 => "0000000001010111110001",
			1390 => "0000000001010111110001",
			1391 => "0000100010101100001100",
			1392 => "0010101011111000001000",
			1393 => "0001011000000000000100",
			1394 => "0000001001010111110001",
			1395 => "0000000001010111110001",
			1396 => "0000000001010111110001",
			1397 => "0011110011100000001000",
			1398 => "0011010110110100000100",
			1399 => "0000000001010111110001",
			1400 => "1111111001010111110001",
			1401 => "0000111001010100000100",
			1402 => "0000001001010111110001",
			1403 => "0000000001010111110001",
			1404 => "0000100011011100100000",
			1405 => "0011101001011100010100",
			1406 => "0010010101010100001000",
			1407 => "0000001110100000000100",
			1408 => "0000000001011001101101",
			1409 => "0000000001011001101101",
			1410 => "0011100010010100000100",
			1411 => "0000000001011001101101",
			1412 => "0010001001000100000100",
			1413 => "0000000001011001101101",
			1414 => "0000000001011001101101",
			1415 => "0001011100110000000100",
			1416 => "0000000001011001101101",
			1417 => "0000010110010000000100",
			1418 => "0000000001011001101101",
			1419 => "0000000001011001101101",
			1420 => "0001101101010100010000",
			1421 => "0011000111011100000100",
			1422 => "0000000001011001101101",
			1423 => "0011100110111000000100",
			1424 => "0000000001011001101101",
			1425 => "0010010011000000000100",
			1426 => "0000000001011001101101",
			1427 => "0000000001011001101101",
			1428 => "0000111100110000001000",
			1429 => "0000001001101000000100",
			1430 => "0000000001011001101101",
			1431 => "0000000001011001101101",
			1432 => "0001001111011000000100",
			1433 => "0000000001011001101101",
			1434 => "0000000001011001101101",
			1435 => "0010010110000000101000",
			1436 => "0001110001010000011000",
			1437 => "0001110110101100001100",
			1438 => "0011101111000000000100",
			1439 => "1100111001011011100001",
			1440 => "0000000100111100000100",
			1441 => "1110001001011011100001",
			1442 => "1100111001011011100001",
			1443 => "0000001011001000000100",
			1444 => "1110111001011011100001",
			1445 => "0000000110101000000100",
			1446 => "1101001001011011100001",
			1447 => "1100111001011011100001",
			1448 => "0000100111011000000100",
			1449 => "1110111001011011100001",
			1450 => "0000001111001100001000",
			1451 => "0001001100101000000100",
			1452 => "1101110001011011100001",
			1453 => "1101001001011011100001",
			1454 => "1100111001011011100001",
			1455 => "0010011101101000001000",
			1456 => "0001111000101000000100",
			1457 => "1100111001011011100001",
			1458 => "1101100001011011100001",
			1459 => "0010001001000100001000",
			1460 => "0001100110110000000100",
			1461 => "1100111001011011100001",
			1462 => "1101010001011011100001",
			1463 => "1100111001011011100001",
			1464 => "0001011100000000101000",
			1465 => "0000101001110100011000",
			1466 => "0001100010001000001100",
			1467 => "0001011100101000001000",
			1468 => "0010101111111100000100",
			1469 => "0000000001011101100101",
			1470 => "0000000001011101100101",
			1471 => "0000000001011101100101",
			1472 => "0001111011111000001000",
			1473 => "0001111100010000000100",
			1474 => "0000000001011101100101",
			1475 => "0000000001011101100101",
			1476 => "0000000001011101100101",
			1477 => "0000001010010100001000",
			1478 => "0000110011100100000100",
			1479 => "0000000001011101100101",
			1480 => "0000000001011101100101",
			1481 => "0000001110110000000100",
			1482 => "0000000001011101100101",
			1483 => "0000000001011101100101",
			1484 => "0001011001010000010000",
			1485 => "0011110000001000001000",
			1486 => "0001111111101000000100",
			1487 => "0000000001011101100101",
			1488 => "0000000001011101100101",
			1489 => "0010011001000100000100",
			1490 => "0000000001011101100101",
			1491 => "0000000001011101100101",
			1492 => "0011110101111100000100",
			1493 => "0000000001011101100101",
			1494 => "0011000101011100000100",
			1495 => "0000000001011101100101",
			1496 => "0000000001011101100101",
			1497 => "0010000101101100011000",
			1498 => "0001111001010000001100",
			1499 => "0000001110000100001000",
			1500 => "0001101101000100000100",
			1501 => "0000000001011111010001",
			1502 => "0000000001011111010001",
			1503 => "0000000001011111010001",
			1504 => "0000001101111000001000",
			1505 => "0010101011111000000100",
			1506 => "0000000001011111010001",
			1507 => "0000000001011111010001",
			1508 => "0000000001011111010001",
			1509 => "0000000011001100011000",
			1510 => "0001100100001000010100",
			1511 => "0000101011101000010000",
			1512 => "0011100101110100001100",
			1513 => "0010110101010100000100",
			1514 => "0000000001011111010001",
			1515 => "0010110101011100000100",
			1516 => "0000000001011111010001",
			1517 => "0000000001011111010001",
			1518 => "0000000001011111010001",
			1519 => "0000000001011111010001",
			1520 => "0000000001011111010001",
			1521 => "0000110011001000000100",
			1522 => "0000000001011111010001",
			1523 => "0000000001011111010001",
			1524 => "0001100101110100001100",
			1525 => "0010010101010100001000",
			1526 => "0001100001111100000100",
			1527 => "1111111001100000110101",
			1528 => "0000001001100000110101",
			1529 => "1111111001100000110101",
			1530 => "0000100011011100010100",
			1531 => "0001010001010000010000",
			1532 => "0010001001000100001100",
			1533 => "0010001111111100001000",
			1534 => "0011011011101100000100",
			1535 => "0000001001100000110101",
			1536 => "0000001001100000110101",
			1537 => "0000010001100000110101",
			1538 => "0000001001100000110101",
			1539 => "1111111001100000110101",
			1540 => "0001100100001000000100",
			1541 => "1111111001100000110101",
			1542 => "0000001101111000001100",
			1543 => "0010001111001000001000",
			1544 => "0010111011101100000100",
			1545 => "0000000001100000110101",
			1546 => "0000010001100000110101",
			1547 => "0000000001100000110101",
			1548 => "1111111001100000110101",
			1549 => "0010011101101000101000",
			1550 => "0001111101001000001100",
			1551 => "0011101111000000000100",
			1552 => "1111111001100010101001",
			1553 => "0000100000001100000100",
			1554 => "0000010001100010101001",
			1555 => "1111111001100010101001",
			1556 => "0000000000101000010100",
			1557 => "0001011101001000010000",
			1558 => "0000111100110000001100",
			1559 => "0000001001110100001000",
			1560 => "0010001001000100000100",
			1561 => "0000010001100010101001",
			1562 => "0000010001100010101001",
			1563 => "0000011001100010101001",
			1564 => "0000001001100010101001",
			1565 => "0000001001100010101001",
			1566 => "0011110011100000000100",
			1567 => "1111111001100010101001",
			1568 => "0000001001100010101001",
			1569 => "0000010000011000001000",
			1570 => "0000000100111100000100",
			1571 => "1111111001100010101001",
			1572 => "0000001001100010101001",
			1573 => "0010110101011100001000",
			1574 => "0001111100101100000100",
			1575 => "1111111001100010101001",
			1576 => "0000001001100010101001",
			1577 => "1111111001100010101001",
			1578 => "0001000101011100011100",
			1579 => "0000101001110100010000",
			1580 => "0001101101000100000100",
			1581 => "0000000001100100110101",
			1582 => "0001000111011100000100",
			1583 => "0000001001100100110101",
			1584 => "0001010011001000000100",
			1585 => "0000000001100100110101",
			1586 => "0000000001100100110101",
			1587 => "0011110011100000001000",
			1588 => "0010001001001100000100",
			1589 => "0000000001100100110101",
			1590 => "0000000001100100110101",
			1591 => "0000000001100100110101",
			1592 => "0011101100011000011000",
			1593 => "0001111111101000010000",
			1594 => "0000110011000000001100",
			1595 => "0000111101101000001000",
			1596 => "0001010101111000000100",
			1597 => "0000000001100100110101",
			1598 => "0000000001100100110101",
			1599 => "0000000001100100110101",
			1600 => "0000000001100100110101",
			1601 => "0001011001010100000100",
			1602 => "0000000001100100110101",
			1603 => "0000000001100100110101",
			1604 => "0011111011110100001000",
			1605 => "0000000010101100000100",
			1606 => "0000000001100100110101",
			1607 => "0000000001100100110101",
			1608 => "0011011010100100000100",
			1609 => "0000000001100100110101",
			1610 => "0000011101000000000100",
			1611 => "0000000001100100110101",
			1612 => "0000000001100100110101",
			1613 => "0011101010001000110000",
			1614 => "0000000011011100100000",
			1615 => "0011101001011100010100",
			1616 => "0001011101101000001100",
			1617 => "0001010101011100000100",
			1618 => "0000000001100110111001",
			1619 => "0011101110010100000100",
			1620 => "0000000001100110111001",
			1621 => "0000000001100110111001",
			1622 => "0001000011010000000100",
			1623 => "0000000001100110111001",
			1624 => "0000000001100110111001",
			1625 => "0001011100010000001000",
			1626 => "0010111110011000000100",
			1627 => "0000000001100110111001",
			1628 => "0000000001100110111001",
			1629 => "0000000001100110111001",
			1630 => "0001001001000100000100",
			1631 => "1111111001100110111001",
			1632 => "0000000011111000001000",
			1633 => "0001100100011100000100",
			1634 => "0000000001100110111001",
			1635 => "0000000001100110111001",
			1636 => "0000000001100110111001",
			1637 => "0010001111001000001100",
			1638 => "0010111011101100000100",
			1639 => "0000000001100110111001",
			1640 => "0000111001010100000100",
			1641 => "0000001001100110111001",
			1642 => "0000000001100110111001",
			1643 => "0011111011110100000100",
			1644 => "0000000001100110111001",
			1645 => "0000000001100110111001",
			1646 => "0001100100001000101000",
			1647 => "0000101011101000011100",
			1648 => "0011100101110100011000",
			1649 => "0010010101010100001000",
			1650 => "0011100101110000000100",
			1651 => "0000000001101000100101",
			1652 => "0000001001101000100101",
			1653 => "0011100010010100000100",
			1654 => "1111111001101000100101",
			1655 => "0000111111011000000100",
			1656 => "0000001001101000100101",
			1657 => "0000010111100100000100",
			1658 => "0000000001101000100101",
			1659 => "1111111001101000100101",
			1660 => "0000001001101000100101",
			1661 => "0000010000011000001000",
			1662 => "0010111010100100000100",
			1663 => "0000000001101000100101",
			1664 => "0000000001101000100101",
			1665 => "1111111001101000100101",
			1666 => "0000001101111000001100",
			1667 => "0001111011111000000100",
			1668 => "0000001001101000100101",
			1669 => "0001101010110000000100",
			1670 => "0000001001101000100101",
			1671 => "0000000001101000100101",
			1672 => "1111111001101000100101",
			1673 => "0011100011101000101000",
			1674 => "0001000011010000001100",
			1675 => "0001101101000100000100",
			1676 => "0000000001101010010001",
			1677 => "0000001100010100000100",
			1678 => "0000000001101010010001",
			1679 => "0000000001101010010001",
			1680 => "0010001001000100011000",
			1681 => "0001110001010000010000",
			1682 => "0000111001000100000100",
			1683 => "0000000001101010010001",
			1684 => "0001100100100000001000",
			1685 => "0001010101111000000100",
			1686 => "0000000001101010010001",
			1687 => "0000000001101010010001",
			1688 => "0000000001101010010001",
			1689 => "0001011000101000000100",
			1690 => "0000000001101010010001",
			1691 => "0000000001101010010001",
			1692 => "0000000001101010010001",
			1693 => "0000001101111000001100",
			1694 => "0000011101000000001000",
			1695 => "0001001100101000000100",
			1696 => "0000000001101010010001",
			1697 => "0000000001101010010001",
			1698 => "0000000001101010010001",
			1699 => "0000000001101010010001",
			1700 => "0010011001001000101000",
			1701 => "0011010110001100010000",
			1702 => "0000001110000100001000",
			1703 => "0001101101000100000100",
			1704 => "0000000001101100110101",
			1705 => "0000000001101100110101",
			1706 => "0010011100101000000100",
			1707 => "0000000001101100110101",
			1708 => "0000000001101100110101",
			1709 => "0001111101001000001100",
			1710 => "0000010111110000001000",
			1711 => "0001100111100000000100",
			1712 => "0000000001101100110101",
			1713 => "0000000001101100110101",
			1714 => "0000000001101100110101",
			1715 => "0010000101011100000100",
			1716 => "0000000001101100110101",
			1717 => "0000000000000000000100",
			1718 => "0000000001101100110101",
			1719 => "0000000001101100110101",
			1720 => "0000011000011000011000",
			1721 => "0001110001010000001100",
			1722 => "0000110011000000001000",
			1723 => "0001010110000000000100",
			1724 => "0000000001101100110101",
			1725 => "0000000001101100110101",
			1726 => "0000000001101100110101",
			1727 => "0011111101001100001000",
			1728 => "0000110001001000000100",
			1729 => "0000000001101100110101",
			1730 => "0000000001101100110101",
			1731 => "0000000001101100110101",
			1732 => "0001011101101000001000",
			1733 => "0000101000110100000100",
			1734 => "0000000001101100110101",
			1735 => "0000000001101100110101",
			1736 => "0000010011000000001000",
			1737 => "0001000011010000000100",
			1738 => "0000000001101100110101",
			1739 => "0000000001101100110101",
			1740 => "0000000001101100110101",
			1741 => "0010000101101100100000",
			1742 => "0001110110101100001100",
			1743 => "0000101010101100001000",
			1744 => "0011101111100100000100",
			1745 => "0000000001101111001001",
			1746 => "0000000001101111001001",
			1747 => "0000000001101111001001",
			1748 => "0000001101111000010000",
			1749 => "0010101011111000001000",
			1750 => "0001011000000000000100",
			1751 => "0000000001101111001001",
			1752 => "0000000001101111001001",
			1753 => "0011011110011000000100",
			1754 => "0000000001101111001001",
			1755 => "0000000001101111001001",
			1756 => "0000000001101111001001",
			1757 => "0011110100110100100000",
			1758 => "0000101011101000010100",
			1759 => "0001110001010000001100",
			1760 => "0001001110011000001000",
			1761 => "0001001011101100000100",
			1762 => "0000000001101111001001",
			1763 => "0000000001101111001001",
			1764 => "0000000001101111001001",
			1765 => "0010010011000000000100",
			1766 => "0000000001101111001001",
			1767 => "0000000001101111001001",
			1768 => "0000111100101100000100",
			1769 => "0000000001101111001001",
			1770 => "0001001100110000000100",
			1771 => "0000000001101111001001",
			1772 => "0000000001101111001001",
			1773 => "0001000101010100000100",
			1774 => "0000000001101111001001",
			1775 => "0000011101000000000100",
			1776 => "0000000001101111001001",
			1777 => "0000000001101111001001",
			1778 => "0010011101101000110000",
			1779 => "0001111101001000010000",
			1780 => "0011101111000000000100",
			1781 => "1111111001110000111101",
			1782 => "0000100000001100000100",
			1783 => "0000011001110000111101",
			1784 => "0001011101101000000100",
			1785 => "0000000001110000111101",
			1786 => "1111111001110000111101",
			1787 => "0000000011001100010100",
			1788 => "0001100100001000010000",
			1789 => "0000000011011100001100",
			1790 => "0011110011101000000100",
			1791 => "0000010001110000111101",
			1792 => "0011110100000100000100",
			1793 => "0000011001110000111101",
			1794 => "0000011001110000111101",
			1795 => "0000001001110000111101",
			1796 => "0000100001110000111101",
			1797 => "0011100101001100001000",
			1798 => "0000111111101000000100",
			1799 => "1111111001110000111101",
			1800 => "0000000001110000111101",
			1801 => "0000011001110000111101",
			1802 => "0010001001000100001000",
			1803 => "0001111011000000000100",
			1804 => "1111111001110000111101",
			1805 => "0000010001110000111101",
			1806 => "1111111001110000111101",
			1807 => "0011101100011000100000",
			1808 => "0001000101011100010000",
			1809 => "0001101101000100000100",
			1810 => "0000000001110011000001",
			1811 => "0000000001110100001000",
			1812 => "0000010111110000000100",
			1813 => "0000000001110011000001",
			1814 => "0000000001110011000001",
			1815 => "0000000001110011000001",
			1816 => "0000110011000000001100",
			1817 => "0000110101101100000100",
			1818 => "0000000001110011000001",
			1819 => "0001011111011000000100",
			1820 => "0000000001110011000001",
			1821 => "0000000001110011000001",
			1822 => "0000000001110011000001",
			1823 => "0000001101111000100000",
			1824 => "0000111100110000001100",
			1825 => "0011100011101000001000",
			1826 => "0000000011011100000100",
			1827 => "0000000001110011000001",
			1828 => "0000000001110011000001",
			1829 => "0000000001110011000001",
			1830 => "0011100100000100010000",
			1831 => "0000111000101000001000",
			1832 => "0011111100111100000100",
			1833 => "0000000001110011000001",
			1834 => "0000000001110011000001",
			1835 => "0001100100001000000100",
			1836 => "0000000001110011000001",
			1837 => "0000000001110011000001",
			1838 => "0000000001110011000001",
			1839 => "0000000001110011000001",
			1840 => "0011101100011000100100",
			1841 => "0010010101010100001100",
			1842 => "0001111000000100000100",
			1843 => "0000000001110101001101",
			1844 => "0000001100010100000100",
			1845 => "0000000001110101001101",
			1846 => "0000000001110101001101",
			1847 => "0001110001010000001100",
			1848 => "0010001010100100000100",
			1849 => "0000000001110101001101",
			1850 => "0000011000111100000100",
			1851 => "0000000001110101001101",
			1852 => "0000000001110101001101",
			1853 => "0010001001000100001000",
			1854 => "0001111011111000000100",
			1855 => "0000000001110101001101",
			1856 => "0000000001110101001101",
			1857 => "0000000001110101001101",
			1858 => "0000001101111000100000",
			1859 => "0000111100110000001100",
			1860 => "0000011001100000001000",
			1861 => "0000101000011100000100",
			1862 => "0000000001110101001101",
			1863 => "0000000001110101001101",
			1864 => "0000000001110101001101",
			1865 => "0010000101101100000100",
			1866 => "0000000001110101001101",
			1867 => "0000111000101000001000",
			1868 => "0001100000001100000100",
			1869 => "0000000001110101001101",
			1870 => "0000000001110101001101",
			1871 => "0000001100001000000100",
			1872 => "0000000001110101001101",
			1873 => "0000000001110101001101",
			1874 => "0000000001110101001101",
			1875 => "0011101100011000100100",
			1876 => "0001000101011100010000",
			1877 => "0001101101000100000100",
			1878 => "1111111001110111010001",
			1879 => "0000000101011000001000",
			1880 => "0010111110011000000100",
			1881 => "0000001001110111010001",
			1882 => "0000000001110111010001",
			1883 => "1111111001110111010001",
			1884 => "0001110001010000001100",
			1885 => "0000110011000000001000",
			1886 => "0010100011000000000100",
			1887 => "0000000001110111010001",
			1888 => "0000000001110111010001",
			1889 => "1111111001110111010001",
			1890 => "0001011100010000000100",
			1891 => "0000000001110111010001",
			1892 => "1111111001110111010001",
			1893 => "0000001101111000011100",
			1894 => "0000110011100100000100",
			1895 => "0000001001110111010001",
			1896 => "0010000101101100001000",
			1897 => "0010111110011000000100",
			1898 => "0000001001110111010001",
			1899 => "0000000001110111010001",
			1900 => "0011011010100100000100",
			1901 => "0000000001110111010001",
			1902 => "0000000011001100001000",
			1903 => "0010101011000000000100",
			1904 => "0000001001110111010001",
			1905 => "1111111001110111010001",
			1906 => "1111111001110111010001",
			1907 => "1111111001110111010001",
			1908 => "0010000101101100011100",
			1909 => "0001101101000100000100",
			1910 => "0000000001111001001101",
			1911 => "0000001101111000010100",
			1912 => "0001010011110100010000",
			1913 => "0011011101000000000100",
			1914 => "0000000001111001001101",
			1915 => "0000010111100100000100",
			1916 => "0000000001111001001101",
			1917 => "0000011001100000000100",
			1918 => "0000000001111001001101",
			1919 => "0000000001111001001101",
			1920 => "0000000001111001001101",
			1921 => "0000000001111001001101",
			1922 => "0000110011100100001000",
			1923 => "0011101111010100000100",
			1924 => "0000000001111001001101",
			1925 => "0000000001111001001101",
			1926 => "0000000011011100001000",
			1927 => "0001011100110000000100",
			1928 => "0000000001111001001101",
			1929 => "0000000001111001001101",
			1930 => "0001001111011000001100",
			1931 => "0001110011000100001000",
			1932 => "0011010101010100000100",
			1933 => "0000000001111001001101",
			1934 => "0000000001111001001101",
			1935 => "0000000001111001001101",
			1936 => "0011000101011100000100",
			1937 => "0000000001111001001101",
			1938 => "0000000001111001001101",
			1939 => "0001000101011100101000",
			1940 => "0001111011111000011100",
			1941 => "0001111100010000001100",
			1942 => "0000100001000000001000",
			1943 => "0000001110100000000100",
			1944 => "0000000001111011110001",
			1945 => "0000000001111011110001",
			1946 => "0000000001111011110001",
			1947 => "0000000110010100001000",
			1948 => "0010011101101000000100",
			1949 => "0000000001111011110001",
			1950 => "0000000001111011110001",
			1951 => "0000001010010100000100",
			1952 => "0000000001111011110001",
			1953 => "0000000001111011110001",
			1954 => "0001111011000000001000",
			1955 => "0010001111001000000100",
			1956 => "0000000001111011110001",
			1957 => "0000000001111011110001",
			1958 => "0000000001111011110001",
			1959 => "0001001111011000100000",
			1960 => "0000000111000100010100",
			1961 => "0011100100001100010000",
			1962 => "0010110101010100001100",
			1963 => "0000110011000000001000",
			1964 => "0000110110000000000100",
			1965 => "0000000001111011110001",
			1966 => "0000000001111011110001",
			1967 => "0000000001111011110001",
			1968 => "0000000001111011110001",
			1969 => "0000000001111011110001",
			1970 => "0001111000100000000100",
			1971 => "0000000001111011110001",
			1972 => "0001110000111100000100",
			1973 => "0000000001111011110001",
			1974 => "0000000001111011110001",
			1975 => "0011100110111000000100",
			1976 => "0000000001111011110001",
			1977 => "0000000100010100000100",
			1978 => "0000000001111011110001",
			1979 => "0000000001111011110001",
			1980 => "0010011101101000110000",
			1981 => "0001111001010000010100",
			1982 => "0001010011001000010000",
			1983 => "0011101111111000000100",
			1984 => "1111111001111101100101",
			1985 => "0000000101011000001000",
			1986 => "0011101110111100000100",
			1987 => "0000001001111101100101",
			1988 => "0000010001111101100101",
			1989 => "1111111001111101100101",
			1990 => "1111111001111101100101",
			1991 => "0000001101111000011000",
			1992 => "0011000101010100010100",
			1993 => "0000111100110000001100",
			1994 => "0011111001111000001000",
			1995 => "0010000101101100000100",
			1996 => "0000010001111101100101",
			1997 => "0000001001111101100101",
			1998 => "0000010001111101100101",
			1999 => "0011100100000100000100",
			2000 => "0000001001111101100101",
			2001 => "0000000001111101100101",
			2002 => "0000010001111101100101",
			2003 => "1111111001111101100101",
			2004 => "0010001001000100001000",
			2005 => "0001100100101000000100",
			2006 => "1111111001111101100101",
			2007 => "0000010001111101100101",
			2008 => "1111111001111101100101",
			2009 => "0010000101101100101000",
			2010 => "0011011110011000011100",
			2011 => "0001111001010000010000",
			2012 => "0000001110000100001000",
			2013 => "0001101101000100000100",
			2014 => "0000000010000000011001",
			2015 => "0000000010000000011001",
			2016 => "0010111010100100000100",
			2017 => "0000000010000000011001",
			2018 => "0000000010000000011001",
			2019 => "0000001101111000001000",
			2020 => "0011010110001100000100",
			2021 => "0000000010000000011001",
			2022 => "0000000010000000011001",
			2023 => "0000000010000000011001",
			2024 => "0000001110110100001000",
			2025 => "0011110100010000000100",
			2026 => "0000000010000000011001",
			2027 => "0000000010000000011001",
			2028 => "0000000010000000011001",
			2029 => "0011101100000100100000",
			2030 => "0010111011101100001000",
			2031 => "0001000101010100000100",
			2032 => "0000000010000000011001",
			2033 => "0000000010000000011001",
			2034 => "0000101011101000001100",
			2035 => "0000000101111100000100",
			2036 => "0000000010000000011001",
			2037 => "0001001111011000000100",
			2038 => "0000000010000000011001",
			2039 => "0000000010000000011001",
			2040 => "0000111100101100000100",
			2041 => "0000000010000000011001",
			2042 => "0001000110101100000100",
			2043 => "0000000010000000011001",
			2044 => "0000000010000000011001",
			2045 => "0011110000011100001100",
			2046 => "0011110100110100000100",
			2047 => "0000000010000000011001",
			2048 => "0010101011000000000100",
			2049 => "0000000010000000011001",
			2050 => "0000000010000000011001",
			2051 => "0000111101001000000100",
			2052 => "0000000010000000011001",
			2053 => "0000000010000000011001",
			2054 => "0001100010001000001100",
			2055 => "0010010111011100001000",
			2056 => "0011011101000000000100",
			2057 => "1111111010000010100101",
			2058 => "0000001010000010100101",
			2059 => "1111111010000010100101",
			2060 => "0000000010100100101000",
			2061 => "0010000101101100010100",
			2062 => "0001111100010000000100",
			2063 => "1111111010000010100101",
			2064 => "0010101011111000001100",
			2065 => "0011101100011000001000",
			2066 => "0000000101000100000100",
			2067 => "0000001010000010100101",
			2068 => "0000000010000010100101",
			2069 => "0000001010000010100101",
			2070 => "0000000010000010100101",
			2071 => "0011100010110000001000",
			2072 => "0000010111100100000100",
			2073 => "0000000010000010100101",
			2074 => "1111111010000010100101",
			2075 => "0000101011100000000100",
			2076 => "0000001010000010100101",
			2077 => "0000111000101000000100",
			2078 => "1111111010000010100101",
			2079 => "0000001010000010100101",
			2080 => "0011110011100000001100",
			2081 => "0001000101010100001000",
			2082 => "0010111011101100000100",
			2083 => "1111111010000010100101",
			2084 => "0000000010000010100101",
			2085 => "1111111010000010100101",
			2086 => "0000101010111000000100",
			2087 => "0000001010000010100101",
			2088 => "1111111010000010100101",
			2089 => "0001111001010000011000",
			2090 => "0000010111110000010100",
			2091 => "0001011111011000010000",
			2092 => "0010101010000100000100",
			2093 => "0000000010000100110001",
			2094 => "0000000000100100001000",
			2095 => "0000100100010000000100",
			2096 => "0000000010000100110001",
			2097 => "0000000010000100110001",
			2098 => "0000000010000100110001",
			2099 => "0000000010000100110001",
			2100 => "0000000010000100110001",
			2101 => "0010000101101100010000",
			2102 => "0000000110010100001000",
			2103 => "0010011010000100000100",
			2104 => "0000001010000100110001",
			2105 => "0000000010000100110001",
			2106 => "0000111100010000000100",
			2107 => "0000000010000100110001",
			2108 => "0000000010000100110001",
			2109 => "0011011110011000000100",
			2110 => "0000000010000100110001",
			2111 => "0000111100110000001100",
			2112 => "0010010110000000000100",
			2113 => "0000001010000100110001",
			2114 => "0000010011110000000100",
			2115 => "0000000010000100110001",
			2116 => "0000000010000100110001",
			2117 => "0000111000101000001000",
			2118 => "0011110000001000000100",
			2119 => "0000000010000100110001",
			2120 => "0000000010000100110001",
			2121 => "0010011010000100000100",
			2122 => "0000000010000100110001",
			2123 => "0000000010000100110001",
			2124 => "0011101100011000101100",
			2125 => "0001000101011100010100",
			2126 => "0011100000010100001100",
			2127 => "0010010101010100001000",
			2128 => "0000111110011000000100",
			2129 => "0000000010000111000101",
			2130 => "0000001010000111000101",
			2131 => "1111111010000111000101",
			2132 => "0000000101011000000100",
			2133 => "0000001010000111000101",
			2134 => "1111111010000111000101",
			2135 => "0001110001010000010000",
			2136 => "0000110011000000001100",
			2137 => "0001011111011000001000",
			2138 => "0010100101101100000100",
			2139 => "0000000010000111000101",
			2140 => "0000000010000111000101",
			2141 => "0000000010000111000101",
			2142 => "1111111010000111000101",
			2143 => "0001011100010000000100",
			2144 => "0000000010000111000101",
			2145 => "1111111010000111000101",
			2146 => "0000001101111000011100",
			2147 => "0000110011100100000100",
			2148 => "0000001010000111000101",
			2149 => "0010000101101100001000",
			2150 => "0010111110011000000100",
			2151 => "0000001010000111000101",
			2152 => "0000000010000111000101",
			2153 => "0011011010100100000100",
			2154 => "0000000010000111000101",
			2155 => "0000011101000000000100",
			2156 => "0000001010000111000101",
			2157 => "0000001011010000000100",
			2158 => "0000000010000111000101",
			2159 => "1111111010000111000101",
			2160 => "1111111010000111000101",
			2161 => "0010011010000100101000",
			2162 => "0011101111000000000100",
			2163 => "1111111010001000101001",
			2164 => "0000001101111000100000",
			2165 => "0001010011000000001000",
			2166 => "0000101011001000000100",
			2167 => "0000001010001000101001",
			2168 => "0000000010001000101001",
			2169 => "0001111001010000001000",
			2170 => "0000001101001100000100",
			2171 => "0000000010001000101001",
			2172 => "1111111010001000101001",
			2173 => "0010000101101100001000",
			2174 => "0000000110010100000100",
			2175 => "0000001010001000101001",
			2176 => "0000000010001000101001",
			2177 => "0011010011010000000100",
			2178 => "0000000010001000101001",
			2179 => "0000001010001000101001",
			2180 => "1111111010001000101001",
			2181 => "0000010111100100001000",
			2182 => "0001111011000000000100",
			2183 => "1111111010001000101001",
			2184 => "0000001010001000101001",
			2185 => "1111111010001000101001",
			2186 => "0011101100011000100000",
			2187 => "0000011000011000011100",
			2188 => "0001011100010000011000",
			2189 => "0001111100010000001100",
			2190 => "0001011100101000001000",
			2191 => "0010101111111100000100",
			2192 => "1111111010001010011101",
			2193 => "0000001010001010011101",
			2194 => "1111111010001010011101",
			2195 => "0000001110110100001000",
			2196 => "0001100010001000000100",
			2197 => "0000000010001010011101",
			2198 => "0000001010001010011101",
			2199 => "1111111010001010011101",
			2200 => "1111111010001010011101",
			2201 => "1111111010001010011101",
			2202 => "0000001101111000011000",
			2203 => "0000110011100100000100",
			2204 => "0000001010001010011101",
			2205 => "0010000101101100000100",
			2206 => "0000001010001010011101",
			2207 => "0011011010100100000100",
			2208 => "0000000010001010011101",
			2209 => "0000100010101100001000",
			2210 => "0010101011000000000100",
			2211 => "0000001010001010011101",
			2212 => "1111111010001010011101",
			2213 => "1111111010001010011101",
			2214 => "1111111010001010011101",
			2215 => "0001100000100100111100",
			2216 => "0000000011001100101100",
			2217 => "0001000011010000001100",
			2218 => "0001101101000100000100",
			2219 => "0000000010001100100001",
			2220 => "0000010110010000000100",
			2221 => "0000000010001100100001",
			2222 => "0000001010001100100001",
			2223 => "0011100111001000010100",
			2224 => "0001011101101000001000",
			2225 => "0001000101011100000100",
			2226 => "0000000010001100100001",
			2227 => "0000000010001100100001",
			2228 => "0001110001010000000100",
			2229 => "1111111010001100100001",
			2230 => "0010110101011100000100",
			2231 => "0000000010001100100001",
			2232 => "0000000010001100100001",
			2233 => "0011011010100100000100",
			2234 => "0000000010001100100001",
			2235 => "0010101011000000000100",
			2236 => "0000000010001100100001",
			2237 => "0000000010001100100001",
			2238 => "0011010110110100001000",
			2239 => "0001011001010000000100",
			2240 => "0000000010001100100001",
			2241 => "0000000010001100100001",
			2242 => "0001010101111000000100",
			2243 => "0000000010001100100001",
			2244 => "1111111010001100100001",
			2245 => "0000111001010100000100",
			2246 => "0000000010001100100001",
			2247 => "0000000010001100100001",
			2248 => "0011101010001001000000",
			2249 => "0000101011101000100100",
			2250 => "0011101110111100011000",
			2251 => "0010010101010100001100",
			2252 => "0011011101000000000100",
			2253 => "0000000010001111000101",
			2254 => "0000111110011000000100",
			2255 => "0000000010001111000101",
			2256 => "0000000010001111000101",
			2257 => "0011010110110100000100",
			2258 => "0000000010001111000101",
			2259 => "0010000011010000000100",
			2260 => "0000000010001111000101",
			2261 => "0000000010001111000101",
			2262 => "0001011001010100001000",
			2263 => "0001101111010100000100",
			2264 => "0000000010001111000101",
			2265 => "0000000010001111000101",
			2266 => "0000000010001111000101",
			2267 => "0001001001000100000100",
			2268 => "0000000010001111000101",
			2269 => "0001100100001000010000",
			2270 => "0010000101101100001100",
			2271 => "0011111101010100001000",
			2272 => "0001100100011100000100",
			2273 => "0000000010001111000101",
			2274 => "0000000010001111000101",
			2275 => "0000000010001111000101",
			2276 => "0000000010001111000101",
			2277 => "0001101110101100000100",
			2278 => "0000000010001111000101",
			2279 => "0000000010001111000101",
			2280 => "0010001111001000001100",
			2281 => "0000000110101000000100",
			2282 => "0000000010001111000101",
			2283 => "0011110011100000000100",
			2284 => "0000000010001111000101",
			2285 => "0000000010001111000101",
			2286 => "0011111011110100000100",
			2287 => "0000000010001111000101",
			2288 => "0000000010001111000101",
			2289 => "0010011101101000110000",
			2290 => "0001111100010000001100",
			2291 => "0010010101010100001000",
			2292 => "0001111000000100000100",
			2293 => "1111111010010000111001",
			2294 => "0000001010010000111001",
			2295 => "1111111010010000111001",
			2296 => "0000001101111000100000",
			2297 => "0010101011000000011100",
			2298 => "0001000101011100001100",
			2299 => "0010111011101100000100",
			2300 => "0000001010010000111001",
			2301 => "0011111000001000000100",
			2302 => "0000001010010000111001",
			2303 => "0000010010010000111001",
			2304 => "0001110001010000001000",
			2305 => "0010011001001000000100",
			2306 => "0000000010010000111001",
			2307 => "1111111010010000111001",
			2308 => "0011100010110100000100",
			2309 => "0000001010010000111001",
			2310 => "0000000010010000111001",
			2311 => "1111111010010000111001",
			2312 => "1111111010010000111001",
			2313 => "0010001001000100001000",
			2314 => "0001111011000000000100",
			2315 => "1111111010010000111001",
			2316 => "0000010010010000111001",
			2317 => "1111111010010000111001",
			2318 => "0010011101101000111100",
			2319 => "0001111101001000011000",
			2320 => "0001000101011100010000",
			2321 => "0001101101000100000100",
			2322 => "1111111010010011000101",
			2323 => "0000001110000100000100",
			2324 => "0000001010010011000101",
			2325 => "0010010101011100000100",
			2326 => "1111111010010011000101",
			2327 => "0000000010010011000101",
			2328 => "0000111001000100000100",
			2329 => "0000000010010011000101",
			2330 => "1111111010010011000101",
			2331 => "0000001101111000100000",
			2332 => "0000111100110000010100",
			2333 => "0010001001000100001100",
			2334 => "0011100100010000001000",
			2335 => "0011111010101100000100",
			2336 => "0000001010010011000101",
			2337 => "0000000010010011000101",
			2338 => "0000001010010011000101",
			2339 => "0001110001010000000100",
			2340 => "1111111010010011000101",
			2341 => "0000001010010011000101",
			2342 => "0011011011101100000100",
			2343 => "1111111010010011000101",
			2344 => "0000000110101000000100",
			2345 => "0000001010010011000101",
			2346 => "0000000010010011000101",
			2347 => "1111111010010011000101",
			2348 => "0010010011000000001000",
			2349 => "0001111100101100000100",
			2350 => "1111111010010011000101",
			2351 => "0000001010010011000101",
			2352 => "1111111010010011000101",
			2353 => "0011110011010100001100",
			2354 => "0010110110001100001000",
			2355 => "0010111101000000000100",
			2356 => "1111111010010101010001",
			2357 => "0000000010010101010001",
			2358 => "1111111010010101010001",
			2359 => "0000000011001100101000",
			2360 => "0001010011110100100100",
			2361 => "0001000111011100001100",
			2362 => "0011001110011000000100",
			2363 => "0000001010010101010001",
			2364 => "0000000101011000000100",
			2365 => "0000001010010101010001",
			2366 => "0000001010010101010001",
			2367 => "0001110001010000001100",
			2368 => "0011011110011000001000",
			2369 => "0000000111000100000100",
			2370 => "0000001010010101010001",
			2371 => "1111111010010101010001",
			2372 => "1111111010010101010001",
			2373 => "0000010111100100000100",
			2374 => "0000001010010101010001",
			2375 => "0011011010100100000100",
			2376 => "0000000010010101010001",
			2377 => "0000001010010101010001",
			2378 => "1111111010010101010001",
			2379 => "0001101011010100001100",
			2380 => "0011010110110100001000",
			2381 => "0001011001010000000100",
			2382 => "1111111010010101010001",
			2383 => "0000001010010101010001",
			2384 => "1111111010010101010001",
			2385 => "0000111100110000000100",
			2386 => "0000001010010101010001",
			2387 => "1111111010010101010001",
			2388 => "0011100011101000110100",
			2389 => "0000001011111100110000",
			2390 => "0010001001000100011100",
			2391 => "0011101101000100010000",
			2392 => "0010010101010100001000",
			2393 => "0010100101101100000100",
			2394 => "0000000010010111110101",
			2395 => "0000000010010111110101",
			2396 => "0011010110110100000100",
			2397 => "0000000010010111110101",
			2398 => "0000000010010111110101",
			2399 => "0000111111101000001000",
			2400 => "0001111101001000000100",
			2401 => "0000000010010111110101",
			2402 => "0000001010010111110101",
			2403 => "0000000010010111110101",
			2404 => "0001000011010000001000",
			2405 => "0000101100111000000100",
			2406 => "0000000010010111110101",
			2407 => "0000000010010111110101",
			2408 => "0001001010000100000100",
			2409 => "1111111010010111110101",
			2410 => "0001000101111000000100",
			2411 => "0000000010010111110101",
			2412 => "0000000010010111110101",
			2413 => "1111111010010111110101",
			2414 => "0000111000101000010100",
			2415 => "0000111001010100010000",
			2416 => "0001100000100100001100",
			2417 => "0000000110101000000100",
			2418 => "0000000010010111110101",
			2419 => "0010101001010100000100",
			2420 => "0000000010010111110101",
			2421 => "1111111010010111110101",
			2422 => "0000000010010111110101",
			2423 => "1111111010010111110101",
			2424 => "0011100100000100001000",
			2425 => "0000000000000000000100",
			2426 => "0000001010010111110101",
			2427 => "0000000010010111110101",
			2428 => "0000000010010111110101",
			2429 => "0011100010010100001100",
			2430 => "0010010101010100001000",
			2431 => "0000001110100100000100",
			2432 => "1111111010011001100001",
			2433 => "0000001010011001100001",
			2434 => "1111111010011001100001",
			2435 => "0000001101111000101000",
			2436 => "0010010101111000100100",
			2437 => "0000000011001100010100",
			2438 => "0011101010001000010000",
			2439 => "0010001001000100001000",
			2440 => "0000001011111100000100",
			2441 => "0000001010011001100001",
			2442 => "1111111010011001100001",
			2443 => "0000000001110100000100",
			2444 => "0000000010011001100001",
			2445 => "1111111010011001100001",
			2446 => "0000001010011001100001",
			2447 => "0000101101011100001100",
			2448 => "0001000111011100000100",
			2449 => "1111111010011001100001",
			2450 => "0001001001000100000100",
			2451 => "0000001010011001100001",
			2452 => "1111111010011001100001",
			2453 => "0000001010011001100001",
			2454 => "1111111010011001100001",
			2455 => "1111111010011001100001",
			2456 => "0011100110000101000000",
			2457 => "0001011010000100001100",
			2458 => "0001101101000100000100",
			2459 => "0000000010011011111101",
			2460 => "0000001100010100000100",
			2461 => "0000000010011011111101",
			2462 => "0000000010011011111101",
			2463 => "0010010101011100001100",
			2464 => "0000001110110100001000",
			2465 => "0001101010110100000100",
			2466 => "0000000010011011111101",
			2467 => "0000000010011011111101",
			2468 => "0000000010011011111101",
			2469 => "0001111100101100011000",
			2470 => "0010001001001100001100",
			2471 => "0010000011010000000100",
			2472 => "0000000010011011111101",
			2473 => "0011000111011100000100",
			2474 => "0000000010011011111101",
			2475 => "0000000010011011111101",
			2476 => "0011001110011000000100",
			2477 => "0000000010011011111101",
			2478 => "0011000101011100000100",
			2479 => "0000000010011011111101",
			2480 => "0000000010011011111101",
			2481 => "0000011000011000001000",
			2482 => "0001100001000000000100",
			2483 => "0000000010011011111101",
			2484 => "0000000010011011111101",
			2485 => "0010001010000100000100",
			2486 => "0000000010011011111101",
			2487 => "0000000010011011111101",
			2488 => "0010111011101100000100",
			2489 => "0000000010011011111101",
			2490 => "0000011101000000001000",
			2491 => "0000011001100000000100",
			2492 => "0000000010011011111101",
			2493 => "0000000010011011111101",
			2494 => "0000000010011011111101",
			2495 => "0010011010000101001100",
			2496 => "0001111001010000101100",
			2497 => "0001011010000100010100",
			2498 => "0001101111000100001100",
			2499 => "0010110110001100001000",
			2500 => "0001010011010000000100",
			2501 => "0000000010011110101001",
			2502 => "0000001010011110101001",
			2503 => "1111111010011110101001",
			2504 => "0000001100010100000100",
			2505 => "0000001010011110101001",
			2506 => "1111111010011110101001",
			2507 => "0001000011010000001000",
			2508 => "0011110000000100000100",
			2509 => "0000000010011110101001",
			2510 => "1111111010011110101001",
			2511 => "0001111101001000001000",
			2512 => "0010001010100100000100",
			2513 => "0000000010011110101001",
			2514 => "1111111010011110101001",
			2515 => "0001011000111000000100",
			2516 => "0000000010011110101001",
			2517 => "1111111010011110101001",
			2518 => "0000001101111000011100",
			2519 => "0000010111100100001000",
			2520 => "0001111011111000000100",
			2521 => "0000000010011110101001",
			2522 => "0000001010011110101001",
			2523 => "0011011010100100001100",
			2524 => "0010001001000100001000",
			2525 => "0000001010000000000100",
			2526 => "0000001010011110101001",
			2527 => "0000000010011110101001",
			2528 => "0000000010011110101001",
			2529 => "0011101111010100000100",
			2530 => "1111111010011110101001",
			2531 => "0000001010011110101001",
			2532 => "1111111010011110101001",
			2533 => "0000010000011000001000",
			2534 => "0001000110000000000100",
			2535 => "0000000010011110101001",
			2536 => "1111111010011110101001",
			2537 => "1111111010011110101001",
			2538 => "0001101101010100111100",
			2539 => "0011111011000100110000",
			2540 => "0001100100001000101100",
			2541 => "0000000011011100100000",
			2542 => "0011101001011100010000",
			2543 => "0010010101010100001000",
			2544 => "0010100101101100000100",
			2545 => "0000000010100000101111",
			2546 => "0000000010100000101111",
			2547 => "0000011000111100000100",
			2548 => "0000000010100000101111",
			2549 => "0000000010100000101111",
			2550 => "0001011100110000001000",
			2551 => "0000000101111100000100",
			2552 => "0000000010100000101111",
			2553 => "0000000010100000101111",
			2554 => "0010001010000100000100",
			2555 => "0000000010100000101111",
			2556 => "0000000010100000101111",
			2557 => "0001111011000000000100",
			2558 => "0000000010100000101111",
			2559 => "0010001111001000000100",
			2560 => "0000000010100000101111",
			2561 => "0000000010100000101111",
			2562 => "0000000010100000101111",
			2563 => "0001110011000100000100",
			2564 => "0000000010100000101111",
			2565 => "0011100100110000000100",
			2566 => "0000000010100000101111",
			2567 => "0000000010100000101111",
			2568 => "0000001101111000000100",
			2569 => "0000000010100000101111",
			2570 => "0000000010100000101111",
			2571 => "0000111100110000100000",
			2572 => "0011100011101000011000",
			2573 => "0000001011101000010000",
			2574 => "0011100000010100001100",
			2575 => "0001011100101000001000",
			2576 => "0001111000000100000100",
			2577 => "0000000010100010010001",
			2578 => "0000000010100010010001",
			2579 => "0000000010100010010001",
			2580 => "0000000010100010010001",
			2581 => "0000111100010000000100",
			2582 => "0000000010100010010001",
			2583 => "0000000010100010010001",
			2584 => "0000001011001100000100",
			2585 => "0000000010100010010001",
			2586 => "0000000010100010010001",
			2587 => "0000100011011100001000",
			2588 => "0011100011010100000100",
			2589 => "0000000010100010010001",
			2590 => "0000000010100010010001",
			2591 => "0001001111011000000100",
			2592 => "0000000010100010010001",
			2593 => "0010011010000100000100",
			2594 => "0000000010100010010001",
			2595 => "0000000010100010010001",
			2596 => "0010000101101100010100",
			2597 => "0000001101111000010000",
			2598 => "0011111111110000000100",
			2599 => "0000000010100011110101",
			2600 => "0001001111101000001000",
			2601 => "0011011101000000000100",
			2602 => "0000000010100011110101",
			2603 => "0000000010100011110101",
			2604 => "0000000010100011110101",
			2605 => "0000000010100011110101",
			2606 => "0011011010100100010000",
			2607 => "0000110011100100001000",
			2608 => "0010101100010000000100",
			2609 => "0000000010100011110101",
			2610 => "0000000010100011110101",
			2611 => "0010110111011100000100",
			2612 => "0000000010100011110101",
			2613 => "0000000010100011110101",
			2614 => "0000000011001100001100",
			2615 => "0011101111010100000100",
			2616 => "0000000010100011110101",
			2617 => "0000010110001100000100",
			2618 => "0000000010100011110101",
			2619 => "0000000010100011110101",
			2620 => "0000000010100011110101",
			2621 => "0011101100011000100100",
			2622 => "0001011101101000001100",
			2623 => "0011111111110000000100",
			2624 => "0000000010100101101001",
			2625 => "0000001110000100000100",
			2626 => "0000000010100101101001",
			2627 => "0000000010100101101001",
			2628 => "0001000011010000001000",
			2629 => "0001111100110000000100",
			2630 => "0000000010100101101001",
			2631 => "0000000010100101101001",
			2632 => "0001110001010000001000",
			2633 => "0000111001000100000100",
			2634 => "0000000010100101101001",
			2635 => "0000000010100101101001",
			2636 => "0010110101011100000100",
			2637 => "0000000010100101101001",
			2638 => "0000000010100101101001",
			2639 => "0000100010101100001000",
			2640 => "0011010101011100000100",
			2641 => "0000000010100101101001",
			2642 => "0000000010100101101001",
			2643 => "0001100000100100001000",
			2644 => "0010001001001100000100",
			2645 => "0000000010100101101001",
			2646 => "0000000010100101101001",
			2647 => "0000111001010100000100",
			2648 => "0000000010100101101001",
			2649 => "0000000010100101101001",
			2650 => "0000001110110100100000",
			2651 => "0011100101110100011000",
			2652 => "0001000101011100001100",
			2653 => "0001101101000100000100",
			2654 => "0000000010100111011101",
			2655 => "0000001011011100000100",
			2656 => "0000000010100111011101",
			2657 => "0000000010100111011101",
			2658 => "0000110011000000001000",
			2659 => "0000111101101000000100",
			2660 => "0000000010100111011101",
			2661 => "0000000010100111011101",
			2662 => "0000000010100111011101",
			2663 => "0000010110010000000100",
			2664 => "0000000010100111011101",
			2665 => "0000000010100111011101",
			2666 => "0011100101001100010100",
			2667 => "0000111000101000001100",
			2668 => "0001001000000100001000",
			2669 => "0001111000100000000100",
			2670 => "0000000010100111011101",
			2671 => "0000000010100111011101",
			2672 => "0000000010100111011101",
			2673 => "0010011010000100000100",
			2674 => "0000000010100111011101",
			2675 => "0000000010100111011101",
			2676 => "0000111001010100000100",
			2677 => "0000000010100111011101",
			2678 => "0000000010100111011101",
			2679 => "0011100010110100101000",
			2680 => "0000001011001000010000",
			2681 => "0011111111110000000100",
			2682 => "0000000010101001001001",
			2683 => "0001011100110000001000",
			2684 => "0000011000011000000100",
			2685 => "0000000010101001001001",
			2686 => "0000000010101001001001",
			2687 => "0000000010101001001001",
			2688 => "0001001000000100001100",
			2689 => "0001110110011100000100",
			2690 => "0000000010101001001001",
			2691 => "0001110001001000000100",
			2692 => "0000000010101001001001",
			2693 => "0000000010101001001001",
			2694 => "0011000101011100001000",
			2695 => "0001001100010000000100",
			2696 => "0000000010101001001001",
			2697 => "0000000010101001001001",
			2698 => "0000000010101001001001",
			2699 => "0000001101111000001100",
			2700 => "0010001111001000001000",
			2701 => "0000111100110000000100",
			2702 => "0000000010101001001001",
			2703 => "0000000010101001001001",
			2704 => "0000000010101001001001",
			2705 => "0000000010101001001001",
			2706 => "0010000101101100011100",
			2707 => "0001101101000100000100",
			2708 => "0000000010101010111101",
			2709 => "0011011110011000001100",
			2710 => "0000001101111000001000",
			2711 => "0011011101000000000100",
			2712 => "0000000010101010111101",
			2713 => "0000000010101010111101",
			2714 => "0000000010101010111101",
			2715 => "0000001110110100001000",
			2716 => "0011110100010000000100",
			2717 => "0000000010101010111101",
			2718 => "0000000010101010111101",
			2719 => "0000000010101010111101",
			2720 => "0011011010100100010000",
			2721 => "0000110011100100001000",
			2722 => "0001101010111100000100",
			2723 => "0000000010101010111101",
			2724 => "0000000010101010111101",
			2725 => "0000000011011100000100",
			2726 => "0000000010101010111101",
			2727 => "0000000010101010111101",
			2728 => "0010011101101000001100",
			2729 => "0000001111101100001000",
			2730 => "0011101111010100000100",
			2731 => "0000000010101010111101",
			2732 => "0000000010101010111101",
			2733 => "0000000010101010111101",
			2734 => "0000000010101010111101",
			2735 => "0010000101101100011000",
			2736 => "0001111001010000001100",
			2737 => "0000001110000100001000",
			2738 => "0001101101000100000100",
			2739 => "0000000010101100101001",
			2740 => "0000000010101100101001",
			2741 => "0000000010101100101001",
			2742 => "0000001101111000001000",
			2743 => "0010101011111000000100",
			2744 => "0000000010101100101001",
			2745 => "0000000010101100101001",
			2746 => "0000000010101100101001",
			2747 => "0000000011001100011000",
			2748 => "0001100100001000010100",
			2749 => "0000101011101000010000",
			2750 => "0011100101110100001100",
			2751 => "0010110101010100000100",
			2752 => "0000000010101100101001",
			2753 => "0010110101011100000100",
			2754 => "0000000010101100101001",
			2755 => "0000000010101100101001",
			2756 => "0000000010101100101001",
			2757 => "0000000010101100101001",
			2758 => "0000000010101100101001",
			2759 => "0000110011001000000100",
			2760 => "0000000010101100101001",
			2761 => "0000000010101100101001",
			2762 => "0011101001011100010100",
			2763 => "0010111011101100001000",
			2764 => "0001110011000000000100",
			2765 => "1111111010101110001101",
			2766 => "0000001010101110001101",
			2767 => "0011101001110000000100",
			2768 => "1111111010101110001101",
			2769 => "0000011000011000000100",
			2770 => "0000000010101110001101",
			2771 => "1111111010101110001101",
			2772 => "0000001101111000011100",
			2773 => "0010010101111000011000",
			2774 => "0000100011011100001100",
			2775 => "0011100001101100001000",
			2776 => "0001000101011100000100",
			2777 => "0000001010101110001101",
			2778 => "0000000010101110001101",
			2779 => "0000001010101110001101",
			2780 => "0011100110111000000100",
			2781 => "1111111010101110001101",
			2782 => "0000111100110000000100",
			2783 => "0000001010101110001101",
			2784 => "0000000010101110001101",
			2785 => "1111111010101110001101",
			2786 => "1111111010101110001101",
			2787 => "0010011101101000101100",
			2788 => "0001111001010000010100",
			2789 => "0000001110000100010000",
			2790 => "0000010111110000001000",
			2791 => "0001101101000100000100",
			2792 => "1111111010110000000001",
			2793 => "0000001010110000000001",
			2794 => "0010000101011100000100",
			2795 => "0000000010110000000001",
			2796 => "1111111010110000000001",
			2797 => "1111111010110000000001",
			2798 => "0000000011001100010000",
			2799 => "0001000101010100000100",
			2800 => "0000001010110000000001",
			2801 => "0011011010100100001000",
			2802 => "0001001001000100000100",
			2803 => "0000000010110000000001",
			2804 => "0000001010110000000001",
			2805 => "0000001010110000000001",
			2806 => "0001101011010100000100",
			2807 => "1111111010110000000001",
			2808 => "0000000010110000000001",
			2809 => "0000010000011000001100",
			2810 => "0001001100000000001000",
			2811 => "0001000001100100000100",
			2812 => "0000000010110000000001",
			2813 => "0000001010110000000001",
			2814 => "1111111010110000000001",
			2815 => "1111111010110000000001",
			2816 => "0001110001010000011100",
			2817 => "0010011001001000011000",
			2818 => "0000001110110100010100",
			2819 => "0001111100010000001100",
			2820 => "0001011100101000001000",
			2821 => "0000101101000100000100",
			2822 => "0000000010110001110101",
			2823 => "0000001010110001110101",
			2824 => "1111111010110001110101",
			2825 => "0001111101001000000100",
			2826 => "0000000010110001110101",
			2827 => "0000001010110001110101",
			2828 => "1111111010110001110101",
			2829 => "1111111010110001110101",
			2830 => "0000100011011100001000",
			2831 => "0010010101111000000100",
			2832 => "0000001010110001110101",
			2833 => "1111111010110001110101",
			2834 => "0010001111001000010000",
			2835 => "0000011001100000001000",
			2836 => "0000010111100100000100",
			2837 => "0000000010110001110101",
			2838 => "1111111010110001110101",
			2839 => "0011101100000100000100",
			2840 => "0000000010110001110101",
			2841 => "0000001010110001110101",
			2842 => "0000000011111000000100",
			2843 => "0000000010110001110101",
			2844 => "1111111010110001110101",
			2845 => "0000111100110000101100",
			2846 => "0011100011101000100000",
			2847 => "0000001011101000010100",
			2848 => "0011100010010100001100",
			2849 => "0010010101010100001000",
			2850 => "0010101111111100000100",
			2851 => "0000000010110100001001",
			2852 => "0000000010110100001001",
			2853 => "0000000010110100001001",
			2854 => "0010010101101100000100",
			2855 => "0000000010110100001001",
			2856 => "0000000010110100001001",
			2857 => "0010101000101000000100",
			2858 => "0000000010110100001001",
			2859 => "0010101111101000000100",
			2860 => "0000000010110100001001",
			2861 => "0000000010110100001001",
			2862 => "0010001111001000001000",
			2863 => "0000001011001100000100",
			2864 => "0000000010110100001001",
			2865 => "0000000010110100001001",
			2866 => "0000000010110100001001",
			2867 => "0010010101101100010000",
			2868 => "0000001010010100001000",
			2869 => "0000000111101100000100",
			2870 => "0000000010110100001001",
			2871 => "0000000010110100001001",
			2872 => "0000000101101000000100",
			2873 => "0000000010110100001001",
			2874 => "0000000010110100001001",
			2875 => "0011100011101000001000",
			2876 => "0001011001010000000100",
			2877 => "0000000010110100001001",
			2878 => "0000000010110100001001",
			2879 => "0000000110111100000100",
			2880 => "0000000010110100001001",
			2881 => "0000000010110100001001",
			2882 => "0001100100001000101000",
			2883 => "0000101011101000011100",
			2884 => "0011100101110100011000",
			2885 => "0010010101010100001000",
			2886 => "0011100101110000000100",
			2887 => "0000000010110101110101",
			2888 => "0000001010110101110101",
			2889 => "0011100010010100000100",
			2890 => "1111111010110101110101",
			2891 => "0000111111011000000100",
			2892 => "0000000010110101110101",
			2893 => "0000010111100100000100",
			2894 => "0000000010110101110101",
			2895 => "1111111010110101110101",
			2896 => "0000001010110101110101",
			2897 => "0010001001001100001000",
			2898 => "0001000101111000000100",
			2899 => "0000000010110101110101",
			2900 => "0000000010110101110101",
			2901 => "1111111010110101110101",
			2902 => "0000001101111000001100",
			2903 => "0001111011111000000100",
			2904 => "0000001010110101110101",
			2905 => "0001101010110000000100",
			2906 => "0000001010110101110101",
			2907 => "0000000010110101110101",
			2908 => "1111111010110101110101",
			2909 => "0001011100000000101100",
			2910 => "0000101001110100011100",
			2911 => "0001111100010000001100",
			2912 => "0001011100101000001000",
			2913 => "0001111000000100000100",
			2914 => "0000000010111000010001",
			2915 => "0000000010111000010001",
			2916 => "0000000010111000010001",
			2917 => "0001111011111000001000",
			2918 => "0001100010001000000100",
			2919 => "0000000010111000010001",
			2920 => "0000000010111000010001",
			2921 => "0001111100101100000100",
			2922 => "0000000010111000010001",
			2923 => "0000000010111000010001",
			2924 => "0000001010010100001000",
			2925 => "0000110011100100000100",
			2926 => "0000000010111000010001",
			2927 => "0000000010111000010001",
			2928 => "0000001110110000000100",
			2929 => "0000000010111000010001",
			2930 => "0000000010111000010001",
			2931 => "0001011001010000011000",
			2932 => "0011110000001000010000",
			2933 => "0001100100101000001000",
			2934 => "0010110111011100000100",
			2935 => "0000000010111000010001",
			2936 => "0000000010111000010001",
			2937 => "0000011000011000000100",
			2938 => "0000000010111000010001",
			2939 => "0000000010111000010001",
			2940 => "0010011001000100000100",
			2941 => "0000000010111000010001",
			2942 => "0000000010111000010001",
			2943 => "0001100000010000000100",
			2944 => "0000000010111000010001",
			2945 => "0011000101011100000100",
			2946 => "0000000010111000010001",
			2947 => "0000000010111000010001",
			2948 => "0001100010001000001100",
			2949 => "0010010101010100001000",
			2950 => "0001101110010100000100",
			2951 => "1111111010111001111101",
			2952 => "0000001010111001111101",
			2953 => "1111111010111001111101",
			2954 => "0000100011011100010100",
			2955 => "0001011001010000010000",
			2956 => "0010001001000100001100",
			2957 => "0010001111111100001000",
			2958 => "0000000101000100000100",
			2959 => "0000001010111001111101",
			2960 => "0000001010111001111101",
			2961 => "0000001010111001111101",
			2962 => "0000000010111001111101",
			2963 => "1111111010111001111101",
			2964 => "0011100110111000000100",
			2965 => "1111111010111001111101",
			2966 => "0000001101111000010000",
			2967 => "0001011001010000001000",
			2968 => "0011101100000100000100",
			2969 => "1111111010111001111101",
			2970 => "0000001010111001111101",
			2971 => "0011001010000100000100",
			2972 => "0000010010111001111101",
			2973 => "1111111010111001111101",
			2974 => "1111111010111001111101",
			2975 => "0010011101101000110000",
			2976 => "0001111100010000001100",
			2977 => "0010010101010100001000",
			2978 => "0001111000000100000100",
			2979 => "1111111010111100000001",
			2980 => "0000001010111100000001",
			2981 => "1111111010111100000001",
			2982 => "0000000011001100011000",
			2983 => "0001011100010000010000",
			2984 => "0000100011011100001100",
			2985 => "0001011000000100001000",
			2986 => "0010101000000100000100",
			2987 => "0000010010111100000001",
			2988 => "0000010010111100000001",
			2989 => "0000010010111100000001",
			2990 => "0000001010111100000001",
			2991 => "0001111111101000000100",
			2992 => "1111111010111100000001",
			2993 => "0000010010111100000001",
			2994 => "0011100101100000001000",
			2995 => "0001110100101100000100",
			2996 => "1111111010111100000001",
			2997 => "0000000010111100000001",
			2998 => "0000010010111100000001",
			2999 => "0000010000011000001000",
			3000 => "0001111001010100000100",
			3001 => "1111111010111100000001",
			3002 => "0000001010111100000001",
			3003 => "0010010011000000001000",
			3004 => "0001111100101100000100",
			3005 => "1111111010111100000001",
			3006 => "0000001010111100000001",
			3007 => "1111111010111100000001",
			3008 => "0010000101101100100000",
			3009 => "0001110110101100001100",
			3010 => "0000000001111000001000",
			3011 => "0011100101110000000100",
			3012 => "0000000010111110010101",
			3013 => "0000000010111110010101",
			3014 => "0000000010111110010101",
			3015 => "0000001101111000010000",
			3016 => "0010101011111000001000",
			3017 => "0001011000000000000100",
			3018 => "0000000010111110010101",
			3019 => "0000000010111110010101",
			3020 => "0010101100001100000100",
			3021 => "0000000010111110010101",
			3022 => "0000000010111110010101",
			3023 => "0000000010111110010101",
			3024 => "0011101100000100100000",
			3025 => "0010111011101100001000",
			3026 => "0001010011001000000100",
			3027 => "0000000010111110010101",
			3028 => "0000000010111110010101",
			3029 => "0000101011101000001100",
			3030 => "0001110001010000000100",
			3031 => "0000000010111110010101",
			3032 => "0001011100110000000100",
			3033 => "0000000010111110010101",
			3034 => "0000000010111110010101",
			3035 => "0000111100101100000100",
			3036 => "0000000010111110010101",
			3037 => "0001010000111100000100",
			3038 => "0000000010111110010101",
			3039 => "0000000010111110010101",
			3040 => "0010101111101000000100",
			3041 => "0000000010111110010101",
			3042 => "0011010101010100000100",
			3043 => "0000000010111110010101",
			3044 => "0000000010111110010101",
			3045 => "0001101101010100110000",
			3046 => "0000100011011100100000",
			3047 => "0011100101110100011000",
			3048 => "0000010111110000010100",
			3049 => "0000001110000100001100",
			3050 => "0000001110100000000100",
			3051 => "0000000011000000001001",
			3052 => "0010111010100100000100",
			3053 => "0000000011000000001001",
			3054 => "0000000011000000001001",
			3055 => "0000011001100100000100",
			3056 => "0000000011000000001001",
			3057 => "0000000011000000001001",
			3058 => "0000000011000000001001",
			3059 => "0001111011111000000100",
			3060 => "0000000011000000001001",
			3061 => "0000000011000000001001",
			3062 => "0011000111011100000100",
			3063 => "0000000011000000001001",
			3064 => "0011100110111000000100",
			3065 => "0000000011000000001001",
			3066 => "0010110101011100000100",
			3067 => "0000000011000000001001",
			3068 => "0000000011000000001001",
			3069 => "0010111011101100000100",
			3070 => "0000000011000000001001",
			3071 => "0000011101000000000100",
			3072 => "0000000011000000001001",
			3073 => "0000000011000000001001",
			3074 => "0010000101101100101000",
			3075 => "0011011110011000011100",
			3076 => "0001111001010000010000",
			3077 => "0000001110000100001000",
			3078 => "0001101101000100000100",
			3079 => "0000000011000010101101",
			3080 => "0000000011000010101101",
			3081 => "0010111010100100000100",
			3082 => "0000000011000010101101",
			3083 => "0000000011000010101101",
			3084 => "0000001101111000001000",
			3085 => "0011010110001100000100",
			3086 => "0000000011000010101101",
			3087 => "0000000011000010101101",
			3088 => "0000000011000010101101",
			3089 => "0000001110110100001000",
			3090 => "0011110100010000000100",
			3091 => "0000000011000010101101",
			3092 => "0000000011000010101101",
			3093 => "0000000011000010101101",
			3094 => "0010101000101000010100",
			3095 => "0011100010110100010000",
			3096 => "0000001011001000001100",
			3097 => "0000000101111100000100",
			3098 => "0000000011000010101101",
			3099 => "0001111000101000000100",
			3100 => "0000000011000010101101",
			3101 => "0000000011000010101101",
			3102 => "0000000011000010101101",
			3103 => "0000000011000010101101",
			3104 => "0011010101010100010000",
			3105 => "0000111100101100001000",
			3106 => "0000001101110100000100",
			3107 => "0000000011000010101101",
			3108 => "0000000011000010101101",
			3109 => "0001011110010100000100",
			3110 => "0000000011000010101101",
			3111 => "0000000011000010101101",
			3112 => "0010001111001000000100",
			3113 => "0000000011000010101101",
			3114 => "0000000011000010101101",
			3115 => "0001011100000000101000",
			3116 => "0000101001110100011100",
			3117 => "0011100111001000010100",
			3118 => "0000011000011000010000",
			3119 => "0001101101000100000100",
			3120 => "0000000011000100110001",
			3121 => "0000001110000100000100",
			3122 => "0000000011000100110001",
			3123 => "0000000011111100000100",
			3124 => "0000000011000100110001",
			3125 => "0000000011000100110001",
			3126 => "0000000011000100110001",
			3127 => "0011001010100100000100",
			3128 => "0000001011000100110001",
			3129 => "0000000011000100110001",
			3130 => "0010111011101100000100",
			3131 => "0000000011000100110001",
			3132 => "0010011001001000000100",
			3133 => "0000000011000100110001",
			3134 => "0000000011000100110001",
			3135 => "0001111011111000000100",
			3136 => "0000000011000100110001",
			3137 => "0010001001000100001000",
			3138 => "0000111001000000000100",
			3139 => "0000000011000100110001",
			3140 => "0000000011000100110001",
			3141 => "0000000011111000001100",
			3142 => "0000010110110100001000",
			3143 => "0000110001101000000100",
			3144 => "0000000011000100110001",
			3145 => "0000000011000100110001",
			3146 => "0000000011000100110001",
			3147 => "0000000011000100110001",
			3148 => "0001101101010100111000",
			3149 => "0000001110110100100000",
			3150 => "0011100010001000010100",
			3151 => "0000010111110000010000",
			3152 => "0011111111110000000100",
			3153 => "0000000011000110110101",
			3154 => "0000001110000100000100",
			3155 => "0000001011000110110101",
			3156 => "0001110110101100000100",
			3157 => "0000000011000110110101",
			3158 => "0000000011000110110101",
			3159 => "1111111011000110110101",
			3160 => "0010111110011000000100",
			3161 => "0000000011000110110101",
			3162 => "0011100100001100000100",
			3163 => "0000000011000110110101",
			3164 => "0000001011000110110101",
			3165 => "0000110011000100010000",
			3166 => "0011101100000100001100",
			3167 => "0000010000011000001000",
			3168 => "0001000101111000000100",
			3169 => "0000000011000110110101",
			3170 => "0000000011000110110101",
			3171 => "1111111011000110110101",
			3172 => "0000000011000110110101",
			3173 => "0000110001001000000100",
			3174 => "0000000011000110110101",
			3175 => "0000000011000110110101",
			3176 => "0010111011101100000100",
			3177 => "0000000011000110110101",
			3178 => "0000011101000000000100",
			3179 => "0000001011000110110101",
			3180 => "0000000011000110110101",
			3181 => "0001000101011100101000",
			3182 => "0001111011111000011100",
			3183 => "0001111100010000001100",
			3184 => "0000100001000000001000",
			3185 => "0000001110100000000100",
			3186 => "0000000011001001011001",
			3187 => "0000000011001001011001",
			3188 => "0000000011001001011001",
			3189 => "0000000110010100001000",
			3190 => "0010011101101000000100",
			3191 => "0000000011001001011001",
			3192 => "0000000011001001011001",
			3193 => "0000001010010100000100",
			3194 => "0000000011001001011001",
			3195 => "0000000011001001011001",
			3196 => "0001111011000000001000",
			3197 => "0010001111001000000100",
			3198 => "0000000011001001011001",
			3199 => "0000000011001001011001",
			3200 => "0000000011001001011001",
			3201 => "0001001111011000100000",
			3202 => "0000000111000100010100",
			3203 => "0011100100001100010000",
			3204 => "0010110101010100001100",
			3205 => "0000110011000000001000",
			3206 => "0000110110000000000100",
			3207 => "0000000011001001011001",
			3208 => "0000000011001001011001",
			3209 => "0000000011001001011001",
			3210 => "0000000011001001011001",
			3211 => "0000000011001001011001",
			3212 => "0001111000100000000100",
			3213 => "0000000011001001011001",
			3214 => "0001110000111100000100",
			3215 => "0000000011001001011001",
			3216 => "0000000011001001011001",
			3217 => "0011100110111000000100",
			3218 => "0000000011001001011001",
			3219 => "0000000100010100000100",
			3220 => "0000000011001001011001",
			3221 => "0000000011001001011001",
			3222 => "0011100011101000110000",
			3223 => "0000001011111100101100",
			3224 => "0011101001011100011000",
			3225 => "0010010101010100001000",
			3226 => "0000001110100000000100",
			3227 => "0000000011001011101101",
			3228 => "0000000011001011101101",
			3229 => "0011010110110100001000",
			3230 => "0010001001001100000100",
			3231 => "0000000011001011101101",
			3232 => "0000000011001011101101",
			3233 => "0010000011010000000100",
			3234 => "0000000011001011101101",
			3235 => "1111111011001011101101",
			3236 => "0010001001000100001000",
			3237 => "0000111011111000000100",
			3238 => "0000001011001011101101",
			3239 => "0000000011001011101101",
			3240 => "0000001000011100001000",
			3241 => "0000100011111100000100",
			3242 => "0000000011001011101101",
			3243 => "0000000011001011101101",
			3244 => "1111111011001011101101",
			3245 => "1111111011001011101101",
			3246 => "0010001111001000010000",
			3247 => "0000111100110000001000",
			3248 => "0010111011101100000100",
			3249 => "0000000011001011101101",
			3250 => "0000001011001011101101",
			3251 => "0011100100000100000100",
			3252 => "0000000011001011101101",
			3253 => "0000000011001011101101",
			3254 => "0011111101001100001000",
			3255 => "0010001100110000000100",
			3256 => "0000000011001011101101",
			3257 => "0000000011001011101101",
			3258 => "1111111011001011101101",
			3259 => "0011100011101000110100",
			3260 => "0000000011011100011100",
			3261 => "0011100011010100011000",
			3262 => "0000010111110000010000",
			3263 => "0011111111110000000100",
			3264 => "0000000011001110001001",
			3265 => "0000001110000100000100",
			3266 => "0000000011001110001001",
			3267 => "0010110101010100000100",
			3268 => "0000000011001110001001",
			3269 => "0000000011001110001001",
			3270 => "0010001001001100000100",
			3271 => "0000000011001110001001",
			3272 => "1111111011001110001001",
			3273 => "0000000011001110001001",
			3274 => "0000010000011000001000",
			3275 => "0010111010100100000100",
			3276 => "0000000011001110001001",
			3277 => "0000000011001110001001",
			3278 => "0010000101011100001100",
			3279 => "0010001001001100000100",
			3280 => "0000000011001110001001",
			3281 => "0011110110011000000100",
			3282 => "0000000011001110001001",
			3283 => "0000000011001110001001",
			3284 => "1111111011001110001001",
			3285 => "0000111100110000001000",
			3286 => "0000001011001100000100",
			3287 => "0000000011001110001001",
			3288 => "0000000011001110001001",
			3289 => "0000111000101000001000",
			3290 => "0010000101101100000100",
			3291 => "0000000011001110001001",
			3292 => "1111111011001110001001",
			3293 => "0011100100000100001000",
			3294 => "0000100110101000000100",
			3295 => "0000001011001110001001",
			3296 => "0000000011001110001001",
			3297 => "0000000011001110001001",
			3298 => "0001100010001000001100",
			3299 => "0010010111011100001000",
			3300 => "0011011101000000000100",
			3301 => "1111111011010000010101",
			3302 => "0000001011010000010101",
			3303 => "1111111011010000010101",
			3304 => "0000000010100100101000",
			3305 => "0010000101101100010100",
			3306 => "0001111100010000000100",
			3307 => "1111111011010000010101",
			3308 => "0010101011111000001100",
			3309 => "0011101100011000001000",
			3310 => "0000000101000100000100",
			3311 => "0000001011010000010101",
			3312 => "0000000011010000010101",
			3313 => "0000001011010000010101",
			3314 => "0000000011010000010101",
			3315 => "0011100010110000001000",
			3316 => "0000010111100100000100",
			3317 => "0000000011010000010101",
			3318 => "1111111011010000010101",
			3319 => "0000101011100000000100",
			3320 => "0000001011010000010101",
			3321 => "0000111000101000000100",
			3322 => "0000000011010000010101",
			3323 => "0000001011010000010101",
			3324 => "0001101011010100001100",
			3325 => "0000010111100100001000",
			3326 => "0011100110111000000100",
			3327 => "1111111011010000010101",
			3328 => "0000001011010000010101",
			3329 => "1111111011010000010101",
			3330 => "0000111001010100000100",
			3331 => "0000001011010000010101",
			3332 => "1111111011010000010101",
			3333 => "0001100010001000001100",
			3334 => "0010010101010100001000",
			3335 => "0000110111011100000100",
			3336 => "1111111011010010000001",
			3337 => "0000001011010010000001",
			3338 => "1111111011010010000001",
			3339 => "0000001101111000101000",
			3340 => "0011101100011000010000",
			3341 => "0000011000011000001100",
			3342 => "0000100111111100001000",
			3343 => "0001011100110000000100",
			3344 => "0000001011010010000001",
			3345 => "1111111011010010000001",
			3346 => "1111111011010010000001",
			3347 => "1111111011010010000001",
			3348 => "0011010101011100010100",
			3349 => "0011011010100100001100",
			3350 => "0010000101101100001000",
			3351 => "0010000101011100000100",
			3352 => "0000000011010010000001",
			3353 => "0000001011010010000001",
			3354 => "0000000011010010000001",
			3355 => "0000111001010000000100",
			3356 => "0000001011010010000001",
			3357 => "0000001011010010000001",
			3358 => "1111111011010010000001",
			3359 => "1111111011010010000001",
			3360 => "0010011010000100110100",
			3361 => "0011101111111000001100",
			3362 => "0010110110001100001000",
			3363 => "0001111001001000000100",
			3364 => "1111111011010011111101",
			3365 => "0000000011010011111101",
			3366 => "1111111011010011111101",
			3367 => "0000000011001100100000",
			3368 => "0011100010110000010000",
			3369 => "0000011000011000001100",
			3370 => "0000101000100100001000",
			3371 => "0001010011000000000100",
			3372 => "0000001011010011111101",
			3373 => "0000001011010011111101",
			3374 => "1111111011010011111101",
			3375 => "1111111011010011111101",
			3376 => "0000111100110000001100",
			3377 => "0010001001000100001000",
			3378 => "0000000011100000000100",
			3379 => "0000001011010011111101",
			3380 => "0000010011010011111101",
			3381 => "0000001011010011111101",
			3382 => "0000001011010011111101",
			3383 => "0001101011010100000100",
			3384 => "1111111011010011111101",
			3385 => "0000001011010011111101",
			3386 => "0011001100101000001000",
			3387 => "0001011100110000000100",
			3388 => "0000000011010011111101",
			3389 => "1111111011010011111101",
			3390 => "1111111011010011111101",
			3391 => "0011100011101000110100",
			3392 => "0000001011111100110000",
			3393 => "0011101001011100011000",
			3394 => "0010010101010100001000",
			3395 => "0000001110100000000100",
			3396 => "0000000011010110011001",
			3397 => "0000000011010110011001",
			3398 => "0011010110110100001000",
			3399 => "0010001001001100000100",
			3400 => "0000000011010110011001",
			3401 => "0000000011010110011001",
			3402 => "0000011000111100000100",
			3403 => "0000000011010110011001",
			3404 => "1111111011010110011001",
			3405 => "0010001001000100001100",
			3406 => "0000111011111000001000",
			3407 => "0001111001010100000100",
			3408 => "0000000011010110011001",
			3409 => "0000001011010110011001",
			3410 => "0000000011010110011001",
			3411 => "0000001000011100001000",
			3412 => "0000100011111100000100",
			3413 => "0000000011010110011001",
			3414 => "0000000011010110011001",
			3415 => "1111111011010110011001",
			3416 => "1111111011010110011001",
			3417 => "0010001111001000010000",
			3418 => "0001000111011100001000",
			3419 => "0001011111011000000100",
			3420 => "0000001011010110011001",
			3421 => "0000000011010110011001",
			3422 => "0000011001100000000100",
			3423 => "0000000011010110011001",
			3424 => "0000001011010110011001",
			3425 => "0011111101001100001000",
			3426 => "0010001100110000000100",
			3427 => "0000000011010110011001",
			3428 => "0000000011010110011001",
			3429 => "1111111011010110011001",
			3430 => "0001111001010000011100",
			3431 => "0001011101101000010000",
			3432 => "0010100101101100000100",
			3433 => "0000000011011001001101",
			3434 => "0000001110000100001000",
			3435 => "0000001110100000000100",
			3436 => "0000000011011001001101",
			3437 => "0000000011011001001101",
			3438 => "0000000011011001001101",
			3439 => "0000111001000100000100",
			3440 => "0000000011011001001101",
			3441 => "0001001010100100000100",
			3442 => "0000000011011001001101",
			3443 => "0000000011011001001101",
			3444 => "0010101111101000011100",
			3445 => "0001011100010000010000",
			3446 => "0011010101010100001100",
			3447 => "0011011110011000001000",
			3448 => "0001100100001000000100",
			3449 => "0000000011011001001101",
			3450 => "0000000011011001001101",
			3451 => "0000000011011001001101",
			3452 => "0000000011011001001101",
			3453 => "0011111000001000001000",
			3454 => "0001101000110100000100",
			3455 => "0000000011011001001101",
			3456 => "0000000011011001001101",
			3457 => "0000000011011001001101",
			3458 => "0000010111100100001000",
			3459 => "0001011010011100000100",
			3460 => "0000000011011001001101",
			3461 => "0000000011011001001101",
			3462 => "0011100101001100010000",
			3463 => "0001001111011000001000",
			3464 => "0011110000000100000100",
			3465 => "0000000011011001001101",
			3466 => "0000000011011001001101",
			3467 => "0011111000100100000100",
			3468 => "0000000011011001001101",
			3469 => "0000000011011001001101",
			3470 => "0011101000010100001000",
			3471 => "0000111111101000000100",
			3472 => "0000000011011001001101",
			3473 => "0000000011011001001101",
			3474 => "0000000011011001001101",
			3475 => "0011101111010100101000",
			3476 => "0000011000011000100100",
			3477 => "0001001101101000011100",
			3478 => "0001111100010000010000",
			3479 => "0001011100101000001100",
			3480 => "0001111000000100000100",
			3481 => "0000000011011011110001",
			3482 => "0001011011101100000100",
			3483 => "0000000011011011110001",
			3484 => "0000000011011011110001",
			3485 => "0000000011011011110001",
			3486 => "0000001010101000001000",
			3487 => "0001100010001000000100",
			3488 => "0000000011011011110001",
			3489 => "0000000011011011110001",
			3490 => "0000000011011011110001",
			3491 => "0001010110101100000100",
			3492 => "0000000011011011110001",
			3493 => "0000000011011011110001",
			3494 => "0000000011011011110001",
			3495 => "0010101111101000011000",
			3496 => "0001011100010000010000",
			3497 => "0011011110011000001100",
			3498 => "0011001110011000001000",
			3499 => "0000100000000000000100",
			3500 => "0000000011011011110001",
			3501 => "0000000011011011110001",
			3502 => "0000000011011011110001",
			3503 => "0000001011011011110001",
			3504 => "0001100000001100000100",
			3505 => "0000000011011011110001",
			3506 => "0000000011011011110001",
			3507 => "0001011001010000001000",
			3508 => "0001111100101100000100",
			3509 => "0000000011011011110001",
			3510 => "0000000011011011110001",
			3511 => "0010011010000100001000",
			3512 => "0000001110110000000100",
			3513 => "0000000011011011110001",
			3514 => "0000000011011011110001",
			3515 => "0000000011011011110001",
			3516 => "0011101101100100110000",
			3517 => "0001011100101000001000",
			3518 => "0000001110100000000100",
			3519 => "0000000011011110010101",
			3520 => "0000000011011110010101",
			3521 => "0001111111101000100000",
			3522 => "0011101111010100011000",
			3523 => "0001011101101000010000",
			3524 => "0001010101101100001000",
			3525 => "0001001011101100000100",
			3526 => "0000000011011110010101",
			3527 => "0000000011011110010101",
			3528 => "0001001011101100000100",
			3529 => "0000000011011110010101",
			3530 => "0000000011011110010101",
			3531 => "0001000011010000000100",
			3532 => "0000000011011110010101",
			3533 => "0000000011011110010101",
			3534 => "0001001010000100000100",
			3535 => "0000000011011110010101",
			3536 => "0000000011011110010101",
			3537 => "0001000110000000000100",
			3538 => "0000000011011110010101",
			3539 => "0000000011011110010101",
			3540 => "0000000011001100001100",
			3541 => "0001011000000000000100",
			3542 => "0000000011011110010101",
			3543 => "0001011101001000000100",
			3544 => "0000000011011110010101",
			3545 => "0000000011011110010101",
			3546 => "0001100000100100010000",
			3547 => "0000111111101000001000",
			3548 => "0000110011001000000100",
			3549 => "0000000011011110010101",
			3550 => "0000000011011110010101",
			3551 => "0010101001011000000100",
			3552 => "0000000011011110010101",
			3553 => "0000000011011110010101",
			3554 => "0000111001010100000100",
			3555 => "0000000011011110010101",
			3556 => "0000000011011110010101",
			3557 => "0001100010001000001100",
			3558 => "0010010111011100001000",
			3559 => "0010110110110100000100",
			3560 => "0000000011100000001001",
			3561 => "0000000011100000001001",
			3562 => "1111111011100000001001",
			3563 => "0000001101111000101100",
			3564 => "0001011111011000001100",
			3565 => "0010011100101000001000",
			3566 => "0010100011000000000100",
			3567 => "0000000011100000001001",
			3568 => "0000001011100000001001",
			3569 => "0000000011100000001001",
			3570 => "0001110001010000001100",
			3571 => "0000000111000100001000",
			3572 => "0001111101001000000100",
			3573 => "1111111011100000001001",
			3574 => "0000000011100000001001",
			3575 => "1111111011100000001001",
			3576 => "0000010111110000000100",
			3577 => "0000001011100000001001",
			3578 => "0000101011100000001000",
			3579 => "0011100011010100000100",
			3580 => "0000000011100000001001",
			3581 => "0000001011100000001001",
			3582 => "0001100100001000000100",
			3583 => "1111111011100000001001",
			3584 => "0000000011100000001001",
			3585 => "1111111011100000001001",
			3586 => "0010000101101100100100",
			3587 => "0001101101000100000100",
			3588 => "0000000011100010100101",
			3589 => "0000001101111000011100",
			3590 => "0001000101011100001000",
			3591 => "0010000011010000000100",
			3592 => "0000000011100010100101",
			3593 => "0000000011100010100101",
			3594 => "0000111100110000001000",
			3595 => "0001110110101100000100",
			3596 => "0000000011100010100101",
			3597 => "0000000011100010100101",
			3598 => "0010010110000000000100",
			3599 => "0000000011100010100101",
			3600 => "0010000101011100000100",
			3601 => "0000000011100010100101",
			3602 => "0000000011100010100101",
			3603 => "0000000011100010100101",
			3604 => "0011110100110100100000",
			3605 => "0000101011101000010100",
			3606 => "0001110001010000001100",
			3607 => "0001001110011000001000",
			3608 => "0001001011101100000100",
			3609 => "0000000011100010100101",
			3610 => "0000000011100010100101",
			3611 => "0000000011100010100101",
			3612 => "0010010011000000000100",
			3613 => "0000000011100010100101",
			3614 => "0000000011100010100101",
			3615 => "0000111100101100000100",
			3616 => "0000000011100010100101",
			3617 => "0001001100110000000100",
			3618 => "0000000011100010100101",
			3619 => "0000000011100010100101",
			3620 => "0001000101010100000100",
			3621 => "0000000011100010100101",
			3622 => "0000011101000000000100",
			3623 => "0000000011100010100101",
			3624 => "0000000011100010100101",
			3625 => "0011110011010100001100",
			3626 => "0010110110001100001000",
			3627 => "0010111101000000000100",
			3628 => "1111111011100100110001",
			3629 => "0000000011100100110001",
			3630 => "1111111011100100110001",
			3631 => "0000000011001100101000",
			3632 => "0001010011110100100100",
			3633 => "0001000111011100001100",
			3634 => "0011001110011000000100",
			3635 => "0000001011100100110001",
			3636 => "0000000101011000000100",
			3637 => "0000001011100100110001",
			3638 => "0000001011100100110001",
			3639 => "0001110001010000001100",
			3640 => "0011011110011000001000",
			3641 => "0000000111000100000100",
			3642 => "0000001011100100110001",
			3643 => "1111111011100100110001",
			3644 => "1111111011100100110001",
			3645 => "0011010101011100001000",
			3646 => "0000010111100100000100",
			3647 => "0000001011100100110001",
			3648 => "0000001011100100110001",
			3649 => "1111111011100100110001",
			3650 => "1111111011100100110001",
			3651 => "0001101011010100001100",
			3652 => "0011010110110100001000",
			3653 => "0001011001010000000100",
			3654 => "1111111011100100110001",
			3655 => "0000001011100100110001",
			3656 => "1111111011100100110001",
			3657 => "0000111100110000000100",
			3658 => "0000001011100100110001",
			3659 => "1111111011100100110001",
			3660 => "0011101100011000110100",
			3661 => "0001000101011100011100",
			3662 => "0000010110010000010000",
			3663 => "0001101101000100000100",
			3664 => "0000000011100111010101",
			3665 => "0000001110000100000100",
			3666 => "0000001011100111010101",
			3667 => "0010010101011100000100",
			3668 => "0000000011100111010101",
			3669 => "0000000011100111010101",
			3670 => "0001111101001000000100",
			3671 => "0000000011100111010101",
			3672 => "0010101010000100000100",
			3673 => "0000000011100111010101",
			3674 => "0000000011100111010101",
			3675 => "0001111100101100010000",
			3676 => "0000110011000000001100",
			3677 => "0000111101101000001000",
			3678 => "0001010101111000000100",
			3679 => "0000000011100111010101",
			3680 => "0000000011100111010101",
			3681 => "0000000011100111010101",
			3682 => "1111111011100111010101",
			3683 => "0001011100010000000100",
			3684 => "0000000011100111010101",
			3685 => "0000000011100111010101",
			3686 => "0000001101111000011100",
			3687 => "0001011111011000000100",
			3688 => "0000001011100111010101",
			3689 => "0001011000000100000100",
			3690 => "0000000011100111010101",
			3691 => "0000100011011100000100",
			3692 => "0000001011100111010101",
			3693 => "0000111000101000001000",
			3694 => "0011101000110100000100",
			3695 => "0000000011100111010101",
			3696 => "0000000011100111010101",
			3697 => "0001100100001000000100",
			3698 => "0000000011100111010101",
			3699 => "0000001011100111010101",
			3700 => "1111111011100111010101",
			3701 => "0011111111110000000100",
			3702 => "1111111011101001000001",
			3703 => "0001010001010000101000",
			3704 => "0000001101111000100100",
			3705 => "0000010111110000010000",
			3706 => "0000101001110100001000",
			3707 => "0010111011101100000100",
			3708 => "0000000011101001000001",
			3709 => "0000001011101001000001",
			3710 => "0001011000000100000100",
			3711 => "0000000011101001000001",
			3712 => "1111111011101001000001",
			3713 => "0011100100001100001000",
			3714 => "0000011000011000000100",
			3715 => "0000000011101001000001",
			3716 => "1111111011101001000001",
			3717 => "0000000011011100000100",
			3718 => "0000001011101001000001",
			3719 => "0001100100001000000100",
			3720 => "1111111011101001000001",
			3721 => "0000000011101001000001",
			3722 => "1111111011101001000001",
			3723 => "0011100110000100000100",
			3724 => "1111111011101001000001",
			3725 => "0011111101001100000100",
			3726 => "0000001011101001000001",
			3727 => "1111111011101001000001",
			3728 => "0011000110001100001000",
			3729 => "0010001111111100000100",
			3730 => "0000000011101011010101",
			3731 => "0000001011101011010101",
			3732 => "0001011010000100010000",
			3733 => "0001101111000100001000",
			3734 => "0010111011101100000100",
			3735 => "0000000011101011010101",
			3736 => "1111111011101011010101",
			3737 => "0010111011101100000100",
			3738 => "0000000011101011010101",
			3739 => "0000001011101011010101",
			3740 => "0001111001010000010000",
			3741 => "0001000011010000000100",
			3742 => "0000000011101011010101",
			3743 => "0010001010100100000100",
			3744 => "0000000011101011010101",
			3745 => "0010101111011000000100",
			3746 => "0000000011101011010101",
			3747 => "1111111011101011010101",
			3748 => "0000000011001100010100",
			3749 => "0010101011111000001100",
			3750 => "0001010011001000000100",
			3751 => "0000000011101011010101",
			3752 => "0000100011011100000100",
			3753 => "0000001011101011010101",
			3754 => "0000000011101011010101",
			3755 => "0000010111110000000100",
			3756 => "0000000011101011010101",
			3757 => "1111111011101011010101",
			3758 => "0000010111100100001000",
			3759 => "0011011011101100000100",
			3760 => "0000000011101011010101",
			3761 => "0000000011101011010101",
			3762 => "0000110011100100000100",
			3763 => "0000000011101011010101",
			3764 => "1111111011101011010101",
			3765 => "0011000110001100001000",
			3766 => "0010001111111100000100",
			3767 => "0000000011101101110001",
			3768 => "0000001011101101110001",
			3769 => "0001011010000100010000",
			3770 => "0001101111000100001000",
			3771 => "0010111011101100000100",
			3772 => "0000000011101101110001",
			3773 => "0000000011101101110001",
			3774 => "0010111011101100000100",
			3775 => "0000000011101101110001",
			3776 => "0000001011101101110001",
			3777 => "0001111001010000010000",
			3778 => "0001000011010000000100",
			3779 => "0000000011101101110001",
			3780 => "0010001010100100000100",
			3781 => "0000000011101101110001",
			3782 => "0010101111011000000100",
			3783 => "0000000011101101110001",
			3784 => "1111111011101101110001",
			3785 => "0000000011001100011000",
			3786 => "0010101011111000010000",
			3787 => "0011011010100100001000",
			3788 => "0010001111111100000100",
			3789 => "0000001011101101110001",
			3790 => "0000000011101101110001",
			3791 => "0011100010110000000100",
			3792 => "0000000011101101110001",
			3793 => "0000001011101101110001",
			3794 => "0000010111110000000100",
			3795 => "0000000011101101110001",
			3796 => "1111111011101101110001",
			3797 => "0000010111100100001000",
			3798 => "0000000101101000000100",
			3799 => "0000000011101101110001",
			3800 => "0000000011101101110001",
			3801 => "0000110011100100000100",
			3802 => "0000000011101101110001",
			3803 => "1111111011101101110001",
			3804 => "0011111111110000000100",
			3805 => "1111111011101111010111",
			3806 => "0000001101111000101100",
			3807 => "0001010011110100101000",
			3808 => "0000010111100100010100",
			3809 => "0000100011011100001000",
			3810 => "0001011000000000000100",
			3811 => "0000001011101111010111",
			3812 => "0000001011101111010111",
			3813 => "0010101001010100000100",
			3814 => "1111111011101111010111",
			3815 => "0011100111001000000100",
			3816 => "1111111011101111010111",
			3817 => "0000001011101111010111",
			3818 => "0011101100011000001000",
			3819 => "0001111011111000000100",
			3820 => "1111111011101111010111",
			3821 => "0000000011101111010111",
			3822 => "0001011111011000000100",
			3823 => "0000001011101111010111",
			3824 => "0000000011111000000100",
			3825 => "0000001011101111010111",
			3826 => "0000000011101111010111",
			3827 => "1111111011101111010111",
			3828 => "1111111011101111010111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1331, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2571, initial_addr_3'length));
	end generate gen_rom_1;

	gen_rom_2: if SELECT_ROM = 2 generate
		bank <= (
			0 => "0010011001000100101100",
			1 => "0000001111101100010000",
			2 => "0010101001011000001100",
			3 => "0010101111101000000100",
			4 => "1100111000000001111101",
			5 => "0000010111110000000100",
			6 => "1101010000000001111101",
			7 => "1100111000000001111101",
			8 => "1101101000000001111101",
			9 => "0001011000111000001100",
			10 => "0001011000000100000100",
			11 => "1100111000000001111101",
			12 => "0010001111111100000100",
			13 => "1101110000000001111101",
			14 => "1100111000000001111101",
			15 => "0000010111100100001000",
			16 => "0001011101001000000100",
			17 => "1110011000000001111101",
			18 => "1110111000000001111101",
			19 => "0011110010101000000100",
			20 => "1101111000000001111101",
			21 => "1100111000000001111101",
			22 => "0011001100101000010000",
			23 => "0010101001000000000100",
			24 => "1100111000000001111101",
			25 => "0000010110010000001000",
			26 => "0001101111000100000100",
			27 => "1100111000000001111101",
			28 => "1101000000000001111101",
			29 => "1101011000000001111101",
			30 => "1100111000000001111101",
			31 => "0010010101101100101000",
			32 => "0001011000000000001100",
			33 => "0010001010100100000100",
			34 => "0000000000000100000001",
			35 => "0000111100110000000100",
			36 => "0000000000000100000001",
			37 => "0000000000000100000001",
			38 => "0011001110011000001000",
			39 => "0001100101001100000100",
			40 => "0000000000000100000001",
			41 => "0000000000000100000001",
			42 => "0000011000011000010000",
			43 => "0000001011111100000100",
			44 => "0000000000000100000001",
			45 => "0001100101001100000100",
			46 => "0000000000000100000001",
			47 => "0011111011010100000100",
			48 => "0000000000000100000001",
			49 => "0000000000000100000001",
			50 => "0000000000000100000001",
			51 => "0010001001001100001000",
			52 => "0011111001011100000100",
			53 => "0000000000000100000001",
			54 => "0000000000000100000001",
			55 => "0011100010001100001000",
			56 => "0000000100110000000100",
			57 => "0000000000000100000001",
			58 => "0000000000000100000001",
			59 => "0010101100110100000100",
			60 => "0000000000000100000001",
			61 => "0010100000111000000100",
			62 => "0000000000000100000001",
			63 => "0000000000000100000001",
			64 => "0010011001000100101000",
			65 => "0000001101110100001000",
			66 => "0000111111101000000100",
			67 => "1111111000000101110101",
			68 => "0000000000000101110101",
			69 => "0001011000000000001000",
			70 => "0001001100101000000100",
			71 => "1111111000000101110101",
			72 => "0000000000000101110101",
			73 => "0000011000011000010000",
			74 => "0010000101101100001100",
			75 => "0011111110101100000100",
			76 => "0000101000000101110101",
			77 => "0000100111111000000100",
			78 => "0000010000000101110101",
			79 => "0000100000000101110101",
			80 => "0000001000000101110101",
			81 => "0001111111101000000100",
			82 => "1111111000000101110101",
			83 => "0000000000000101110101",
			84 => "0011001100101000010000",
			85 => "0010101001000000000100",
			86 => "1111111000000101110101",
			87 => "0001011001101100001000",
			88 => "0001101010011000000100",
			89 => "0000000000000101110101",
			90 => "0000011000000101110101",
			91 => "1111111000000101110101",
			92 => "1111111000000101110101",
			93 => "0010011001000100100000",
			94 => "0000000111101100000100",
			95 => "1111111000000111011001",
			96 => "0011100001000000011000",
			97 => "0001011000000100000100",
			98 => "1111111000000111011001",
			99 => "0010101011111000001100",
			100 => "0010000101101100001000",
			101 => "0000101101110000000100",
			102 => "0000000000000111011001",
			103 => "0000001000000111011001",
			104 => "1111111000000111011001",
			105 => "0011010110001100000100",
			106 => "0000001000000111011001",
			107 => "0000001000000111011001",
			108 => "1111111000000111011001",
			109 => "0011001100101000010000",
			110 => "0010101001000000000100",
			111 => "1111111000000111011001",
			112 => "0000010110010000001000",
			113 => "0001001100001100000100",
			114 => "1111111000000111011001",
			115 => "0000001000000111011001",
			116 => "0000001000000111011001",
			117 => "1111111000000111011001",
			118 => "0010011001000100110000",
			119 => "0000001101110100001100",
			120 => "0000000111101100000100",
			121 => "1111111000001001011101",
			122 => "0000001011001000000100",
			123 => "0000000000001001011101",
			124 => "1111111000001001011101",
			125 => "0001001001000100010000",
			126 => "0000111000000000001000",
			127 => "0000101111001100000100",
			128 => "1111111000001001011101",
			129 => "0000000000001001011101",
			130 => "0011101110010000000100",
			131 => "0000010000001001011101",
			132 => "1111111000001001011101",
			133 => "0011100111100000010000",
			134 => "0000101001110100000100",
			135 => "0000100000001001011101",
			136 => "0010000101101100001000",
			137 => "0001001010000100000100",
			138 => "0000010000001001011101",
			139 => "0000010000001001011101",
			140 => "0000001000001001011101",
			141 => "1111111000001001011101",
			142 => "0010110101010100010000",
			143 => "0010101001000000000100",
			144 => "1111111000001001011101",
			145 => "0001000110011100000100",
			146 => "0000010000001001011101",
			147 => "0001001100001100000100",
			148 => "1111111000001001011101",
			149 => "0000000000001001011101",
			150 => "1111111000001001011101",
			151 => "0011001100101000101000",
			152 => "0001100101001000001100",
			153 => "0010000101101100000100",
			154 => "1111111000001010110001",
			155 => "0011011011101100000100",
			156 => "0000001000001010110001",
			157 => "1111111000001010110001",
			158 => "0011100001000000011000",
			159 => "0001011000000100000100",
			160 => "1111111000001010110001",
			161 => "0011010011010000010000",
			162 => "0010101011111000001000",
			163 => "0010010101101100000100",
			164 => "0000000000001010110001",
			165 => "1111111000001010110001",
			166 => "0001011001101100000100",
			167 => "0000001000001010110001",
			168 => "1111111000001010110001",
			169 => "1111111000001010110001",
			170 => "1111111000001010110001",
			171 => "1111111000001010110001",
			172 => "0001110110101100011100",
			173 => "0000100010100100010100",
			174 => "0010101001000000001000",
			175 => "0010001010100100000100",
			176 => "0000000000001101000101",
			177 => "0000000000001101000101",
			178 => "0000000100110000000100",
			179 => "0000000000001101000101",
			180 => "0001011001101100000100",
			181 => "0000000000001101000101",
			182 => "0000000000001101000101",
			183 => "0000010111110000000100",
			184 => "0000000000001101000101",
			185 => "0000000000001101000101",
			186 => "0000101101110000101000",
			187 => "0001101000110100010100",
			188 => "0011111110001000001100",
			189 => "0000011001100000000100",
			190 => "0000000000001101000101",
			191 => "0000010001100100000100",
			192 => "0000000000001101000101",
			193 => "0000000000001101000101",
			194 => "0000011000011000000100",
			195 => "0000000000001101000101",
			196 => "0000000000001101000101",
			197 => "0001111001010000000100",
			198 => "0000000000001101000101",
			199 => "0001110100101100001100",
			200 => "0010001111001000001000",
			201 => "0001001001000100000100",
			202 => "0000000000001101000101",
			203 => "0000000000001101000101",
			204 => "0000000000001101000101",
			205 => "0000000000001101000101",
			206 => "0001111000101000000100",
			207 => "0000000000001101000101",
			208 => "0000000000001101000101",
			209 => "0011100110110000111100",
			210 => "0000001101110000101000",
			211 => "0010010101011100001100",
			212 => "0010001001001100000100",
			213 => "0000000000001111100001",
			214 => "0010001111111100000100",
			215 => "0000000000001111100001",
			216 => "0000000000001111100001",
			217 => "0011001010100100001000",
			218 => "0010101001010100000100",
			219 => "0000000000001111100001",
			220 => "0000000000001111100001",
			221 => "0000000100010100010000",
			222 => "0010101100001100001000",
			223 => "0011100010001100000100",
			224 => "0000000000001111100001",
			225 => "0000000000001111100001",
			226 => "0001011001101100000100",
			227 => "0000000000001111100001",
			228 => "0000000000001111100001",
			229 => "0000000000001111100001",
			230 => "0011011011101100001100",
			231 => "0010000101011100001000",
			232 => "0011111011000100000100",
			233 => "0000000000001111100001",
			234 => "0000000000001111100001",
			235 => "0000000000001111100001",
			236 => "0011111011110100000100",
			237 => "0000000000001111100001",
			238 => "0000000000001111100001",
			239 => "0010111011101100001000",
			240 => "0010101000101000000100",
			241 => "0000000000001111100001",
			242 => "0000000000001111100001",
			243 => "0000010110010000000100",
			244 => "0000000000001111100001",
			245 => "0000011000011000000100",
			246 => "0000000000001111100001",
			247 => "0000000000001111100001",
			248 => "0010000101101100101100",
			249 => "0000101101110000100100",
			250 => "0000100000101000100000",
			251 => "0000001101110000011000",
			252 => "0010111010100100001100",
			253 => "0011010011110000000100",
			254 => "0000000000010001100101",
			255 => "0010101011111000000100",
			256 => "0000000000010001100101",
			257 => "0000000000010001100101",
			258 => "0000001011111100001000",
			259 => "0000110000111100000100",
			260 => "0000000000010001100101",
			261 => "0000000000010001100101",
			262 => "0000000000010001100101",
			263 => "0001001101101000000100",
			264 => "0000000000010001100101",
			265 => "0000000000010001100101",
			266 => "0000000000010001100101",
			267 => "0001011000000000000100",
			268 => "0000000000010001100101",
			269 => "0000000000010001100101",
			270 => "0000111011111000001000",
			271 => "0001011110111000000100",
			272 => "0000000000010001100101",
			273 => "0000000000010001100101",
			274 => "0011001100101000001100",
			275 => "0010101001011000000100",
			276 => "0000000000010001100101",
			277 => "0000010110010000000100",
			278 => "0000000000010001100101",
			279 => "0000000000010001100101",
			280 => "0000000000010001100101",
			281 => "0010011001000100110100",
			282 => "0000001101110100001100",
			283 => "0000000111101100000100",
			284 => "1111111000010011110001",
			285 => "0011001010100100000100",
			286 => "0000000000010011110001",
			287 => "1111111000010011110001",
			288 => "0001001001000100010000",
			289 => "0000111000000000001000",
			290 => "0000101111001100000100",
			291 => "1111111000010011110001",
			292 => "0000000000010011110001",
			293 => "0011111011011000000100",
			294 => "0000010000010011110001",
			295 => "1111111000010011110001",
			296 => "0011100111100000010100",
			297 => "0010000101101100010000",
			298 => "0001001010000100001000",
			299 => "0011111011110100000100",
			300 => "0000001000010011110001",
			301 => "0000010000010011110001",
			302 => "0011110010111100000100",
			303 => "0000010000010011110001",
			304 => "0000010000010011110001",
			305 => "0000001000010011110001",
			306 => "1111111000010011110001",
			307 => "0010110101010100010000",
			308 => "0010101001000000000100",
			309 => "1111111000010011110001",
			310 => "0000010110010000001000",
			311 => "0001001100001100000100",
			312 => "1111111000010011110001",
			313 => "0000000000010011110001",
			314 => "0000001000010011110001",
			315 => "1111111000010011110001",
			316 => "0011011011101100110000",
			317 => "0011100110110000101000",
			318 => "0000001101110000100000",
			319 => "0010101011111000010000",
			320 => "0010110110001100000100",
			321 => "0000000000010110000101",
			322 => "0010110011010000001000",
			323 => "0001000101010100000100",
			324 => "0000000000010110000101",
			325 => "0000000000010110000101",
			326 => "0000000000010110000101",
			327 => "0010011010000100001100",
			328 => "0001100100000000000100",
			329 => "0000000000010110000101",
			330 => "0001011001101100000100",
			331 => "0000000000010110000101",
			332 => "0000000000010110000101",
			333 => "0000000000010110000101",
			334 => "0000010111110000000100",
			335 => "0000000000010110000101",
			336 => "0000000000010110000101",
			337 => "0010111011101100000100",
			338 => "0000000000010110000101",
			339 => "0000000000010110000101",
			340 => "0010001001001100001000",
			341 => "0011110101001100000100",
			342 => "0000000000010110000101",
			343 => "0000000000010110000101",
			344 => "0010101100110100001100",
			345 => "0010111110011000001000",
			346 => "0011001110011000000100",
			347 => "0000000000010110000101",
			348 => "0000000000010110000101",
			349 => "0000000000010110000101",
			350 => "0000110011110100000100",
			351 => "0000000000010110000101",
			352 => "0000000000010110000101",
			353 => "0011100110110001000000",
			354 => "0011001110011000010000",
			355 => "0001100101001100001100",
			356 => "0001001010000100001000",
			357 => "0010001010100100000100",
			358 => "0000000000011000101001",
			359 => "0000000000011000101001",
			360 => "0000000000011000101001",
			361 => "0000000000011000101001",
			362 => "0000001101110100010100",
			363 => "0001010001111100001100",
			364 => "0011100010001100001000",
			365 => "0000000100110000000100",
			366 => "0000000000011000101001",
			367 => "0000000000011000101001",
			368 => "0000000000011000101001",
			369 => "0001011001101100000100",
			370 => "0000000000011000101001",
			371 => "0000000000011000101001",
			372 => "0000010110010000001100",
			373 => "0001001100010000001000",
			374 => "0011111000001000000100",
			375 => "0000000000011000101001",
			376 => "0000000000011000101001",
			377 => "0000000000011000101001",
			378 => "0001011111101000001000",
			379 => "0000000101101000000100",
			380 => "0000000000011000101001",
			381 => "0000000000011000101001",
			382 => "0010010110000000000100",
			383 => "0000000000011000101001",
			384 => "0000000000011000101001",
			385 => "0010111011101100001000",
			386 => "0011110000011100000100",
			387 => "0000000000011000101001",
			388 => "0000000000011000101001",
			389 => "0000010110010000000100",
			390 => "0000000000011000101001",
			391 => "0000011000011000000100",
			392 => "0000000000011000101001",
			393 => "0000000000011000101001",
			394 => "0010010101101100110000",
			395 => "0001011000000000001000",
			396 => "0000111100110000000100",
			397 => "1111111000011010111101",
			398 => "0000000000011010111101",
			399 => "0010000101101100100000",
			400 => "0000011001100100001000",
			401 => "0011110101111100000100",
			402 => "1111111000011010111101",
			403 => "0000000000011010111101",
			404 => "0001011101001000001100",
			405 => "0011110000100100001000",
			406 => "0001110110101100000100",
			407 => "0000000000011010111101",
			408 => "0000000000011010111101",
			409 => "0000001000011010111101",
			410 => "0010101001010100000100",
			411 => "0000000000011010111101",
			412 => "0001100001001100000100",
			413 => "0000000000011010111101",
			414 => "0000001000011010111101",
			415 => "0011110000001000000100",
			416 => "0000000000011010111101",
			417 => "1111111000011010111101",
			418 => "0010101001011000001000",
			419 => "0010001001001100000100",
			420 => "0000000000011010111101",
			421 => "1111111000011010111101",
			422 => "0010010011000000010000",
			423 => "0011101010011000001000",
			424 => "0001101101101100000100",
			425 => "0000001000011010111101",
			426 => "1111111000011010111101",
			427 => "0010001111111100000100",
			428 => "0000000000011010111101",
			429 => "0000001000011010111101",
			430 => "1111111000011010111101",
			431 => "0000100111000100011000",
			432 => "0010101011111000000100",
			433 => "1111111000011101100001",
			434 => "0001001000000000000100",
			435 => "0000001000011101100001",
			436 => "0000011000111100001000",
			437 => "0010000101011100000100",
			438 => "1111111000011101100001",
			439 => "0000001000011101100001",
			440 => "0010001001001100000100",
			441 => "0000000000011101100001",
			442 => "1111111000011101100001",
			443 => "0010000101101100101100",
			444 => "0000111000000000010100",
			445 => "0011010110001100001100",
			446 => "0001001001000100001000",
			447 => "0010010101010100000100",
			448 => "1111111000011101100001",
			449 => "0000000000011101100001",
			450 => "0000001000011101100001",
			451 => "0001111001010100000100",
			452 => "1111111000011101100001",
			453 => "0000000000011101100001",
			454 => "0011100110110000010000",
			455 => "0011001110011000000100",
			456 => "0000001000011101100001",
			457 => "0001100100110000000100",
			458 => "0000001000011101100001",
			459 => "0011111100111100000100",
			460 => "0000001000011101100001",
			461 => "0000001000011101100001",
			462 => "0000101011100100000100",
			463 => "1111111000011101100001",
			464 => "0000001000011101100001",
			465 => "0010101001011000001000",
			466 => "0001111001010000000100",
			467 => "1111111000011101100001",
			468 => "1111111000011101100001",
			469 => "0011101110100100000100",
			470 => "0000001000011101100001",
			471 => "1111111000011101100001",
			472 => "0000010001100100101000",
			473 => "0000011000111100001000",
			474 => "0011010110110100000100",
			475 => "1111111000011110110101",
			476 => "0000000000011110110101",
			477 => "0000110101111000000100",
			478 => "1111111000011110110101",
			479 => "0011100001000000011000",
			480 => "0000000101101000010000",
			481 => "0010101011111000001000",
			482 => "0000010110010000000100",
			483 => "0000000000011110110101",
			484 => "1111111000011110110101",
			485 => "0001011001101100000100",
			486 => "0000001000011110110101",
			487 => "1111111000011110110101",
			488 => "0011011011101100000100",
			489 => "0000001000011110110101",
			490 => "0000000000011110110101",
			491 => "1111111000011110110101",
			492 => "1111111000011110110101",
			493 => "0010101001010100011100",
			494 => "0001111001010000010000",
			495 => "0011101111110100001000",
			496 => "0011110111000000000100",
			497 => "0000000000100001110001",
			498 => "0000000000100001110001",
			499 => "0000000101010000000100",
			500 => "1111111000100001110001",
			501 => "0000000000100001110001",
			502 => "0010111010100100001000",
			503 => "0011100110111000000100",
			504 => "0000000000100001110001",
			505 => "0000000000100001110001",
			506 => "0000000000100001110001",
			507 => "0000011000011000101100",
			508 => "0001100111101000011100",
			509 => "0001110110101100010100",
			510 => "0011101010110100001100",
			511 => "0010000101101100000100",
			512 => "0000000000100001110001",
			513 => "0001101101101100000100",
			514 => "0000000000100001110001",
			515 => "0000000000100001110001",
			516 => "0011010110001100000100",
			517 => "0000000000100001110001",
			518 => "0000000000100001110001",
			519 => "0010100100101100000100",
			520 => "0000000000100001110001",
			521 => "0000000000100001110001",
			522 => "0011101101100100001000",
			523 => "0001011011000000000100",
			524 => "0000001000100001110001",
			525 => "0000000000100001110001",
			526 => "0010111110011000000100",
			527 => "0000000000100001110001",
			528 => "0000000000100001110001",
			529 => "0000001011000100001000",
			530 => "0000100100100000000100",
			531 => "0000000000100001110001",
			532 => "0000000000100001110001",
			533 => "0001111111101000000100",
			534 => "0000000000100001110001",
			535 => "0001111011111000001000",
			536 => "0011110000000100000100",
			537 => "0000000000100001110001",
			538 => "0000000000100001110001",
			539 => "0000000000100001110001",
			540 => "0011100110110000111100",
			541 => "0000001101110000101100",
			542 => "0001011101001000010100",
			543 => "0011000111011100001100",
			544 => "0010110110001100001000",
			545 => "0001100111010100000100",
			546 => "0000000000100100000101",
			547 => "0000001000100100000101",
			548 => "1111111000100100000101",
			549 => "0010010101101100000100",
			550 => "0000001000100100000101",
			551 => "0000000000100100000101",
			552 => "0001000011000100010100",
			553 => "0001010001111100010000",
			554 => "0011101001011100001000",
			555 => "0001111100000000000100",
			556 => "0000000000100100000101",
			557 => "1111111000100100000101",
			558 => "0000111101001000000100",
			559 => "0000000000100100000101",
			560 => "0000001000100100000101",
			561 => "0000001000100100000101",
			562 => "1111111000100100000101",
			563 => "0011010110001100000100",
			564 => "0000001000100100000101",
			565 => "0010101001010100000100",
			566 => "1111111000100100000101",
			567 => "0000010111100100000100",
			568 => "0000001000100100000101",
			569 => "0000000000100100000101",
			570 => "0010011001001000001100",
			571 => "0000000101010000001000",
			572 => "0011111101001100000100",
			573 => "0000000000100100000101",
			574 => "1111111000100100000101",
			575 => "0000000000100100000101",
			576 => "1111111000100100000101",
			577 => "0011011011101100111000",
			578 => "0001001001000100010000",
			579 => "0000111000000000001100",
			580 => "0000111111011000001000",
			581 => "0000110011000000000100",
			582 => "0000000000100110100001",
			583 => "0000000000100110100001",
			584 => "0000000000100110100001",
			585 => "0000000000100110100001",
			586 => "0011111011110100100000",
			587 => "0001110110101100010100",
			588 => "0000010111100100010000",
			589 => "0011000011010000001000",
			590 => "0001111000000100000100",
			591 => "0000000000100110100001",
			592 => "0000000000100110100001",
			593 => "0000111011000000000100",
			594 => "0000000000100110100001",
			595 => "0000000000100110100001",
			596 => "0000000000100110100001",
			597 => "0001000101111000000100",
			598 => "0000000000100110100001",
			599 => "0000000010101100000100",
			600 => "0000000000100110100001",
			601 => "0000000000100110100001",
			602 => "0000010001110000000100",
			603 => "0000000000100110100001",
			604 => "0000000000100110100001",
			605 => "0010001001001100000100",
			606 => "0000000000100110100001",
			607 => "0010111110011000001000",
			608 => "0000111101001000000100",
			609 => "0000000000100110100001",
			610 => "0000000000100110100001",
			611 => "0010101100110100000100",
			612 => "0000000000100110100001",
			613 => "0000110011110100000100",
			614 => "0000000000100110100001",
			615 => "0000000000100110100001",
			616 => "0010101001010100100100",
			617 => "0011111011010100011000",
			618 => "0001010110101100001100",
			619 => "0000111111011000001000",
			620 => "0000110011000000000100",
			621 => "0000000000101001011101",
			622 => "0000000000101001011101",
			623 => "1111111000101001011101",
			624 => "0001001101101000000100",
			625 => "0000000000101001011101",
			626 => "0000110011100100000100",
			627 => "0000000000101001011101",
			628 => "0000000000101001011101",
			629 => "0011100110110000000100",
			630 => "0000000000101001011101",
			631 => "0010111011101100000100",
			632 => "0000000000101001011101",
			633 => "0000000000101001011101",
			634 => "0000101101011100101000",
			635 => "0001010001111100100000",
			636 => "0011101001011100001100",
			637 => "0011100010001100001000",
			638 => "0010000101101100000100",
			639 => "0000000000101001011101",
			640 => "0000000000101001011101",
			641 => "1111111000101001011101",
			642 => "0000101111101100010000",
			643 => "0001111101001000001000",
			644 => "0011100101110100000100",
			645 => "0000000000101001011101",
			646 => "0000000000101001011101",
			647 => "0011011011101100000100",
			648 => "0000000000101001011101",
			649 => "0000000000101001011101",
			650 => "0000000000101001011101",
			651 => "0001011001101100000100",
			652 => "0000000000101001011101",
			653 => "0000000000101001011101",
			654 => "0010000101101100001000",
			655 => "0011101110100000000100",
			656 => "0000001000101001011101",
			657 => "0000000000101001011101",
			658 => "0010100000111100000100",
			659 => "0000000000101001011101",
			660 => "0000111100101100000100",
			661 => "0000000000101001011101",
			662 => "0000000000101001011101",
			663 => "0000010111100100111100",
			664 => "0000011000111100001000",
			665 => "0011010110110100000100",
			666 => "1111111000101100000001",
			667 => "0000000000101100000001",
			668 => "0001100101000000011000",
			669 => "0011010110001100001000",
			670 => "0000010111110000000100",
			671 => "1111111000101100000001",
			672 => "0000000000101100000001",
			673 => "0001000110011100001100",
			674 => "0010101111101000000100",
			675 => "1111111000101100000001",
			676 => "0000111011000000000100",
			677 => "0000000000101100000001",
			678 => "0000001000101100000001",
			679 => "1111111000101100000001",
			680 => "0010111110011000001100",
			681 => "0001011000000100000100",
			682 => "0000000000101100000001",
			683 => "0000111100010000000100",
			684 => "0000000000101100000001",
			685 => "0000001000101100000001",
			686 => "0011100010110000000100",
			687 => "0000000000101100000001",
			688 => "0011100111001000000100",
			689 => "1111111000101100000001",
			690 => "0011100110110000000100",
			691 => "0000001000101100000001",
			692 => "0000000000101100000001",
			693 => "0011010110001100001000",
			694 => "0010000101011100000100",
			695 => "0000000000101100000001",
			696 => "0000000000101100000001",
			697 => "0010111011101100001000",
			698 => "0001101110101100000100",
			699 => "0000000000101100000001",
			700 => "0000000000101100000001",
			701 => "0011001110011000000100",
			702 => "0000000000101100000001",
			703 => "1111111000101100000001",
			704 => "0011100110110001001000",
			705 => "0000000011001100100100",
			706 => "0001010001111100011100",
			707 => "0001111100000000001100",
			708 => "0000000100110000000100",
			709 => "0000000000101110101101",
			710 => "0010001111111100000100",
			711 => "0000000000101110101101",
			712 => "0000000000101110101101",
			713 => "0000001011111100000100",
			714 => "0000000000101110101101",
			715 => "0011011110011000000100",
			716 => "0000000000101110101101",
			717 => "0011110100001000000100",
			718 => "0000000000101110101101",
			719 => "0000000000101110101101",
			720 => "0001011001101100000100",
			721 => "0000000000101110101101",
			722 => "0000000000101110101101",
			723 => "0000010110010000010000",
			724 => "0000110011100100001000",
			725 => "0000100110111100000100",
			726 => "0000000000101110101101",
			727 => "0000000000101110101101",
			728 => "0010101001010100000100",
			729 => "0000000000101110101101",
			730 => "0000001000101110101101",
			731 => "0000111101001000001000",
			732 => "0000000101101000000100",
			733 => "0000000000101110101101",
			734 => "0000000000101110101101",
			735 => "0001010110011100000100",
			736 => "0000000000101110101101",
			737 => "0001001100010000000100",
			738 => "0000000000101110101101",
			739 => "0000000000101110101101",
			740 => "0000010110010000000100",
			741 => "0000000000101110101101",
			742 => "0010011100101000001000",
			743 => "0011110100110100000100",
			744 => "0000000000101110101101",
			745 => "0000000000101110101101",
			746 => "0000000000101110101101",
			747 => "0000001101110001000100",
			748 => "0010101011111000100100",
			749 => "0010110110001100001000",
			750 => "0011001011101100000100",
			751 => "0000000000110001101001",
			752 => "0000000000110001101001",
			753 => "0001000101011100001100",
			754 => "0001100001100000001000",
			755 => "0011100010000000000100",
			756 => "0000000000110001101001",
			757 => "0000000000110001101001",
			758 => "0000000000110001101001",
			759 => "0001010001010000001000",
			760 => "0001101010111100000100",
			761 => "0000000000110001101001",
			762 => "0000000000110001101001",
			763 => "0001100110111000000100",
			764 => "0000000000110001101001",
			765 => "0000000000110001101001",
			766 => "0010010110000000001000",
			767 => "0001001111101000000100",
			768 => "0000000000110001101001",
			769 => "0000000000110001101001",
			770 => "0011110001101100010100",
			771 => "0001000011000100001100",
			772 => "0000010110010000000100",
			773 => "0000000000110001101001",
			774 => "0000110011000100000100",
			775 => "0000000000110001101001",
			776 => "0000000000110001101001",
			777 => "0001101110111100000100",
			778 => "0000000000110001101001",
			779 => "0000000000110001101001",
			780 => "0000000000110001101001",
			781 => "0010000101011100001100",
			782 => "0011011011101100001000",
			783 => "0001001001000100000100",
			784 => "0000000000110001101001",
			785 => "0000000000110001101001",
			786 => "0000000000110001101001",
			787 => "0010000101101100001000",
			788 => "0010101001010100000100",
			789 => "0000000000110001101001",
			790 => "0000000000110001101001",
			791 => "0010100000111100000100",
			792 => "0000000000110001101001",
			793 => "0000000000110001101001",
			794 => "0011001110011000010100",
			795 => "0001100101001100001100",
			796 => "0010001010100100000100",
			797 => "0000000000110100010101",
			798 => "0011011011101100000100",
			799 => "1111111000110100010101",
			800 => "0000000000110100010101",
			801 => "0000010111110000000100",
			802 => "0000001000110100010101",
			803 => "0000000000110100010101",
			804 => "0011100110110000111000",
			805 => "0000010110010000100000",
			806 => "0011101111110000010000",
			807 => "0001001100001100001000",
			808 => "0011001010100100000100",
			809 => "0000000000110100010101",
			810 => "1111111000110100010101",
			811 => "0000010000011000000100",
			812 => "0000000000110100010101",
			813 => "0000000000110100010101",
			814 => "0000110011100100001000",
			815 => "0011010110001100000100",
			816 => "0000000000110100010101",
			817 => "0000000000110100010101",
			818 => "0000001111101100000100",
			819 => "0000000000110100010101",
			820 => "0000001000110100010101",
			821 => "0001011111101000001000",
			822 => "0011111000001000000100",
			823 => "1111111000110100010101",
			824 => "0000000000110100010101",
			825 => "0011010011010000001100",
			826 => "0001000011000100001000",
			827 => "0000010001100100000100",
			828 => "0000000000110100010101",
			829 => "0000000000110100010101",
			830 => "0000000000110100010101",
			831 => "0000000000110100010101",
			832 => "0011000011010000001000",
			833 => "0001101010110000000100",
			834 => "0000000000110100010101",
			835 => "0000000000110100010101",
			836 => "1111111000110100010101",
			837 => "0000010001100100101000",
			838 => "0001011000000100000100",
			839 => "1111111000110101101001",
			840 => "0010001010100100000100",
			841 => "0000001000110101101001",
			842 => "0001010001111100010100",
			843 => "0001001100101100010000",
			844 => "0010101001011000001000",
			845 => "0010000101101100000100",
			846 => "0000000000110101101001",
			847 => "1111111000110101101001",
			848 => "0000001010101000000100",
			849 => "0000000000110101101001",
			850 => "0000001000110101101001",
			851 => "1111111000110101101001",
			852 => "0001010001011100001000",
			853 => "0011110110100000000100",
			854 => "0000000000110101101001",
			855 => "0000001000110101101001",
			856 => "1111111000110101101001",
			857 => "1111111000110101101001",
			858 => "0011010011010000111100",
			859 => "0010101001011000100100",
			860 => "0010000101101100100000",
			861 => "0000101101110000010100",
			862 => "0000010110010000001100",
			863 => "0000100110100100001000",
			864 => "0011001110011000000100",
			865 => "0000000000110111100101",
			866 => "0000000000110111100101",
			867 => "1111111000110111100101",
			868 => "0001011111101000000100",
			869 => "1111111000110111100101",
			870 => "0000001000110111100101",
			871 => "0001101010110000001000",
			872 => "0000001001101000000100",
			873 => "0000000000110111100101",
			874 => "0000001000110111100101",
			875 => "1111111000110111100101",
			876 => "1111111000110111100101",
			877 => "0000010110010000010000",
			878 => "0011101010011000000100",
			879 => "1111111000110111100101",
			880 => "0000011001100100000100",
			881 => "0000001000110111100101",
			882 => "0000001001110100000100",
			883 => "1111111000110111100101",
			884 => "0000000000110111100101",
			885 => "0001000011000100000100",
			886 => "0000001000110111100101",
			887 => "1111111000110111100101",
			888 => "1111111000110111100101",
			889 => "0011011011101101000000",
			890 => "0000001101110000101100",
			891 => "0010101011111000011000",
			892 => "0010110110001100000100",
			893 => "0000000000111010011001",
			894 => "0011100111001000010000",
			895 => "0001000101010100001000",
			896 => "0001111100010000000100",
			897 => "0000000000111010011001",
			898 => "0000000000111010011001",
			899 => "0001111000111000000100",
			900 => "0000000000111010011001",
			901 => "0000000000111010011001",
			902 => "0000000000111010011001",
			903 => "0010011010000100010000",
			904 => "0001011001101100001100",
			905 => "0001100100000000000100",
			906 => "0000000000111010011001",
			907 => "0011010110001100000100",
			908 => "0000000000111010011001",
			909 => "0000000000111010011001",
			910 => "0000000000111010011001",
			911 => "0000000000111010011001",
			912 => "0001000101011100000100",
			913 => "0000000000111010011001",
			914 => "0010001111111100001100",
			915 => "0000000101101000000100",
			916 => "0000000000111010011001",
			917 => "0000001001101000000100",
			918 => "0000000000111010011001",
			919 => "0000000000111010011001",
			920 => "0000000000111010011001",
			921 => "0010001001001100001000",
			922 => "0001000110011100000100",
			923 => "0000000000111010011001",
			924 => "0000000000111010011001",
			925 => "0010111110011000001000",
			926 => "0000111101001000000100",
			927 => "0000000000111010011001",
			928 => "0000000000111010011001",
			929 => "0010101100110100000100",
			930 => "0000000000111010011001",
			931 => "0000111010011100000100",
			932 => "0000000000111010011001",
			933 => "0000000000111010011001",
			934 => "0010110101010100110000",
			935 => "0011100001000000101100",
			936 => "0010101001011000011000",
			937 => "0010000101101100010100",
			938 => "0000001110110000010000",
			939 => "0010001010100100001000",
			940 => "0000001101001100000100",
			941 => "0000000000111011111101",
			942 => "0000001000111011111101",
			943 => "0011111000001000000100",
			944 => "0000000000111011111101",
			945 => "1111111000111011111101",
			946 => "0000001000111011111101",
			947 => "1111111000111011111101",
			948 => "0001000110011100001100",
			949 => "0000010110010000001000",
			950 => "0000001101110100000100",
			951 => "1111111000111011111101",
			952 => "0000001000111011111101",
			953 => "0000001000111011111101",
			954 => "0001001100001100000100",
			955 => "1111111000111011111101",
			956 => "0000001000111011111101",
			957 => "1111111000111011111101",
			958 => "1111111000111011111101",
			959 => "0010001010100100001000",
			960 => "0010010101010100000100",
			961 => "0000000000111110000001",
			962 => "0000000000111110000001",
			963 => "0001011000000000001000",
			964 => "0000111101001000000100",
			965 => "0000000000111110000001",
			966 => "0000000000111110000001",
			967 => "0000000101101000101000",
			968 => "0001111100110000010100",
			969 => "0000011001100100001000",
			970 => "0010001001001100000100",
			971 => "0000000000111110000001",
			972 => "0000000000111110000001",
			973 => "0000000100110000000100",
			974 => "0000000000111110000001",
			975 => "0010101110111000000100",
			976 => "0000000000111110000001",
			977 => "0000000000111110000001",
			978 => "0000111101001000001000",
			979 => "0011100001101100000100",
			980 => "0000000000111110000001",
			981 => "0000000000111110000001",
			982 => "0010111110011000000100",
			983 => "0000000000111110000001",
			984 => "0010000101011100000100",
			985 => "0000000000111110000001",
			986 => "0000000000111110000001",
			987 => "0011011011101100000100",
			988 => "0000000000111110000001",
			989 => "0001000110000000000100",
			990 => "0000000000111110000001",
			991 => "0000000000111110000001",
			992 => "0001001001000100011100",
			993 => "0000111000000000010000",
			994 => "0000101111001100001100",
			995 => "0000111111011000001000",
			996 => "0000110011000000000100",
			997 => "0000000001000001001101",
			998 => "0000000001000001001101",
			999 => "1111111001000001001101",
			1000 => "0000000001000001001101",
			1001 => "0011101110100000001000",
			1002 => "0001111100010000000100",
			1003 => "0000000001000001001101",
			1004 => "0000000001000001001101",
			1005 => "0000000001000001001101",
			1006 => "0000010111100100101000",
			1007 => "0000000011001100011100",
			1008 => "0011010110001100000100",
			1009 => "0000000001000001001101",
			1010 => "0011011011101100001100",
			1011 => "0010011010000100001000",
			1012 => "0000000100110000000100",
			1013 => "0000000001000001001101",
			1014 => "0000000001000001001101",
			1015 => "0000000001000001001101",
			1016 => "0010001001001100000100",
			1017 => "0000000001000001001101",
			1018 => "0001011001010000000100",
			1019 => "0000000001000001001101",
			1020 => "0000000001000001001101",
			1021 => "0001011100110000000100",
			1022 => "0000000001000001001101",
			1023 => "0010001111111100000100",
			1024 => "0000001001000001001101",
			1025 => "0000000001000001001101",
			1026 => "0000111011111000011000",
			1027 => "0011001110011000000100",
			1028 => "0000000001000001001101",
			1029 => "0011110110011000001100",
			1030 => "0001011000100000000100",
			1031 => "0000000001000001001101",
			1032 => "0001010000111100000100",
			1033 => "0000000001000001001101",
			1034 => "0000000001000001001101",
			1035 => "0001100000010000000100",
			1036 => "0000000001000001001101",
			1037 => "0000000001000001001101",
			1038 => "0011100101001000000100",
			1039 => "0000000001000001001101",
			1040 => "0011010011010000000100",
			1041 => "0000000001000001001101",
			1042 => "0000000001000001001101",
			1043 => "0000110000111100110100",
			1044 => "0010010110000000110000",
			1045 => "0010101011111000100100",
			1046 => "0000011000011000100000",
			1047 => "0011001110011000010000",
			1048 => "0001100101001100001000",
			1049 => "0010001010100100000100",
			1050 => "0000000001000011010001",
			1051 => "1111111001000011010001",
			1052 => "0001101101010000000100",
			1053 => "0000001001000011010001",
			1054 => "0000000001000011010001",
			1055 => "0011100110110000001000",
			1056 => "0011101111110000000100",
			1057 => "1111111001000011010001",
			1058 => "0000000001000011010001",
			1059 => "0001100000001100000100",
			1060 => "1111111001000011010001",
			1061 => "0000000001000011010001",
			1062 => "1111111001000011010001",
			1063 => "0001001001010000001000",
			1064 => "0000010001110000000100",
			1065 => "0000000001000011010001",
			1066 => "0000001001000011010001",
			1067 => "0000000001000011010001",
			1068 => "1111111001000011010001",
			1069 => "0001011001101100001100",
			1070 => "0011111001011100000100",
			1071 => "0000000001000011010001",
			1072 => "0001100101100000000100",
			1073 => "0000001001000011010001",
			1074 => "0000000001000011010001",
			1075 => "0000000001000011010001",
			1076 => "0001110110101100101100",
			1077 => "0000111000000000010000",
			1078 => "0001001001000100000100",
			1079 => "1111111001000110010101",
			1080 => "0000010001110000000100",
			1081 => "0000000001000110010101",
			1082 => "0001000110000000000100",
			1083 => "0000000001000110010101",
			1084 => "0000000001000110010101",
			1085 => "0000011000011000011000",
			1086 => "0001011011000000001000",
			1087 => "0011110001000100000100",
			1088 => "0000000001000110010101",
			1089 => "0000001001000110010101",
			1090 => "0010101001000000001000",
			1091 => "0010001001001100000100",
			1092 => "0000000001000110010101",
			1093 => "0000000001000110010101",
			1094 => "0001011001101100000100",
			1095 => "0000000001000110010101",
			1096 => "0000000001000110010101",
			1097 => "0000000001000110010101",
			1098 => "0000001110110000101100",
			1099 => "0010010101011100001000",
			1100 => "0000010111100100000100",
			1101 => "1111111001000110010101",
			1102 => "0000000001000110010101",
			1103 => "0010001001001100001000",
			1104 => "0000001000010000000100",
			1105 => "0000000001000110010101",
			1106 => "0000000001000110010101",
			1107 => "0010101001010100001100",
			1108 => "0011100011010100001000",
			1109 => "0001100011011000000100",
			1110 => "0000000001000110010101",
			1111 => "0000000001000110010101",
			1112 => "1111111001000110010101",
			1113 => "0010011001000100001000",
			1114 => "0000000011001100000100",
			1115 => "0000000001000110010101",
			1116 => "0000000001000110010101",
			1117 => "0010101100110100000100",
			1118 => "0000000001000110010101",
			1119 => "0000000001000110010101",
			1120 => "0011100001000000001000",
			1121 => "0011000111011100000100",
			1122 => "0000001001000110010101",
			1123 => "0000000001000110010101",
			1124 => "0000000001000110010101",
			1125 => "0001101100100000000100",
			1126 => "0000000001001000100001",
			1127 => "0011101101100100111000",
			1128 => "0000010110010000100100",
			1129 => "0010010101011100010000",
			1130 => "0010001001001100001000",
			1131 => "0010111011101100000100",
			1132 => "0000000001001000100001",
			1133 => "1111111001001000100001",
			1134 => "0001011000000100000100",
			1135 => "0000000001001000100001",
			1136 => "0000000001001000100001",
			1137 => "0001001100010000001000",
			1138 => "0000110011001000000100",
			1139 => "0000000001001000100001",
			1140 => "0000001001001000100001",
			1141 => "0000110000111100000100",
			1142 => "0000000001001000100001",
			1143 => "0010101100110100000100",
			1144 => "0000000001001000100001",
			1145 => "0000000001001000100001",
			1146 => "0000111011111000001100",
			1147 => "0000100111111000001000",
			1148 => "0001011000100000000100",
			1149 => "1111111001001000100001",
			1150 => "0000000001001000100001",
			1151 => "0000000001001000100001",
			1152 => "0011010111011100000100",
			1153 => "0000000001001000100001",
			1154 => "0000000001001000100001",
			1155 => "0010010101011100001000",
			1156 => "0010101001010100000100",
			1157 => "0000000001001000100001",
			1158 => "0000000001001000100001",
			1159 => "0000000001001000100001",
			1160 => "0011100110110001010000",
			1161 => "0011100111001000111000",
			1162 => "0001010110101100010100",
			1163 => "0001001100101000001100",
			1164 => "0001000101010100000100",
			1165 => "0000000001001011011101",
			1166 => "0010101000000000000100",
			1167 => "0000000001001011011101",
			1168 => "0000000001001011011101",
			1169 => "0001001010000100000100",
			1170 => "1111111001001011011101",
			1171 => "0000000001001011011101",
			1172 => "0001001111011000001100",
			1173 => "0010000101101100001000",
			1174 => "0000000011001100000100",
			1175 => "0000000001001011011101",
			1176 => "0000001001001011011101",
			1177 => "0000000001001011011101",
			1178 => "0010101001000000001100",
			1179 => "0010011001001000000100",
			1180 => "0000000001001011011101",
			1181 => "0010001001001100000100",
			1182 => "0000000001001011011101",
			1183 => "0000000001001011011101",
			1184 => "0011010110001100000100",
			1185 => "0000000001001011011101",
			1186 => "0001011001101100000100",
			1187 => "0000000001001011011101",
			1188 => "0000000001001011011101",
			1189 => "0000010110010000000100",
			1190 => "0000001001001011011101",
			1191 => "0000111101001000001000",
			1192 => "0001011100010000000100",
			1193 => "0000000001001011011101",
			1194 => "0000000001001011011101",
			1195 => "0001011011000000000100",
			1196 => "0000000001001011011101",
			1197 => "0010101001011000000100",
			1198 => "0000000001001011011101",
			1199 => "0000000001001011011101",
			1200 => "0000010001110000000100",
			1201 => "0000000001001011011101",
			1202 => "0001011100110000000100",
			1203 => "0000000001001011011101",
			1204 => "0010010101101100000100",
			1205 => "0000000001001011011101",
			1206 => "0000000001001011011101",
			1207 => "0001110110101100110000",
			1208 => "0010101001010100011000",
			1209 => "0011001010100100001100",
			1210 => "0001001001000100000100",
			1211 => "0000000001001111000001",
			1212 => "0000011000011000000100",
			1213 => "0000000001001111000001",
			1214 => "0000000001001111000001",
			1215 => "0001111100010000000100",
			1216 => "0000000001001111000001",
			1217 => "0000111111011000000100",
			1218 => "0000000001001111000001",
			1219 => "0000000001001111000001",
			1220 => "0011101010110100001100",
			1221 => "0010000101101100000100",
			1222 => "0000000001001111000001",
			1223 => "0011100010001100000100",
			1224 => "0000000001001111000001",
			1225 => "0000000001001111000001",
			1226 => "0001011001101100001000",
			1227 => "0000100111000100000100",
			1228 => "0000000001001111000001",
			1229 => "0000000001001111000001",
			1230 => "0000000001001111000001",
			1231 => "0000001110110000111000",
			1232 => "0000100000101000101100",
			1233 => "0000000000000000100000",
			1234 => "0011111010110000010000",
			1235 => "0011111110001000001000",
			1236 => "0000011001100000000100",
			1237 => "0000000001001111000001",
			1238 => "0000000001001111000001",
			1239 => "0010011001000100000100",
			1240 => "0000000001001111000001",
			1241 => "0000000001001111000001",
			1242 => "0000111000101000001000",
			1243 => "0001010001010000000100",
			1244 => "0000000001001111000001",
			1245 => "0000000001001111000001",
			1246 => "0000111111101000000100",
			1247 => "0000000001001111000001",
			1248 => "0000000001001111000001",
			1249 => "0000010110010000000100",
			1250 => "0000000001001111000001",
			1251 => "0000111100101100000100",
			1252 => "0000000001001111000001",
			1253 => "0000000001001111000001",
			1254 => "0001011111101000000100",
			1255 => "0000000001001111000001",
			1256 => "0001010000111100000100",
			1257 => "0000000001001111000001",
			1258 => "0000000001001111000001",
			1259 => "0011100001000000001000",
			1260 => "0010000101101100000100",
			1261 => "0000000001001111000001",
			1262 => "0000000001001111000001",
			1263 => "0000000001001111000001",
			1264 => "0001011000000000001000",
			1265 => "0000111101001000000100",
			1266 => "0000000001010001010101",
			1267 => "0000000001010001010101",
			1268 => "0010000011010000001000",
			1269 => "0010010101011100000100",
			1270 => "0000000001010001010101",
			1271 => "0000000001010001010101",
			1272 => "0000010111100100100000",
			1273 => "0001111101001000010000",
			1274 => "0000110011100100000100",
			1275 => "0000000001010001010101",
			1276 => "0011110000000100001000",
			1277 => "0011010110001100000100",
			1278 => "0000000001010001010101",
			1279 => "0000000001010001010101",
			1280 => "0000001001010001010101",
			1281 => "0000000101101000001100",
			1282 => "0010000101011100000100",
			1283 => "0000000001010001010101",
			1284 => "0000111111101000000100",
			1285 => "1111111001010001010101",
			1286 => "0000000001010001010101",
			1287 => "0000000001010001010101",
			1288 => "0000111011111000010000",
			1289 => "0011001110011000000100",
			1290 => "0000000001010001010101",
			1291 => "0001011000100000000100",
			1292 => "0000000001010001010101",
			1293 => "0001010001001000000100",
			1294 => "0000000001010001010101",
			1295 => "0000000001010001010101",
			1296 => "0011100101001000000100",
			1297 => "0000000001010001010101",
			1298 => "0011010011010000000100",
			1299 => "0000000001010001010101",
			1300 => "0000000001010001010101",
			1301 => "0011100110110001010100",
			1302 => "0011011011101100110000",
			1303 => "0011101101100000101000",
			1304 => "0010010101011100010100",
			1305 => "0010110110001100001000",
			1306 => "0010110110110100000100",
			1307 => "0000000001010100100001",
			1308 => "0000000001010100100001",
			1309 => "0010001010100100000100",
			1310 => "0000000001010100100001",
			1311 => "0010001001001100000100",
			1312 => "0000000001010100100001",
			1313 => "0000000001010100100001",
			1314 => "0010101100010000001000",
			1315 => "0010011100101000000100",
			1316 => "0000000001010100100001",
			1317 => "0000000001010100100001",
			1318 => "0010011010000100001000",
			1319 => "0000000100110000000100",
			1320 => "0000000001010100100001",
			1321 => "0000000001010100100001",
			1322 => "0000000001010100100001",
			1323 => "0000010110010000000100",
			1324 => "0000000001010100100001",
			1325 => "0000000001010100100001",
			1326 => "0010001001001100001000",
			1327 => "0001100101001000000100",
			1328 => "0000000001010100100001",
			1329 => "0000000001010100100001",
			1330 => "0000111101001000000100",
			1331 => "0000000001010100100001",
			1332 => "0000001011111100001100",
			1333 => "0010101100110100000100",
			1334 => "0000000001010100100001",
			1335 => "0001011001101100000100",
			1336 => "0000000001010100100001",
			1337 => "0000000001010100100001",
			1338 => "0011110010111100001000",
			1339 => "0000111100101100000100",
			1340 => "0000000001010100100001",
			1341 => "0000000001010100100001",
			1342 => "0000000001010100100001",
			1343 => "0010111011101100001000",
			1344 => "0011110011111100000100",
			1345 => "0000000001010100100001",
			1346 => "0000000001010100100001",
			1347 => "0000010110010000000100",
			1348 => "0000000001010100100001",
			1349 => "0000011000011000000100",
			1350 => "0000000001010100100001",
			1351 => "0000000001010100100001",
			1352 => "0000011001100100011100",
			1353 => "0010001111111100010100",
			1354 => "0010010101011100001000",
			1355 => "0011001110011000000100",
			1356 => "1111111001011000000101",
			1357 => "0000000001011000000101",
			1358 => "0010011001001000000100",
			1359 => "0000000001011000000101",
			1360 => "0001000101101100000100",
			1361 => "0000000001011000000101",
			1362 => "1111111001011000000101",
			1363 => "0010011010000100000100",
			1364 => "0000001001011000000101",
			1365 => "0000000001011000000101",
			1366 => "0010000101011100101000",
			1367 => "0000011000011000100100",
			1368 => "0001001001000100010000",
			1369 => "0001001100101000001100",
			1370 => "0001000101010100001000",
			1371 => "0011011011101100000100",
			1372 => "0000000001011000000101",
			1373 => "0000000001011000000101",
			1374 => "0000001001011000000101",
			1375 => "0000000001011000000101",
			1376 => "0001000110011100010000",
			1377 => "0000101011100100001000",
			1378 => "0000001001110100000100",
			1379 => "0000000001011000000101",
			1380 => "0000001001011000000101",
			1381 => "0011101100011000000100",
			1382 => "0000001001011000000101",
			1383 => "0000000001011000000101",
			1384 => "0000000001011000000101",
			1385 => "1111111001011000000101",
			1386 => "0000111101001000010000",
			1387 => "0000001001101000001000",
			1388 => "0010100100101100000100",
			1389 => "1111111001011000000101",
			1390 => "0000000001011000000101",
			1391 => "0000001101011000000100",
			1392 => "0000001001011000000101",
			1393 => "0000000001011000000101",
			1394 => "0010010101101100001000",
			1395 => "0010000101101100000100",
			1396 => "0000001001011000000101",
			1397 => "0000000001011000000101",
			1398 => "0000111011111000001000",
			1399 => "0010110011010000000100",
			1400 => "0000000001011000000101",
			1401 => "1111111001011000000101",
			1402 => "0011100101001000001000",
			1403 => "0011100010001100000100",
			1404 => "0000000001011000000101",
			1405 => "1111111001011000000101",
			1406 => "0011010011010000000100",
			1407 => "0000001001011000000101",
			1408 => "1111111001011000000101",
			1409 => "0001101100100000000100",
			1410 => "0000000001011010010001",
			1411 => "0011101101100100111000",
			1412 => "0000001110110000110000",
			1413 => "0011101111110100010100",
			1414 => "0000101111101100010000",
			1415 => "0001101111110000001000",
			1416 => "0011001001001000000100",
			1417 => "0000000001011010010001",
			1418 => "0000000001011010010001",
			1419 => "0001000101011100000100",
			1420 => "0000000001011010010001",
			1421 => "0000000001011010010001",
			1422 => "0000001001011010010001",
			1423 => "0001001010000100010000",
			1424 => "0000100110101000001000",
			1425 => "0010101101001000000100",
			1426 => "0000000001011010010001",
			1427 => "0000000001011010010001",
			1428 => "0011100111001000000100",
			1429 => "1111111001011010010001",
			1430 => "0000000001011010010001",
			1431 => "0000001111001100001000",
			1432 => "0000010001100100000100",
			1433 => "0000000001011010010001",
			1434 => "0000000001011010010001",
			1435 => "0000000001011010010001",
			1436 => "0010000101101100000100",
			1437 => "0000001001011010010001",
			1438 => "0000000001011010010001",
			1439 => "0010010101011100001000",
			1440 => "0010101001010100000100",
			1441 => "0000000001011010010001",
			1442 => "0000000001011010010001",
			1443 => "0000000001011010010001",
			1444 => "0000010001100101011000",
			1445 => "0000011000111100001000",
			1446 => "0011010110110100000100",
			1447 => "1111111001011101000111",
			1448 => "0000000001011101000111",
			1449 => "0000001101110000110000",
			1450 => "0010101011111000011100",
			1451 => "0011100010110000010000",
			1452 => "0001000101010100001000",
			1453 => "0000111000000000000100",
			1454 => "1111111001011101000111",
			1455 => "0000001001011101000111",
			1456 => "0011011110011000000100",
			1457 => "1111111001011101000111",
			1458 => "0000000001011101000111",
			1459 => "0011001110011000000100",
			1460 => "1111111001011101000111",
			1461 => "0000010111100100000100",
			1462 => "0000001001011101000111",
			1463 => "1111111001011101000111",
			1464 => "0001011001101100010000",
			1465 => "0000010001110000001000",
			1466 => "0000011000111100000100",
			1467 => "0000001001011101000111",
			1468 => "0000000001011101000111",
			1469 => "0001000011000100000100",
			1470 => "0000001001011101000111",
			1471 => "1111111001011101000111",
			1472 => "1111111001011101000111",
			1473 => "0001111101001000001100",
			1474 => "0011111101001100000100",
			1475 => "0000001001011101000111",
			1476 => "0011110101000100000100",
			1477 => "0000000001011101000111",
			1478 => "0000001001011101000111",
			1479 => "0000000101101000001000",
			1480 => "0000001011001100000100",
			1481 => "0000000001011101000111",
			1482 => "1111111001011101000111",
			1483 => "0011100001000000001000",
			1484 => "0011011011101100000100",
			1485 => "0000001001011101000111",
			1486 => "0000000001011101000111",
			1487 => "1111111001011101000111",
			1488 => "1111111001011101000111",
			1489 => "0010011001000100100000",
			1490 => "0000001101110100001000",
			1491 => "0000111111101000000100",
			1492 => "1111111001011110101001",
			1493 => "0000000001011110101001",
			1494 => "0000011000011000010100",
			1495 => "0001011000000100000100",
			1496 => "1111111001011110101001",
			1497 => "0011100110110000001100",
			1498 => "0000110011100100000100",
			1499 => "0000001001011110101001",
			1500 => "0011001110011000000100",
			1501 => "0000001001011110101001",
			1502 => "0000010001011110101001",
			1503 => "0000000001011110101001",
			1504 => "1111111001011110101001",
			1505 => "0011001100101000010000",
			1506 => "0010101001000000000100",
			1507 => "1111111001011110101001",
			1508 => "0000010110010000001000",
			1509 => "0001001100001100000100",
			1510 => "1111111001011110101001",
			1511 => "0000000001011110101001",
			1512 => "0000001001011110101001",
			1513 => "1111111001011110101001",
			1514 => "0000000011001100100000",
			1515 => "0010101001000000010100",
			1516 => "0010001010100100000100",
			1517 => "0000000001100000111101",
			1518 => "0011001010100100001100",
			1519 => "0001111100000000000100",
			1520 => "0000000001100000111101",
			1521 => "0011001110011000000100",
			1522 => "0000000001100000111101",
			1523 => "0000000001100000111101",
			1524 => "0000000001100000111101",
			1525 => "0000010110010000000100",
			1526 => "0000000001100000111101",
			1527 => "0010010011000000000100",
			1528 => "0000000001100000111101",
			1529 => "0000000001100000111101",
			1530 => "0011100110110000011000",
			1531 => "0000010110010000001100",
			1532 => "0011001110011000000100",
			1533 => "0000000001100000111101",
			1534 => "0001011000000000000100",
			1535 => "0000000001100000111101",
			1536 => "0000000001100000111101",
			1537 => "0011110010111100000100",
			1538 => "0000000001100000111101",
			1539 => "0000000101010000000100",
			1540 => "0000000001100000111101",
			1541 => "0000000001100000111101",
			1542 => "0010111011101100001000",
			1543 => "0011110011100000000100",
			1544 => "0000000001100000111101",
			1545 => "0000000001100000111101",
			1546 => "0000010110010000000100",
			1547 => "0000000001100000111101",
			1548 => "0000011000011000000100",
			1549 => "0000000001100000111101",
			1550 => "0000000001100000111101",
			1551 => "0001011000000000001000",
			1552 => "0000111101001000000100",
			1553 => "1111111001100010010001",
			1554 => "0000000001100010010001",
			1555 => "0000001110110000011100",
			1556 => "0011111101001100011000",
			1557 => "0011010011010000010100",
			1558 => "0000001111001100010000",
			1559 => "0010101001010100001000",
			1560 => "0010001001001100000100",
			1561 => "0000000001100010010001",
			1562 => "1111111001100010010001",
			1563 => "0000011001100100000100",
			1564 => "0000000001100010010001",
			1565 => "0000000001100010010001",
			1566 => "0000001001100010010001",
			1567 => "1111111001100010010001",
			1568 => "1111111001100010010001",
			1569 => "0001111000101000000100",
			1570 => "0000001001100010010001",
			1571 => "1111111001100010010001",
			1572 => "0010011001000100100100",
			1573 => "0000001101110100001000",
			1574 => "0000111111101000000100",
			1575 => "1111111001100011111101",
			1576 => "0000000001100011111101",
			1577 => "0000011000011000011000",
			1578 => "0001011000000100000100",
			1579 => "1111111001100011111101",
			1580 => "0011100110110000010000",
			1581 => "0010101001010100001000",
			1582 => "0011010110001100000100",
			1583 => "0000001001100011111101",
			1584 => "0000000001100011111101",
			1585 => "0011010110001100000100",
			1586 => "0000001001100011111101",
			1587 => "0000010001100011111101",
			1588 => "0000000001100011111101",
			1589 => "1111111001100011111101",
			1590 => "0011001100101000010000",
			1591 => "0010101001000000000100",
			1592 => "1111111001100011111101",
			1593 => "0001011001101100001000",
			1594 => "0010001111111100000100",
			1595 => "0000000001100011111101",
			1596 => "0000010001100011111101",
			1597 => "1111111001100011111101",
			1598 => "1111111001100011111101",
			1599 => "0010011001000100101000",
			1600 => "0000001011111100001000",
			1601 => "0000111111101000000100",
			1602 => "1111111001100101110001",
			1603 => "0000000001100101110001",
			1604 => "0011100110110000011000",
			1605 => "0000110101111000000100",
			1606 => "1111111001100101110001",
			1607 => "0000011000011000010000",
			1608 => "0010101001010100001000",
			1609 => "0011010110001100000100",
			1610 => "0000001001100101110001",
			1611 => "0000000001100101110001",
			1612 => "0011111101001100000100",
			1613 => "0000001001100101110001",
			1614 => "0000001001100101110001",
			1615 => "0000000001100101110001",
			1616 => "0001111001010000000100",
			1617 => "0000000001100101110001",
			1618 => "1111111001100101110001",
			1619 => "0011001100101000010000",
			1620 => "0010101001000000000100",
			1621 => "1111111001100101110001",
			1622 => "0011101010011000001000",
			1623 => "0000000100001000000100",
			1624 => "0000001001100101110001",
			1625 => "1111111001100101110001",
			1626 => "0000010001100101110001",
			1627 => "1111111001100101110001",
			1628 => "0011001100101000101000",
			1629 => "0001100101001000001100",
			1630 => "0010000101101100000100",
			1631 => "1111111001100111000101",
			1632 => "0001010010111000000100",
			1633 => "1111111001100111000101",
			1634 => "0000001001100111000101",
			1635 => "0011100001000000011000",
			1636 => "0001011000000100000100",
			1637 => "1111111001100111000101",
			1638 => "0000010001100100010000",
			1639 => "0001010001111100001000",
			1640 => "0010010110000000000100",
			1641 => "0000000001100111000101",
			1642 => "1111111001100111000101",
			1643 => "0001010111010100000100",
			1644 => "0000010001100111000101",
			1645 => "1111111001100111000101",
			1646 => "1111111001100111000101",
			1647 => "1111111001100111000101",
			1648 => "1111111001100111000101",
			1649 => "0001001001000100011100",
			1650 => "0000111000000000001100",
			1651 => "0010101000111000001000",
			1652 => "0010101000000000000100",
			1653 => "0000000001101001011001",
			1654 => "0000000001101001011001",
			1655 => "0000000001101001011001",
			1656 => "0010011100101000001000",
			1657 => "0001101101010100000100",
			1658 => "0000000001101001011001",
			1659 => "0000000001101001011001",
			1660 => "0001100100000100000100",
			1661 => "0000000001101001011001",
			1662 => "0000000001101001011001",
			1663 => "0010000101101100100000",
			1664 => "0011011010100100011100",
			1665 => "0010101100010000001000",
			1666 => "0001001010000100000100",
			1667 => "0000000001101001011001",
			1668 => "0000000001101001011001",
			1669 => "0000011000011000010000",
			1670 => "0011101001011100001000",
			1671 => "0001010001111100000100",
			1672 => "0000000001101001011001",
			1673 => "0000000001101001011001",
			1674 => "0011100110110000000100",
			1675 => "0000000001101001011001",
			1676 => "0000000001101001011001",
			1677 => "0000000001101001011001",
			1678 => "0000000001101001011001",
			1679 => "0010101001011000000100",
			1680 => "0000000001101001011001",
			1681 => "0011001100101000001000",
			1682 => "0011100101001000000100",
			1683 => "0000000001101001011001",
			1684 => "0000000001101001011001",
			1685 => "0000000001101001011001",
			1686 => "0001011101001000101000",
			1687 => "0000001001101000100000",
			1688 => "0011010110110100010000",
			1689 => "0000010001110000001100",
			1690 => "0010010101011100001000",
			1691 => "0011010011110000000100",
			1692 => "0000000001101011110101",
			1693 => "0000000001101011110101",
			1694 => "0000000001101011110101",
			1695 => "0000000001101011110101",
			1696 => "0010000011010000000100",
			1697 => "0000000001101011110101",
			1698 => "0001111100110000001000",
			1699 => "0000111000000000000100",
			1700 => "0000000001101011110101",
			1701 => "0000000001101011110101",
			1702 => "0000000001101011110101",
			1703 => "0011110100110100000100",
			1704 => "0000000001101011110101",
			1705 => "0000000001101011110101",
			1706 => "0010000101101100011000",
			1707 => "0011111001011100000100",
			1708 => "0000000001101011110101",
			1709 => "0011011010100100010000",
			1710 => "0000011001100100001000",
			1711 => "0001110110101100000100",
			1712 => "0000000001101011110101",
			1713 => "0000000001101011110101",
			1714 => "0001001001011000000100",
			1715 => "0000000001101011110101",
			1716 => "0000000001101011110101",
			1717 => "0000000001101011110101",
			1718 => "0010101001011000000100",
			1719 => "0000000001101011110101",
			1720 => "0010001111001000001000",
			1721 => "0001001000100000000100",
			1722 => "0000000001101011110101",
			1723 => "0000000001101011110101",
			1724 => "0000000001101011110101",
			1725 => "0010000101101100101100",
			1726 => "0000101101110000100100",
			1727 => "0000100000101000100000",
			1728 => "0000001101110000011000",
			1729 => "0010111010100100001100",
			1730 => "0011010011110000000100",
			1731 => "0000000001101101111001",
			1732 => "0010101011111000000100",
			1733 => "0000000001101101111001",
			1734 => "0000000001101101111001",
			1735 => "0000001011111100001000",
			1736 => "0000110000111100000100",
			1737 => "0000000001101101111001",
			1738 => "0000000001101101111001",
			1739 => "0000000001101101111001",
			1740 => "0001001101101000000100",
			1741 => "0000000001101101111001",
			1742 => "0000000001101101111001",
			1743 => "0000000001101101111001",
			1744 => "0001011000000000000100",
			1745 => "0000000001101101111001",
			1746 => "0000000001101101111001",
			1747 => "0000111011111000001000",
			1748 => "0001011110111000000100",
			1749 => "0000000001101101111001",
			1750 => "0000000001101101111001",
			1751 => "0011001100101000001100",
			1752 => "0010101001011000000100",
			1753 => "0000000001101101111001",
			1754 => "0000010110010000000100",
			1755 => "0000000001101101111001",
			1756 => "0000000001101101111001",
			1757 => "0000000001101101111001",
			1758 => "0000011000011000111100",
			1759 => "0001110110101100011100",
			1760 => "0000001101011100010100",
			1761 => "0010101011111000001000",
			1762 => "0010001010100100000100",
			1763 => "0000000001110000000101",
			1764 => "1111111001110000000101",
			1765 => "0000010110010000001000",
			1766 => "0001101110111100000100",
			1767 => "1111111001110000000101",
			1768 => "0000000001110000000101",
			1769 => "0000001001110000000101",
			1770 => "0011110110011000000100",
			1771 => "0000001001110000000101",
			1772 => "0000000001110000000101",
			1773 => "0000001110110000011000",
			1774 => "0000100110100100010100",
			1775 => "0000001011100100001100",
			1776 => "0011001110011000000100",
			1777 => "1111111001110000000101",
			1778 => "0010010101101100000100",
			1779 => "0000000001110000000101",
			1780 => "1111111001110000000101",
			1781 => "0000010110010000000100",
			1782 => "0000000001110000000101",
			1783 => "1111111001110000000101",
			1784 => "1111111001110000000101",
			1785 => "0011101101100100000100",
			1786 => "0000001001110000000101",
			1787 => "0000000001110000000101",
			1788 => "0001111111101000000100",
			1789 => "1111111001110000000101",
			1790 => "0001110100101100000100",
			1791 => "0000001001110000000101",
			1792 => "1111111001110000000101",
			1793 => "0010101001000000111100",
			1794 => "0000000110101000010100",
			1795 => "0011001010100100001100",
			1796 => "0010000101011100000100",
			1797 => "0000000001110010100001",
			1798 => "0010101001010100000100",
			1799 => "0000000001110010100001",
			1800 => "0000000001110010100001",
			1801 => "0010001001001100000100",
			1802 => "0000000001110010100001",
			1803 => "1111111001110010100001",
			1804 => "0011101111110100001000",
			1805 => "0000000110111100000100",
			1806 => "0000000001110010100001",
			1807 => "0000001001110010100001",
			1808 => "0000001110110000010100",
			1809 => "0010101001010100001000",
			1810 => "0001111001010000000100",
			1811 => "1111111001110010100001",
			1812 => "0000000001110010100001",
			1813 => "0011111101001100001000",
			1814 => "0011111100111100000100",
			1815 => "0000000001110010100001",
			1816 => "0000001001110010100001",
			1817 => "1111111001110010100001",
			1818 => "0011100001000000001000",
			1819 => "0010000101101100000100",
			1820 => "0000001001110010100001",
			1821 => "0000000001110010100001",
			1822 => "0000000001110010100001",
			1823 => "0010010011000000010000",
			1824 => "0010001111111100001000",
			1825 => "0010001001001100000100",
			1826 => "0000000001110010100001",
			1827 => "0000000001110010100001",
			1828 => "0001011001101100000100",
			1829 => "0000001001110010100001",
			1830 => "0000000001110010100001",
			1831 => "0000000001110010100001",
			1832 => "0011100110110001000000",
			1833 => "0000001101110100011100",
			1834 => "0001111100000000001100",
			1835 => "0000000100110000000100",
			1836 => "0000000001110101000101",
			1837 => "0010001111111100000100",
			1838 => "0000000001110101000101",
			1839 => "0000000001110101000101",
			1840 => "0001010001111100000100",
			1841 => "0000000001110101000101",
			1842 => "0000010110010000000100",
			1843 => "0000000001110101000101",
			1844 => "0001010001011100000100",
			1845 => "0000000001110101000101",
			1846 => "0000000001110101000101",
			1847 => "0011001110011000001000",
			1848 => "0001100101001100000100",
			1849 => "0000000001110101000101",
			1850 => "0000000001110101000101",
			1851 => "0000011000011000010000",
			1852 => "0010000101101100001100",
			1853 => "0000110011100100001000",
			1854 => "0011010110001100000100",
			1855 => "0000000001110101000101",
			1856 => "0000000001110101000101",
			1857 => "0000000001110101000101",
			1858 => "0000000001110101000101",
			1859 => "0001111111101000000100",
			1860 => "0000000001110101000101",
			1861 => "0001011100101100000100",
			1862 => "0000000001110101000101",
			1863 => "0000000001110101000101",
			1864 => "0010111011101100001000",
			1865 => "0000011001100000000100",
			1866 => "0000000001110101000101",
			1867 => "0000000001110101000101",
			1868 => "0000010110010000000100",
			1869 => "0000000001110101000101",
			1870 => "0000011000011000000100",
			1871 => "0000000001110101000101",
			1872 => "0000000001110101000101",
			1873 => "0000010111100100110100",
			1874 => "0000011000111100001000",
			1875 => "0011010110110100000100",
			1876 => "1111111001110111011001",
			1877 => "0000000001110111011001",
			1878 => "0001100101000000010100",
			1879 => "0010101111101000000100",
			1880 => "1111111001110111011001",
			1881 => "0000010110010000001100",
			1882 => "0011101100100000001000",
			1883 => "0011000011010000000100",
			1884 => "0000000001110111011001",
			1885 => "1111111001110111011001",
			1886 => "0000001001110111011001",
			1887 => "0000001001110111011001",
			1888 => "0001111100110000000100",
			1889 => "0000001001110111011001",
			1890 => "0010111110011000001000",
			1891 => "0000111100010000000100",
			1892 => "0000000001110111011001",
			1893 => "0000001001110111011001",
			1894 => "0001001001000100000100",
			1895 => "1111111001110111011001",
			1896 => "0000001011001100000100",
			1897 => "0000000001110111011001",
			1898 => "0000000001110111011001",
			1899 => "0011010110001100001000",
			1900 => "0010000101011100000100",
			1901 => "0000000001110111011001",
			1902 => "0000000001110111011001",
			1903 => "0010111011101100001000",
			1904 => "0001101110101100000100",
			1905 => "0000000001110111011001",
			1906 => "0000000001110111011001",
			1907 => "0011001110011000000100",
			1908 => "0000000001110111011001",
			1909 => "1111111001110111011001",
			1910 => "0011100110110001000100",
			1911 => "0000000011001100101000",
			1912 => "0010101001000000010000",
			1913 => "0011001010100100001100",
			1914 => "0010001001001100000100",
			1915 => "0000000001111001111101",
			1916 => "0001111000000100000100",
			1917 => "0000000001111001111101",
			1918 => "0000000001111001111101",
			1919 => "0000000001111001111101",
			1920 => "0000010110010000001100",
			1921 => "0001001100001100000100",
			1922 => "0000000001111001111101",
			1923 => "0010001111111100000100",
			1924 => "0000000001111001111101",
			1925 => "0000000001111001111101",
			1926 => "0001000011000100001000",
			1927 => "0000010011110000000100",
			1928 => "0000000001111001111101",
			1929 => "0000000001111001111101",
			1930 => "0000000001111001111101",
			1931 => "0001010110101100010000",
			1932 => "0011011101000000000100",
			1933 => "0000000001111001111101",
			1934 => "0001100000010000001000",
			1935 => "0001110110101100000100",
			1936 => "0000000001111001111101",
			1937 => "0000000001111001111101",
			1938 => "0000000001111001111101",
			1939 => "0010000101101100000100",
			1940 => "0000001001111001111101",
			1941 => "0000111111101000000100",
			1942 => "0000000001111001111101",
			1943 => "0000000001111001111101",
			1944 => "0000010110010000000100",
			1945 => "0000000001111001111101",
			1946 => "0010011100101000001000",
			1947 => "0011110100110100000100",
			1948 => "0000000001111001111101",
			1949 => "0000000001111001111101",
			1950 => "0000000001111001111101",
			1951 => "0011001110011000011100",
			1952 => "0001100101001100010000",
			1953 => "0010001010100100000100",
			1954 => "0000000001111100101001",
			1955 => "0011011011101100001000",
			1956 => "0001111000111000000100",
			1957 => "0000000001111100101001",
			1958 => "1111111001111100101001",
			1959 => "0000000001111100101001",
			1960 => "0010010101011100001000",
			1961 => "0010001111111100000100",
			1962 => "0000001001111100101001",
			1963 => "0000000001111100101001",
			1964 => "0000000001111100101001",
			1965 => "0011100110110000110000",
			1966 => "0000010110010000011000",
			1967 => "0011101111110000001100",
			1968 => "0001001100001100000100",
			1969 => "1111111001111100101001",
			1970 => "0010001111111100000100",
			1971 => "0000000001111100101001",
			1972 => "0000000001111100101001",
			1973 => "0011111000001000001000",
			1974 => "0001011000000000000100",
			1975 => "0000000001111100101001",
			1976 => "0000001001111100101001",
			1977 => "0000000001111100101001",
			1978 => "0001011111101000001000",
			1979 => "0011111000001000000100",
			1980 => "1111111001111100101001",
			1981 => "0000000001111100101001",
			1982 => "0011010011010000001100",
			1983 => "0001000011000100001000",
			1984 => "0000000100110000000100",
			1985 => "0000000001111100101001",
			1986 => "0000001001111100101001",
			1987 => "0000000001111100101001",
			1988 => "0000000001111100101001",
			1989 => "0000010110010000000100",
			1990 => "1111111001111100101001",
			1991 => "0010011001001000000100",
			1992 => "0000000001111100101001",
			1993 => "0000000001111100101001",
			1994 => "0011111001011100000100",
			1995 => "1111111001111110011101",
			1996 => "0011100110110000101000",
			1997 => "0011001110011000001100",
			1998 => "0011010110001100001000",
			1999 => "0011110100011000000100",
			2000 => "1111111001111110011101",
			2001 => "0000000001111110011101",
			2002 => "0000001001111110011101",
			2003 => "0010001001001100001100",
			2004 => "0010111110011000000100",
			2005 => "0000000001111110011101",
			2006 => "0000111001000000000100",
			2007 => "0000001001111110011101",
			2008 => "0000000001111110011101",
			2009 => "0001111100010000000100",
			2010 => "1111111001111110011101",
			2011 => "0000011000111100000100",
			2012 => "0000001001111110011101",
			2013 => "0000111101001000000100",
			2014 => "0000000001111110011101",
			2015 => "0000000001111110011101",
			2016 => "0010111110011000001100",
			2017 => "0010010101011100000100",
			2018 => "1111111001111110011101",
			2019 => "0011111000100100000100",
			2020 => "0000000001111110011101",
			2021 => "0000000001111110011101",
			2022 => "1111111001111110011101",
			2023 => "0010101001000000111000",
			2024 => "0000000110101000010000",
			2025 => "0011001010100100001100",
			2026 => "0010000101011100000100",
			2027 => "0000000010000000110001",
			2028 => "0010101001010100000100",
			2029 => "0000000010000000110001",
			2030 => "0000000010000000110001",
			2031 => "1111111010000000110001",
			2032 => "0011101111110100001000",
			2033 => "0000000110111100000100",
			2034 => "0000000010000000110001",
			2035 => "0000001010000000110001",
			2036 => "0000001110110000010100",
			2037 => "0001110110101100000100",
			2038 => "0000000010000000110001",
			2039 => "0001100000001100001000",
			2040 => "0000111000101000000100",
			2041 => "1111111010000000110001",
			2042 => "0000000010000000110001",
			2043 => "0001001010000100000100",
			2044 => "0000000010000000110001",
			2045 => "0000000010000000110001",
			2046 => "0011100001000000001000",
			2047 => "0010000101101100000100",
			2048 => "0000001010000000110001",
			2049 => "0000000010000000110001",
			2050 => "0000000010000000110001",
			2051 => "0010010011000000010000",
			2052 => "0011010110001100000100",
			2053 => "0000000010000000110001",
			2054 => "0001011001101100001000",
			2055 => "0011111001011100000100",
			2056 => "0000000010000000110001",
			2057 => "0000001010000000110001",
			2058 => "0000000010000000110001",
			2059 => "0000000010000000110001",
			2060 => "0011011011101100111000",
			2061 => "0001001001000100010000",
			2062 => "0000111000000000001100",
			2063 => "0000111111011000001000",
			2064 => "0000110011000000000100",
			2065 => "0000000010000011001101",
			2066 => "0000000010000011001101",
			2067 => "0000000010000011001101",
			2068 => "0000000010000011001101",
			2069 => "0011111011110100100000",
			2070 => "0001110110101100010100",
			2071 => "0000010111100100010000",
			2072 => "0011000011010000001000",
			2073 => "0001111000000100000100",
			2074 => "0000000010000011001101",
			2075 => "0000000010000011001101",
			2076 => "0000111011000000000100",
			2077 => "0000000010000011001101",
			2078 => "0000000010000011001101",
			2079 => "0000000010000011001101",
			2080 => "0001000101111000000100",
			2081 => "0000000010000011001101",
			2082 => "0000000010101100000100",
			2083 => "0000000010000011001101",
			2084 => "0000000010000011001101",
			2085 => "0000010001110000000100",
			2086 => "0000000010000011001101",
			2087 => "0000000010000011001101",
			2088 => "0010001001001100000100",
			2089 => "0000000010000011001101",
			2090 => "0010111110011000001000",
			2091 => "0000111101001000000100",
			2092 => "0000000010000011001101",
			2093 => "0000000010000011001101",
			2094 => "0010101100110100000100",
			2095 => "0000000010000011001101",
			2096 => "0000110011110100000100",
			2097 => "0000000010000011001101",
			2098 => "0000000010000011001101",
			2099 => "0011010011010000100100",
			2100 => "0001011000000100000100",
			2101 => "1111111010000100011001",
			2102 => "0011100001000000011100",
			2103 => "0000000100110000000100",
			2104 => "1111111010000100011001",
			2105 => "0011001110011000001000",
			2106 => "0001100101001100000100",
			2107 => "1111111010000100011001",
			2108 => "0000001010000100011001",
			2109 => "0010001001001100001000",
			2110 => "0010010101011100000100",
			2111 => "0000000010000100011001",
			2112 => "0000001010000100011001",
			2113 => "0011011011101100000100",
			2114 => "0000000010000100011001",
			2115 => "0000000010000100011001",
			2116 => "1111111010000100011001",
			2117 => "1111111010000100011001",
			2118 => "0010101101001000011000",
			2119 => "0010001010100100000100",
			2120 => "0000000010000110111101",
			2121 => "0001011100110000001100",
			2122 => "0011011110011000000100",
			2123 => "1111111010000110111101",
			2124 => "0011110111000000000100",
			2125 => "0000000010000110111101",
			2126 => "0000000010000110111101",
			2127 => "0001000110000000000100",
			2128 => "0000000010000110111101",
			2129 => "0000000010000110111101",
			2130 => "0011011010100100100100",
			2131 => "0000011000011000100000",
			2132 => "0000011001100100001100",
			2133 => "0011010110001100001000",
			2134 => "0010101001011000000100",
			2135 => "0000000010000110111101",
			2136 => "0000000010000110111101",
			2137 => "0000000010000110111101",
			2138 => "0001000110011100010000",
			2139 => "0011101101100100001000",
			2140 => "0000001101110100000100",
			2141 => "0000000010000110111101",
			2142 => "0000001010000110111101",
			2143 => "0011001010100100000100",
			2144 => "0000000010000110111101",
			2145 => "0000000010000110111101",
			2146 => "0000000010000110111101",
			2147 => "0000000010000110111101",
			2148 => "0010101100110100010000",
			2149 => "0011101111010100001000",
			2150 => "0011000111011100000100",
			2151 => "0000000010000110111101",
			2152 => "0000000010000110111101",
			2153 => "0011100110110000000100",
			2154 => "0000000010000110111101",
			2155 => "0000000010000110111101",
			2156 => "0000111010011100000100",
			2157 => "0000000010000110111101",
			2158 => "0000000010000110111101",
			2159 => "0001110110101100101000",
			2160 => "0000100010100100100000",
			2161 => "0010101001000000010100",
			2162 => "0010001010100100000100",
			2163 => "0000000010001001101001",
			2164 => "0001111100000000001000",
			2165 => "0001111000000100000100",
			2166 => "0000000010001001101001",
			2167 => "0000000010001001101001",
			2168 => "0000111011000000000100",
			2169 => "0000000010001001101001",
			2170 => "0000000010001001101001",
			2171 => "0000000100110000000100",
			2172 => "0000000010001001101001",
			2173 => "0001011001101100000100",
			2174 => "0000000010001001101001",
			2175 => "0000000010001001101001",
			2176 => "0000010111110000000100",
			2177 => "0000000010001001101001",
			2178 => "0000000010001001101001",
			2179 => "0000101101110000101000",
			2180 => "0001101000110100010100",
			2181 => "0011111110001000001100",
			2182 => "0000011001100000000100",
			2183 => "0000000010001001101001",
			2184 => "0000010001100100000100",
			2185 => "0000000010001001101001",
			2186 => "0000000010001001101001",
			2187 => "0000011000011000000100",
			2188 => "0000000010001001101001",
			2189 => "0000000010001001101001",
			2190 => "0001111001010000000100",
			2191 => "0000000010001001101001",
			2192 => "0001110100101100001100",
			2193 => "0010001111001000001000",
			2194 => "0001001001000100000100",
			2195 => "0000000010001001101001",
			2196 => "0000000010001001101001",
			2197 => "0000000010001001101001",
			2198 => "0000000010001001101001",
			2199 => "0001111000101000000100",
			2200 => "0000000010001001101001",
			2201 => "0000000010001001101001",
			2202 => "0001011101001000100100",
			2203 => "0000100111111000011100",
			2204 => "0011010011110000000100",
			2205 => "0000000010001100100101",
			2206 => "0000111000000000001100",
			2207 => "0000111111011000001000",
			2208 => "0000110011000000000100",
			2209 => "0000000010001100100101",
			2210 => "0000000010001100100101",
			2211 => "0000000010001100100101",
			2212 => "0001001100101000000100",
			2213 => "0000000010001100100101",
			2214 => "0011100011101100000100",
			2215 => "0000000010001100100101",
			2216 => "0000000010001100100101",
			2217 => "0011110100110100000100",
			2218 => "0000000010001100100101",
			2219 => "0000000010001100100101",
			2220 => "0001011011000000010100",
			2221 => "0011100110110000001100",
			2222 => "0010011001000100001000",
			2223 => "0000000111101100000100",
			2224 => "0000000010001100100101",
			2225 => "0000000010001100100101",
			2226 => "0000000010001100100101",
			2227 => "0000000101010000000100",
			2228 => "0000000010001100100101",
			2229 => "0000000010001100100101",
			2230 => "0000110000111100011100",
			2231 => "0000100111000100001100",
			2232 => "0011100010001100001000",
			2233 => "0001101010100000000100",
			2234 => "0000000010001100100101",
			2235 => "0000000010001100100101",
			2236 => "0000000010001100100101",
			2237 => "0010000101101100000100",
			2238 => "0000000010001100100101",
			2239 => "0010100000111100000100",
			2240 => "0000000010001100100101",
			2241 => "0000111100101100000100",
			2242 => "0000000010001100100101",
			2243 => "0000000010001100100101",
			2244 => "0001011001101100001000",
			2245 => "0011111001011100000100",
			2246 => "0000000010001100100101",
			2247 => "0000000010001100100101",
			2248 => "0000000010001100100101",
			2249 => "0011001100101000110100",
			2250 => "0001100101001000010000",
			2251 => "0010000101101100000100",
			2252 => "1111111010001110010001",
			2253 => "0011011011101100001000",
			2254 => "0000001010001100000100",
			2255 => "1111111010001110010001",
			2256 => "0000010010001110010001",
			2257 => "1111111010001110010001",
			2258 => "0011100001000000100000",
			2259 => "0000110011001000001100",
			2260 => "0011010110110100001000",
			2261 => "0001111100110000000100",
			2262 => "1111111010001110010001",
			2263 => "0000001010001110010001",
			2264 => "1111111010001110010001",
			2265 => "0000010001100100010000",
			2266 => "0010101011111000001000",
			2267 => "0000000101101000000100",
			2268 => "0000000010001110010001",
			2269 => "0000001010001110010001",
			2270 => "0001011001101100000100",
			2271 => "0000001010001110010001",
			2272 => "1111111010001110010001",
			2273 => "1111111010001110010001",
			2274 => "1111111010001110010001",
			2275 => "1111111010001110010001",
			2276 => "0001011000000000001000",
			2277 => "0000111101001000000100",
			2278 => "0000000010010000100101",
			2279 => "0000000010010000100101",
			2280 => "0011100110110000110000",
			2281 => "0011101101100000011100",
			2282 => "0011101111110100010000",
			2283 => "0000000110111100001100",
			2284 => "0010101111101000000100",
			2285 => "0000000010010000100101",
			2286 => "0001011001011000000100",
			2287 => "0000000010010000100101",
			2288 => "0000000010010000100101",
			2289 => "0000000010010000100101",
			2290 => "0010111110011000000100",
			2291 => "0000000010010000100101",
			2292 => "0001000101111000000100",
			2293 => "1111111010010000100101",
			2294 => "0000000010010000100101",
			2295 => "0000010110010000000100",
			2296 => "0000000010010000100101",
			2297 => "0000111100010000000100",
			2298 => "0000000010010000100101",
			2299 => "0001011100101100000100",
			2300 => "0000000010010000100101",
			2301 => "0000001100100100000100",
			2302 => "0000000010010000100101",
			2303 => "0000000010010000100101",
			2304 => "0001000110000000001000",
			2305 => "0001001001001000000100",
			2306 => "0000000010010000100101",
			2307 => "0000000010010000100101",
			2308 => "0000001000001100000100",
			2309 => "0000000010010000100101",
			2310 => "0000001111010000000100",
			2311 => "0000000010010000100101",
			2312 => "0000000010010000100101",
			2313 => "0000101101011100111100",
			2314 => "0000110000111100110000",
			2315 => "0010110110001100001000",
			2316 => "0010110110110100000100",
			2317 => "0000000010010011100001",
			2318 => "0000000010010011100001",
			2319 => "0011011110011000011000",
			2320 => "0011100111001000010000",
			2321 => "0001111100000000001000",
			2322 => "0001001111011000000100",
			2323 => "0000000010010011100001",
			2324 => "0000000010010011100001",
			2325 => "0001000101010100000100",
			2326 => "0000000010010011100001",
			2327 => "0000000010010011100001",
			2328 => "0010101111101000000100",
			2329 => "0000000010010011100001",
			2330 => "0000000010010011100001",
			2331 => "0000001011111100000100",
			2332 => "0000000010010011100001",
			2333 => "0010010110000000001000",
			2334 => "0001100111101000000100",
			2335 => "0000000010010011100001",
			2336 => "0000000010010011100001",
			2337 => "0000000010010011100001",
			2338 => "0001011001101100001000",
			2339 => "0011111001011100000100",
			2340 => "0000000010010011100001",
			2341 => "0000000010010011100001",
			2342 => "0000000010010011100001",
			2343 => "0011100110110000010100",
			2344 => "0000010110010000001000",
			2345 => "0001001101101000000100",
			2346 => "0000000010010011100001",
			2347 => "0000000010010011100001",
			2348 => "0010101001010100000100",
			2349 => "0000000010010011100001",
			2350 => "0001011011111000000100",
			2351 => "0000000010010011100001",
			2352 => "0000000010010011100001",
			2353 => "0010111011101100000100",
			2354 => "0000000010010011100001",
			2355 => "0000010110010000000100",
			2356 => "0000000010010011100001",
			2357 => "0000011001100000000100",
			2358 => "0000000010010011100001",
			2359 => "0000000010010011100001",
			2360 => "0010110101010100111000",
			2361 => "0010000101101100101100",
			2362 => "0001011101001000010100",
			2363 => "0000000110111100000100",
			2364 => "1111111010010101010101",
			2365 => "0010000101011100001000",
			2366 => "0010010101011100000100",
			2367 => "0000000010010101010101",
			2368 => "0000001010010101010101",
			2369 => "0010011100101000000100",
			2370 => "0000000010010101010101",
			2371 => "1111111010010101010101",
			2372 => "0011011010100100010100",
			2373 => "0001100101001000000100",
			2374 => "1111111010010101010101",
			2375 => "0011010110001100001000",
			2376 => "0000001011100100000100",
			2377 => "0000000010010101010101",
			2378 => "0000001010010101010101",
			2379 => "0001011001101100000100",
			2380 => "0000001010010101010101",
			2381 => "0000000010010101010101",
			2382 => "1111111010010101010101",
			2383 => "0010101001011000000100",
			2384 => "1111111010010101010101",
			2385 => "0001001100101100000100",
			2386 => "0000001010010101010101",
			2387 => "1111111010010101010101",
			2388 => "1111111010010101010101",
			2389 => "0001001001000100011100",
			2390 => "0000111000000000010000",
			2391 => "0010101000111000001000",
			2392 => "0000110011001000000100",
			2393 => "0000000010011000010001",
			2394 => "0000000010011000010001",
			2395 => "0000111111011000000100",
			2396 => "0000000010011000010001",
			2397 => "0000000010011000010001",
			2398 => "0010010101101100001000",
			2399 => "0010001111111100000100",
			2400 => "0000000010011000010001",
			2401 => "0000000010011000010001",
			2402 => "0000000010011000010001",
			2403 => "0001000110000000001100",
			2404 => "0001101100000100000100",
			2405 => "0000000010011000010001",
			2406 => "0001111000101000000100",
			2407 => "0000000010011000010001",
			2408 => "0000000010011000010001",
			2409 => "0001110110101100011100",
			2410 => "0011101010110100001100",
			2411 => "0010000101101100000100",
			2412 => "0000000010011000010001",
			2413 => "0001111100000000000100",
			2414 => "0000000010011000010001",
			2415 => "0000000010011000010001",
			2416 => "0000010111100100001100",
			2417 => "0001101110010000001000",
			2418 => "0001101111110000000100",
			2419 => "0000000010011000010001",
			2420 => "0000000010011000010001",
			2421 => "0000000010011000010001",
			2422 => "0000000010011000010001",
			2423 => "0010111110011000000100",
			2424 => "0000000010011000010001",
			2425 => "0011100001000100001100",
			2426 => "0010101100110100000100",
			2427 => "0000000010011000010001",
			2428 => "0000100100011000000100",
			2429 => "0000000010011000010001",
			2430 => "0000000010011000010001",
			2431 => "0011101101100100001000",
			2432 => "0000010001100100000100",
			2433 => "0000000010011000010001",
			2434 => "0000000010011000010001",
			2435 => "0000000010011000010001",
			2436 => "0001011000000000001100",
			2437 => "0000111101001000000100",
			2438 => "1111111010011011000101",
			2439 => "0000111001010100000100",
			2440 => "0000000010011011000101",
			2441 => "0000000010011011000101",
			2442 => "0001100101100000101100",
			2443 => "0000000011001100100000",
			2444 => "0010101001000000010000",
			2445 => "0000010000011000001100",
			2446 => "0010110011010000001000",
			2447 => "0010101111101000000100",
			2448 => "0000000010011011000101",
			2449 => "0000000010011011000101",
			2450 => "0000000010011011000101",
			2451 => "1111111010011011000101",
			2452 => "0001011001101100001100",
			2453 => "0001010001111100001000",
			2454 => "0001011110010100000100",
			2455 => "0000000010011011000101",
			2456 => "0000000010011011000101",
			2457 => "0000001010011011000101",
			2458 => "0000000010011011000101",
			2459 => "0011001010100100000100",
			2460 => "0000000010011011000101",
			2461 => "0010011001000100000100",
			2462 => "0000001010011011000101",
			2463 => "0000000010011011000101",
			2464 => "0000001110110000011000",
			2465 => "0000111101001000001100",
			2466 => "0001000101111000001000",
			2467 => "0011111001111000000100",
			2468 => "0000000010011011000101",
			2469 => "1111111010011011000101",
			2470 => "0000000010011011000101",
			2471 => "0001100100100000001000",
			2472 => "0010011001000100000100",
			2473 => "0000001010011011000101",
			2474 => "0000000010011011000101",
			2475 => "0000000010011011000101",
			2476 => "0001111000101000001000",
			2477 => "0001110110101100000100",
			2478 => "0000000010011011000101",
			2479 => "0000001010011011000101",
			2480 => "0000000010011011000101",
			2481 => "0011000101011101000000",
			2482 => "0000000000101100001100",
			2483 => "0010000101101100000100",
			2484 => "1111111010011101001001",
			2485 => "0011000101010100000100",
			2486 => "1111111010011101001001",
			2487 => "0000001010011101001001",
			2488 => "0001110110101100010100",
			2489 => "0010111010100100010000",
			2490 => "0001100100000100001000",
			2491 => "0001011101001000000100",
			2492 => "1111111010011101001001",
			2493 => "0000000010011101001001",
			2494 => "0000110011001000000100",
			2495 => "0000000010011101001001",
			2496 => "0000001010011101001001",
			2497 => "0000001010011101001001",
			2498 => "0000101101110000010100",
			2499 => "0001000101111000001100",
			2500 => "0011101111110100000100",
			2501 => "0000000010011101001001",
			2502 => "0011100111001000000100",
			2503 => "1111111010011101001001",
			2504 => "0000000010011101001001",
			2505 => "0010011001000100000100",
			2506 => "0000001010011101001001",
			2507 => "1111111010011101001001",
			2508 => "0001111000101000001000",
			2509 => "0010011100101000000100",
			2510 => "0000001010011101001001",
			2511 => "0000000010011101001001",
			2512 => "1111111010011101001001",
			2513 => "1111111010011101001001",
			2514 => "0000110000111101000100",
			2515 => "0000011001100100010100",
			2516 => "0011001110011000000100",
			2517 => "1111111010011111101101",
			2518 => "0010011001001000001000",
			2519 => "0000111111011000000100",
			2520 => "0000000010011111101101",
			2521 => "0000001010011111101101",
			2522 => "0011011011101100000100",
			2523 => "1111111010011111101101",
			2524 => "0000000010011111101101",
			2525 => "0011011010100100100100",
			2526 => "0000011000011000100000",
			2527 => "0010101101001000010000",
			2528 => "0011001110011000001000",
			2529 => "0011001011101100000100",
			2530 => "0000000010011111101101",
			2531 => "1111111010011111101101",
			2532 => "0010000101011100000100",
			2533 => "0000000010011111101101",
			2534 => "0000000010011111101101",
			2535 => "0011111101001100001000",
			2536 => "0001001100101100000100",
			2537 => "0000001010011111101101",
			2538 => "1111111010011111101101",
			2539 => "0000001110110000000100",
			2540 => "1111111010011111101101",
			2541 => "0000000010011111101101",
			2542 => "1111111010011111101101",
			2543 => "0011101111010100000100",
			2544 => "1111111010011111101101",
			2545 => "0001100101100000000100",
			2546 => "0000000010011111101101",
			2547 => "0000000010011111101101",
			2548 => "0001011001101100001100",
			2549 => "0011111001011100000100",
			2550 => "0000000010011111101101",
			2551 => "0001100101100000000100",
			2552 => "0000001010011111101101",
			2553 => "0000000010011111101101",
			2554 => "0000000010011111101101",
			2555 => "0001110110101100110000",
			2556 => "0010101001010100011000",
			2557 => "0011001010100100001100",
			2558 => "0001001001000100000100",
			2559 => "0000000010100011001001",
			2560 => "0000011000011000000100",
			2561 => "0000000010100011001001",
			2562 => "0000000010100011001001",
			2563 => "0001111100010000000100",
			2564 => "0000000010100011001001",
			2565 => "0000111111011000000100",
			2566 => "0000000010100011001001",
			2567 => "0000000010100011001001",
			2568 => "0011101010110100001100",
			2569 => "0010000101101100000100",
			2570 => "0000000010100011001001",
			2571 => "0011100010001100000100",
			2572 => "0000000010100011001001",
			2573 => "0000000010100011001001",
			2574 => "0000100111000100001000",
			2575 => "0011100100100100000100",
			2576 => "0000000010100011001001",
			2577 => "0000000010100011001001",
			2578 => "0000000010100011001001",
			2579 => "0000001110110000110100",
			2580 => "0001000101111000011100",
			2581 => "0001011100101100011000",
			2582 => "0001100000001100010000",
			2583 => "0011100101110100001000",
			2584 => "0010111010100100000100",
			2585 => "0000000010100011001001",
			2586 => "0000000010100011001001",
			2587 => "0000100010100100000100",
			2588 => "0000000010100011001001",
			2589 => "0000000010100011001001",
			2590 => "0010111110011000000100",
			2591 => "0000000010100011001001",
			2592 => "0000000010100011001001",
			2593 => "0000000010100011001001",
			2594 => "0010010101101100000100",
			2595 => "0000000010100011001001",
			2596 => "0000011001100000001000",
			2597 => "0011100010110000000100",
			2598 => "0000000010100011001001",
			2599 => "0000000010100011001001",
			2600 => "0000010001100100001000",
			2601 => "0010001001000100000100",
			2602 => "0000000010100011001001",
			2603 => "0000000010100011001001",
			2604 => "0000000010100011001001",
			2605 => "0011100001000000001000",
			2606 => "0010111010100100000100",
			2607 => "0000000010100011001001",
			2608 => "0000000010100011001001",
			2609 => "0000000010100011001001",
			2610 => "0011100110110001000000",
			2611 => "0001100000010000111100",
			2612 => "0001010110101100011000",
			2613 => "0000111000000000010000",
			2614 => "0011010110110100001100",
			2615 => "0011011111011100000100",
			2616 => "0000000010100101101101",
			2617 => "0000110011000000000100",
			2618 => "0000000010100101101101",
			2619 => "0000000010100101101101",
			2620 => "1111111010100101101101",
			2621 => "0010001111111100000100",
			2622 => "0000000010100101101101",
			2623 => "0000000010100101101101",
			2624 => "0011011010100100010100",
			2625 => "0010000101101100001100",
			2626 => "0000001011100100001000",
			2627 => "0011010110001100000100",
			2628 => "0000000010100101101101",
			2629 => "0000000010100101101101",
			2630 => "0000001010100101101101",
			2631 => "0011100010001100000100",
			2632 => "0000000010100101101101",
			2633 => "0000000010100101101101",
			2634 => "0000011001100000000100",
			2635 => "0000000010100101101101",
			2636 => "0000010001100100001000",
			2637 => "0000111011111000000100",
			2638 => "0000000010100101101101",
			2639 => "0000000010100101101101",
			2640 => "0000000010100101101101",
			2641 => "0000000010100101101101",
			2642 => "0010111011101100001000",
			2643 => "0011110111001100000100",
			2644 => "0000000010100101101101",
			2645 => "0000000010100101101101",
			2646 => "0000010110010000000100",
			2647 => "0000000010100101101101",
			2648 => "0000011000011000000100",
			2649 => "0000000010100101101101",
			2650 => "0000000010100101101101",
			2651 => "0011111001011100000100",
			2652 => "1111111010100111110001",
			2653 => "0011100110110000110000",
			2654 => "0011001110011000001100",
			2655 => "0011010110001100001000",
			2656 => "0011110100011000000100",
			2657 => "1111111010100111110001",
			2658 => "0000000010100111110001",
			2659 => "0000001010100111110001",
			2660 => "0010001001001100010000",
			2661 => "0001011000000100000100",
			2662 => "0000000010100111110001",
			2663 => "0010111110011000000100",
			2664 => "0000000010100111110001",
			2665 => "0000111001000000000100",
			2666 => "0000001010100111110001",
			2667 => "0000000010100111110001",
			2668 => "0000001001101000010000",
			2669 => "0010101001011000001000",
			2670 => "0010011001001000000100",
			2671 => "0000000010100111110001",
			2672 => "1111111010100111110001",
			2673 => "0011101010011000000100",
			2674 => "1111111010100111110001",
			2675 => "0000001010100111110001",
			2676 => "0000001010100111110001",
			2677 => "0010111110011000001100",
			2678 => "0010010101011100000100",
			2679 => "1111111010100111110001",
			2680 => "0011111000100100000100",
			2681 => "0000000010100111110001",
			2682 => "0000000010100111110001",
			2683 => "1111111010100111110001",
			2684 => "0011000101011101000100",
			2685 => "0000000000101100010000",
			2686 => "0010000101101100000100",
			2687 => "1111111010101001111101",
			2688 => "0010001001000100001000",
			2689 => "0011011011101100000100",
			2690 => "0000001010101001111101",
			2691 => "0000000010101001111101",
			2692 => "1111111010101001111101",
			2693 => "0001110110101100010100",
			2694 => "0001000101010100000100",
			2695 => "1111111010101001111101",
			2696 => "0010111010100100001100",
			2697 => "0011101111000100000100",
			2698 => "1111111010101001111101",
			2699 => "0010101101001000000100",
			2700 => "0000000010101001111101",
			2701 => "0000001010101001111101",
			2702 => "0000001010101001111101",
			2703 => "0000001110110000010100",
			2704 => "0010101001011000001100",
			2705 => "0011101111110100000100",
			2706 => "0000000010101001111101",
			2707 => "0000100000101000000100",
			2708 => "0000000010101001111101",
			2709 => "1111111010101001111101",
			2710 => "0010011001000100000100",
			2711 => "0000001010101001111101",
			2712 => "1111111010101001111101",
			2713 => "0001111000101000001000",
			2714 => "0010011100101000000100",
			2715 => "0000001010101001111101",
			2716 => "0000001010101001111101",
			2717 => "1111111010101001111101",
			2718 => "1111111010101001111101",
			2719 => "0010001010100100001000",
			2720 => "0010010101010100000100",
			2721 => "0000000010101100001001",
			2722 => "0000000010101100001001",
			2723 => "0001011000000000001000",
			2724 => "0000111101001000000100",
			2725 => "0000000010101100001001",
			2726 => "0000000010101100001001",
			2727 => "0000000101101000101100",
			2728 => "0001110110101100010000",
			2729 => "0000011000011000001100",
			2730 => "0000100010100100001000",
			2731 => "0010101001000000000100",
			2732 => "0000000010101100001001",
			2733 => "0000000010101100001001",
			2734 => "0000000010101100001001",
			2735 => "0000000010101100001001",
			2736 => "0001101000110100001100",
			2737 => "0001100001100000001000",
			2738 => "0000011001100000000100",
			2739 => "0000000010101100001001",
			2740 => "0000000010101100001001",
			2741 => "0000000010101100001001",
			2742 => "0000111111101000001000",
			2743 => "0001101010111100000100",
			2744 => "0000000010101100001001",
			2745 => "0000000010101100001001",
			2746 => "0011101110100000000100",
			2747 => "0000000010101100001001",
			2748 => "0000000010101100001001",
			2749 => "0011011011101100000100",
			2750 => "0000000010101100001001",
			2751 => "0001000110000000000100",
			2752 => "0000000010101100001001",
			2753 => "0000000010101100001001",
			2754 => "0011010011010001000100",
			2755 => "0000110011001000001100",
			2756 => "0011010110110100001000",
			2757 => "0010111110011000000100",
			2758 => "1111111010101110010101",
			2759 => "0000001010101110010101",
			2760 => "1111111010101110010101",
			2761 => "0011100110110000101000",
			2762 => "0011001110011000001000",
			2763 => "0001100101001100000100",
			2764 => "1111111010101110010101",
			2765 => "0000001010101110010101",
			2766 => "0000100111000100010000",
			2767 => "0000110011000100001000",
			2768 => "0001100100101000000100",
			2769 => "1111111010101110010101",
			2770 => "0000000010101110010101",
			2771 => "0001011001101100000100",
			2772 => "0000001010101110010101",
			2773 => "1111111010101110010101",
			2774 => "0010000101101100001000",
			2775 => "0000111101001000000100",
			2776 => "0000000010101110010101",
			2777 => "0000001010101110010101",
			2778 => "0000111000101000000100",
			2779 => "1111111010101110010101",
			2780 => "0000000010101110010101",
			2781 => "0010111110011000001000",
			2782 => "0000001111001100000100",
			2783 => "1111111010101110010101",
			2784 => "0000001010101110010101",
			2785 => "0000001010111000000100",
			2786 => "1111111010101110010101",
			2787 => "0000000010101110010101",
			2788 => "1111111010101110010101",
			2789 => "0011010011010000110000",
			2790 => "0001011000000100000100",
			2791 => "1111111010101111111001",
			2792 => "0011100001000000101000",
			2793 => "0001111100010000010100",
			2794 => "0001011100010000000100",
			2795 => "1111111010101111111001",
			2796 => "0001011011000000001000",
			2797 => "0000000100110100000100",
			2798 => "1111111010101111111001",
			2799 => "0000001010101111111001",
			2800 => "0010011101101000000100",
			2801 => "1111111010101111111001",
			2802 => "0000000010101111111001",
			2803 => "0000001001101000010000",
			2804 => "0001110110101100001000",
			2805 => "0011011010100100000100",
			2806 => "0000001010101111111001",
			2807 => "1111111010101111111001",
			2808 => "0010010101011100000100",
			2809 => "0000000010101111111001",
			2810 => "0000000010101111111001",
			2811 => "0000001010101111111001",
			2812 => "1111111010101111111001",
			2813 => "1111111010101111111001",
			2814 => "0011010011010001001000",
			2815 => "0001011000000000001000",
			2816 => "0000111101001000000100",
			2817 => "1111111010110010001111",
			2818 => "0000000010110010001111",
			2819 => "0010010101101100011100",
			2820 => "0010000101101100010100",
			2821 => "0000000101101000010000",
			2822 => "0010101011111000001000",
			2823 => "0001111101001000000100",
			2824 => "0000000010110010001111",
			2825 => "0000000010110010001111",
			2826 => "0001001100110000000100",
			2827 => "0000001010110010001111",
			2828 => "0000000010110010001111",
			2829 => "0000001010110010001111",
			2830 => "0011101111010100000100",
			2831 => "0000000010110010001111",
			2832 => "1111111010110010001111",
			2833 => "0010101100001100011000",
			2834 => "0010111010100100001000",
			2835 => "0000010111110000000100",
			2836 => "0000001010110010001111",
			2837 => "1111111010110010001111",
			2838 => "0011100010001100001000",
			2839 => "0010000101101100000100",
			2840 => "1111111010110010001111",
			2841 => "0000001010110010001111",
			2842 => "0001111111101000000100",
			2843 => "1111111010110010001111",
			2844 => "0000000010110010001111",
			2845 => "0010001111111100000100",
			2846 => "1111111010110010001111",
			2847 => "0000111110001100000100",
			2848 => "0000001010110010001111",
			2849 => "0000000010110010001111",
			2850 => "1111111010110010001111",
			2851 => "0010010101101100101000",
			2852 => "0001011000000000001100",
			2853 => "0010001010100100000100",
			2854 => "0000000010110100010001",
			2855 => "0000111100110000000100",
			2856 => "0000000010110100010001",
			2857 => "0000000010110100010001",
			2858 => "0011001110011000001000",
			2859 => "0001100101001100000100",
			2860 => "0000000010110100010001",
			2861 => "0000000010110100010001",
			2862 => "0000011000011000010000",
			2863 => "0000001011111100000100",
			2864 => "0000000010110100010001",
			2865 => "0001100101001100000100",
			2866 => "0000000010110100010001",
			2867 => "0011111011010100000100",
			2868 => "0000000010110100010001",
			2869 => "0000000010110100010001",
			2870 => "0000000010110100010001",
			2871 => "0010001001001100001000",
			2872 => "0011111001011100000100",
			2873 => "0000000010110100010001",
			2874 => "0000000010110100010001",
			2875 => "0011100010001100001000",
			2876 => "0000000100110000000100",
			2877 => "0000000010110100010001",
			2878 => "0000000010110100010001",
			2879 => "0010101100110100000100",
			2880 => "0000000010110100010001",
			2881 => "0010100000111000000100",
			2882 => "0000000010110100010001",
			2883 => "0000000010110100010001",
			2884 => "0000000011001100011100",
			2885 => "0010101001000000010000",
			2886 => "0010001010100100000100",
			2887 => "0000000010110110100101",
			2888 => "0001111100000000001000",
			2889 => "0001111000000100000100",
			2890 => "0000000010110110100101",
			2891 => "0000000010110110100101",
			2892 => "0000000010110110100101",
			2893 => "0000010110010000000100",
			2894 => "0000000010110110100101",
			2895 => "0010010011000000000100",
			2896 => "0000000010110110100101",
			2897 => "0000000010110110100101",
			2898 => "0010101101001000010000",
			2899 => "0001011100110000001100",
			2900 => "0011011110011000001000",
			2901 => "0001100100100000000100",
			2902 => "0000000010110110100101",
			2903 => "0000000010110110100101",
			2904 => "0000000010110110100101",
			2905 => "0000000010110110100101",
			2906 => "0011100110110000010100",
			2907 => "0000010110010000001000",
			2908 => "0000011001100100000100",
			2909 => "0000000010110110100101",
			2910 => "0000000010110110100101",
			2911 => "0011110010111100000100",
			2912 => "0000000010110110100101",
			2913 => "0000100111111000000100",
			2914 => "0000000010110110100101",
			2915 => "0000000010110110100101",
			2916 => "0010111110011000001000",
			2917 => "0011110111001100000100",
			2918 => "0000000010110110100101",
			2919 => "0000000010110110100101",
			2920 => "0000000010110110100101",
			2921 => "0001011000000000001000",
			2922 => "0000111101001000000100",
			2923 => "1111111010111000000001",
			2924 => "0000000010111000000001",
			2925 => "0000001110110000100000",
			2926 => "0011111101001100011100",
			2927 => "0000101100100100010000",
			2928 => "0011111100111100001100",
			2929 => "0010010101011100000100",
			2930 => "0000000010111000000001",
			2931 => "0000000011001100000100",
			2932 => "0000000010111000000001",
			2933 => "0000001010111000000001",
			2934 => "1111111010111000000001",
			2935 => "0000010110010000000100",
			2936 => "0000001010111000000001",
			2937 => "0011111011110100000100",
			2938 => "1111111010111000000001",
			2939 => "0000000010111000000001",
			2940 => "1111111010111000000001",
			2941 => "0001111000101000000100",
			2942 => "0000001010111000000001",
			2943 => "1111111010111000000001",
			2944 => "0010011001000100100100",
			2945 => "0000001011111100001000",
			2946 => "0000111111101000000100",
			2947 => "1111111010111001101101",
			2948 => "0000000010111001101101",
			2949 => "0011100100101000011000",
			2950 => "0001011000000100000100",
			2951 => "1111111010111001101101",
			2952 => "0000011000011000010000",
			2953 => "0010101000101000001000",
			2954 => "0000100111111000000100",
			2955 => "0000000010111001101101",
			2956 => "0000010010111001101101",
			2957 => "0011111101001100000100",
			2958 => "0000001010111001101101",
			2959 => "0000001010111001101101",
			2960 => "0000000010111001101101",
			2961 => "1111111010111001101101",
			2962 => "0011001100101000010000",
			2963 => "0010101001000000000100",
			2964 => "1111111010111001101101",
			2965 => "0001011001101100001000",
			2966 => "0011111101000100000100",
			2967 => "0000000010111001101101",
			2968 => "0000010010111001101101",
			2969 => "1111111010111001101101",
			2970 => "1111111010111001101101",
			2971 => "0011001100101000100100",
			2972 => "0010101000111000001000",
			2973 => "0011101100011000000100",
			2974 => "1111111010111010111001",
			2975 => "0000000010111010111001",
			2976 => "0000011000111100000100",
			2977 => "1111111010111010111001",
			2978 => "0011100001000000010100",
			2979 => "0000010001100100010000",
			2980 => "0000000101101000001000",
			2981 => "0001001010000100000100",
			2982 => "0000000010111010111001",
			2983 => "0000000010111010111001",
			2984 => "0010001111111100000100",
			2985 => "0000001010111010111001",
			2986 => "0000000010111010111001",
			2987 => "1111111010111010111001",
			2988 => "1111111010111010111001",
			2989 => "1111111010111010111001",
			2990 => "0011001100101000101000",
			2991 => "0010101000111000001100",
			2992 => "0011101100011000001000",
			2993 => "0011110100011000000100",
			2994 => "1111111010111100001101",
			2995 => "1111111010111100001101",
			2996 => "0000000010111100001101",
			2997 => "0000011000111100000100",
			2998 => "1111111010111100001101",
			2999 => "0011100001000000010100",
			3000 => "0000010001100100010000",
			3001 => "0001101100100000001000",
			3002 => "0001000110011100000100",
			3003 => "0000000010111100001101",
			3004 => "1111111010111100001101",
			3005 => "0010000101101100000100",
			3006 => "0000001010111100001101",
			3007 => "0000000010111100001101",
			3008 => "1111111010111100001101",
			3009 => "1111111010111100001101",
			3010 => "1111111010111100001101",
			3011 => "0001001001000100010100",
			3012 => "0000111000000000001100",
			3013 => "0010101000111000001000",
			3014 => "0000110011001000000100",
			3015 => "0000000010111110100001",
			3016 => "0000000010111110100001",
			3017 => "0000000010111110100001",
			3018 => "0001111001010000000100",
			3019 => "0000000010111110100001",
			3020 => "0000000010111110100001",
			3021 => "0010000101101100101000",
			3022 => "0000001101110000100000",
			3023 => "0010101011111000010000",
			3024 => "0011011011101100001000",
			3025 => "0011010110110100000100",
			3026 => "0000000010111110100001",
			3027 => "0000000010111110100001",
			3028 => "0000111101001000000100",
			3029 => "0000000010111110100001",
			3030 => "0000000010111110100001",
			3031 => "0001100101001000000100",
			3032 => "0000000010111110100001",
			3033 => "0011011010100100001000",
			3034 => "0010110101010100000100",
			3035 => "0000000010111110100001",
			3036 => "0000000010111110100001",
			3037 => "0000000010111110100001",
			3038 => "0001111101001000000100",
			3039 => "0000000010111110100001",
			3040 => "0000000010111110100001",
			3041 => "0000001101001100001100",
			3042 => "0000000100110000000100",
			3043 => "0000000010111110100001",
			3044 => "0001000011000100000100",
			3045 => "0000000010111110100001",
			3046 => "0000000010111110100001",
			3047 => "0000000010111110100001",
			3048 => "0010000101101101000000",
			3049 => "0000100111000100010100",
			3050 => "0000110000111100001100",
			3051 => "0011001110011000001000",
			3052 => "0010001111111100000100",
			3053 => "1111111011000001000101",
			3054 => "0000001011000001000101",
			3055 => "1111111011000001000101",
			3056 => "0001011001101100000100",
			3057 => "0000001011000001000101",
			3058 => "1111111011000001000101",
			3059 => "0000111000000000010100",
			3060 => "0011010110001100001100",
			3061 => "0001001001000100001000",
			3062 => "0010010101010100000100",
			3063 => "1111111011000001000101",
			3064 => "0000000011000001000101",
			3065 => "0000001011000001000101",
			3066 => "0001111001010100000100",
			3067 => "1111111011000001000101",
			3068 => "0000000011000001000101",
			3069 => "0011100110110000010000",
			3070 => "0011001110011000000100",
			3071 => "0000001011000001000101",
			3072 => "0001100100110000000100",
			3073 => "0000001011000001000101",
			3074 => "0011111100111100000100",
			3075 => "0000001011000001000101",
			3076 => "0000001011000001000101",
			3077 => "0011010110001100000100",
			3078 => "0000000011000001000101",
			3079 => "0000001011000001000101",
			3080 => "0000010000011000001000",
			3081 => "0010011010000100000100",
			3082 => "0000000011000001000101",
			3083 => "1111111011000001000101",
			3084 => "0000111011111000000100",
			3085 => "1111111011000001000101",
			3086 => "0001011001011000000100",
			3087 => "0000001011000001000101",
			3088 => "1111111011000001000101",
			3089 => "0001011101001000101000",
			3090 => "0000111000000000011000",
			3091 => "0001001001000100001100",
			3092 => "0000111111011000001000",
			3093 => "0000110011000000000100",
			3094 => "0000000011000011111001",
			3095 => "0000000011000011111001",
			3096 => "1111111011000011111001",
			3097 => "0011010110001100000100",
			3098 => "0000000011000011111001",
			3099 => "0001111001010000000100",
			3100 => "1111111011000011111001",
			3101 => "0000000011000011111001",
			3102 => "0001001001001000001000",
			3103 => "0000000110111100000100",
			3104 => "0000000011000011111001",
			3105 => "0000000011000011111001",
			3106 => "0001011100110000000100",
			3107 => "0000000011000011111001",
			3108 => "0000000011000011111001",
			3109 => "0001001111011000010000",
			3110 => "0010000101101100001100",
			3111 => "0011101100011000001000",
			3112 => "0011101111110000000100",
			3113 => "0000000011000011111001",
			3114 => "0000001011000011111001",
			3115 => "0000000011000011111001",
			3116 => "0000000011000011111001",
			3117 => "0010101001011000001000",
			3118 => "0010011001001000000100",
			3119 => "0000000011000011111001",
			3120 => "1111111011000011111001",
			3121 => "0001001001010000001000",
			3122 => "0010010110000000000100",
			3123 => "0000000011000011111001",
			3124 => "0000000011000011111001",
			3125 => "0000110000111100001000",
			3126 => "0011100001011100000100",
			3127 => "0000000011000011111001",
			3128 => "1111111011000011111001",
			3129 => "0001011001101100001000",
			3130 => "0011111001011100000100",
			3131 => "0000000011000011111001",
			3132 => "0000000011000011111001",
			3133 => "0000000011000011111001",
			3134 => "0011011011101100110000",
			3135 => "0011100110110000101000",
			3136 => "0000001101110000100000",
			3137 => "0010101011111000010000",
			3138 => "0010110110001100000100",
			3139 => "0000000011000110001101",
			3140 => "0010110011010000001000",
			3141 => "0001000101010100000100",
			3142 => "0000000011000110001101",
			3143 => "0000000011000110001101",
			3144 => "0000000011000110001101",
			3145 => "0010011010000100001100",
			3146 => "0001100100000000000100",
			3147 => "0000000011000110001101",
			3148 => "0001011001101100000100",
			3149 => "0000000011000110001101",
			3150 => "0000000011000110001101",
			3151 => "0000000011000110001101",
			3152 => "0000010111110000000100",
			3153 => "0000000011000110001101",
			3154 => "0000000011000110001101",
			3155 => "0010111011101100000100",
			3156 => "0000000011000110001101",
			3157 => "0000000011000110001101",
			3158 => "0010001001001100001000",
			3159 => "0011110101001100000100",
			3160 => "0000000011000110001101",
			3161 => "0000000011000110001101",
			3162 => "0010101100110100001100",
			3163 => "0010111110011000001000",
			3164 => "0011001110011000000100",
			3165 => "0000000011000110001101",
			3166 => "0000000011000110001101",
			3167 => "0000000011000110001101",
			3168 => "0000110011110100000100",
			3169 => "0000000011000110001101",
			3170 => "0000000011000110001101",
			3171 => "0010011001000100100100",
			3172 => "0000000111101100000100",
			3173 => "1111111011000111111001",
			3174 => "0011100001000000011100",
			3175 => "0001011000000100000100",
			3176 => "1111111011000111111001",
			3177 => "0010101011111000010000",
			3178 => "0000001110110000001000",
			3179 => "0001111101001000000100",
			3180 => "0000001011000111111001",
			3181 => "0000000011000111111001",
			3182 => "0001011101001000000100",
			3183 => "0000001011000111111001",
			3184 => "0000001011000111111001",
			3185 => "0001010011000100000100",
			3186 => "0000001011000111111001",
			3187 => "0000001011000111111001",
			3188 => "1111111011000111111001",
			3189 => "0011001100101000010000",
			3190 => "0010101001000000000100",
			3191 => "1111111011000111111001",
			3192 => "0001011001101100001000",
			3193 => "0010001111111100000100",
			3194 => "0000000011000111111001",
			3195 => "0000001011000111111001",
			3196 => "1111111011000111111001",
			3197 => "1111111011000111111001",
			3198 => "0011100110110000111000",
			3199 => "0001011101001000010000",
			3200 => "0000000110111100000100",
			3201 => "1111111011001010000101",
			3202 => "0000010110010000001000",
			3203 => "0000100110100100000100",
			3204 => "0000000011001010000101",
			3205 => "0000000011001010000101",
			3206 => "1111111011001010000101",
			3207 => "0001011001010000001000",
			3208 => "0011101111110000000100",
			3209 => "0000000011001010000101",
			3210 => "0000001011001010000101",
			3211 => "0001010001010000001000",
			3212 => "0001110110101100000100",
			3213 => "0000000011001010000101",
			3214 => "1111111011001010000101",
			3215 => "0000100111000100001100",
			3216 => "0001101111110000001000",
			3217 => "0001101100100000000100",
			3218 => "0000000011001010000101",
			3219 => "0000001011001010000101",
			3220 => "1111111011001010000101",
			3221 => "0010000101101100000100",
			3222 => "0000001011001010000101",
			3223 => "0000111111101000000100",
			3224 => "1111111011001010000101",
			3225 => "0000001011001010000101",
			3226 => "0000010001110000000100",
			3227 => "1111111011001010000101",
			3228 => "0011100001000000001000",
			3229 => "0010010101101100000100",
			3230 => "0000001011001010000101",
			3231 => "0000000011001010000101",
			3232 => "1111111011001010000101",
			3233 => "0011100110110001000000",
			3234 => "0000001101110100011100",
			3235 => "0001111100000000001100",
			3236 => "0000000100110000000100",
			3237 => "0000000011001100011001",
			3238 => "0010001111111100000100",
			3239 => "0000000011001100011001",
			3240 => "0000000011001100011001",
			3241 => "0001010001111100000100",
			3242 => "0000000011001100011001",
			3243 => "0000010110010000000100",
			3244 => "0000000011001100011001",
			3245 => "0001010001011100000100",
			3246 => "0000000011001100011001",
			3247 => "0000000011001100011001",
			3248 => "0011001110011000001000",
			3249 => "0001100101001100000100",
			3250 => "0000000011001100011001",
			3251 => "0000000011001100011001",
			3252 => "0000011000011000010000",
			3253 => "0010000101101100001100",
			3254 => "0000110011100100001000",
			3255 => "0011010110001100000100",
			3256 => "0000000011001100011001",
			3257 => "0000000011001100011001",
			3258 => "0000000011001100011001",
			3259 => "0000000011001100011001",
			3260 => "0001111111101000000100",
			3261 => "0000000011001100011001",
			3262 => "0001011100101100000100",
			3263 => "0000000011001100011001",
			3264 => "0000000011001100011001",
			3265 => "0010111011101100001000",
			3266 => "0000011001100000000100",
			3267 => "0000000011001100011001",
			3268 => "0000000011001100011001",
			3269 => "0000000011001100011001",
			3270 => "0000101101011100110100",
			3271 => "0011001110011000001000",
			3272 => "0001001010000100000100",
			3273 => "0000000011001110111101",
			3274 => "0000000011001110111101",
			3275 => "0010001001001100010000",
			3276 => "0011111001011100000100",
			3277 => "0000000011001110111101",
			3278 => "0000110011100100000100",
			3279 => "0000000011001110111101",
			3280 => "0001001001011000000100",
			3281 => "0000000011001110111101",
			3282 => "0000000011001110111101",
			3283 => "0010101100001100010000",
			3284 => "0000001011111100000100",
			3285 => "0000000011001110111101",
			3286 => "0001100111101000001000",
			3287 => "0010010110000000000100",
			3288 => "0000000011001110111101",
			3289 => "0000000011001110111101",
			3290 => "0000000011001110111101",
			3291 => "0000000100111100001000",
			3292 => "0011111111110000000100",
			3293 => "0000000011001110111101",
			3294 => "0000000011001110111101",
			3295 => "0000000011001110111101",
			3296 => "0011100110110000010000",
			3297 => "0000010110010000000100",
			3298 => "0000000011001110111101",
			3299 => "0010101001010100000100",
			3300 => "0000000011001110111101",
			3301 => "0001011011111000000100",
			3302 => "0000000011001110111101",
			3303 => "0000000011001110111101",
			3304 => "0010111011101100000100",
			3305 => "0000000011001110111101",
			3306 => "0000010110010000000100",
			3307 => "0000000011001110111101",
			3308 => "0000011001100000000100",
			3309 => "0000000011001110111101",
			3310 => "0000000011001110111101",
			3311 => "0010101001010100011100",
			3312 => "0011111011000100010000",
			3313 => "0001010110101100000100",
			3314 => "1111111011010001101001",
			3315 => "0001001101101000000100",
			3316 => "0000000011010001101001",
			3317 => "0011000011010000000100",
			3318 => "0000000011010001101001",
			3319 => "0000000011010001101001",
			3320 => "0011100110110000000100",
			3321 => "0000000011010001101001",
			3322 => "0010111011101100000100",
			3323 => "0000000011010001101001",
			3324 => "0000000011010001101001",
			3325 => "0000101101011100101000",
			3326 => "0001010001111100100000",
			3327 => "0011101001011100001100",
			3328 => "0011100010001100001000",
			3329 => "0010000101101100000100",
			3330 => "0000000011010001101001",
			3331 => "0000000011010001101001",
			3332 => "1111111011010001101001",
			3333 => "0001110110101100000100",
			3334 => "0000000011010001101001",
			3335 => "0011111010110000001000",
			3336 => "0001001111011000000100",
			3337 => "0000000011010001101001",
			3338 => "0000000011010001101001",
			3339 => "0000000000000000000100",
			3340 => "1111111011010001101001",
			3341 => "0000000011010001101001",
			3342 => "0001011001101100000100",
			3343 => "0000000011010001101001",
			3344 => "0000000011010001101001",
			3345 => "0010000101101100001000",
			3346 => "0011101110100000000100",
			3347 => "0000001011010001101001",
			3348 => "0000000011010001101001",
			3349 => "0010100000111100000100",
			3350 => "0000000011010001101001",
			3351 => "0000111100101100000100",
			3352 => "0000000011010001101001",
			3353 => "0000000011010001101001",
			3354 => "0001011000000000001000",
			3355 => "0000111101001000000100",
			3356 => "0000000011010011101101",
			3357 => "0000000011010011101101",
			3358 => "0010000101101100101100",
			3359 => "0000000101101000100000",
			3360 => "0001110110101100010000",
			3361 => "0011101010110100000100",
			3362 => "0000000011010011101101",
			3363 => "0010101001010100000100",
			3364 => "0000000011010011101101",
			3365 => "0001001001010000000100",
			3366 => "0000000011010011101101",
			3367 => "0000000011010011101101",
			3368 => "0001101000110100001000",
			3369 => "0000001011111100000100",
			3370 => "0000000011010011101101",
			3371 => "0000000011010011101101",
			3372 => "0001101010111100000100",
			3373 => "0000000011010011101101",
			3374 => "0000000011010011101101",
			3375 => "0001001010000100000100",
			3376 => "0000000011010011101101",
			3377 => "0001000101111000000100",
			3378 => "0000000011010011101101",
			3379 => "0000000011010011101101",
			3380 => "0000100100011000001100",
			3381 => "0000110011000100000100",
			3382 => "0000000011010011101101",
			3383 => "0001000011000100000100",
			3384 => "0000000011010011101101",
			3385 => "0000000011010011101101",
			3386 => "0000000011010011101101",
			3387 => "0011100110110001000000",
			3388 => "0000001101110000101100",
			3389 => "0001011101001000010100",
			3390 => "0011000111011100001100",
			3391 => "0010110110001100001000",
			3392 => "0001100111010100000100",
			3393 => "0000000011010110001001",
			3394 => "0000000011010110001001",
			3395 => "1111111011010110001001",
			3396 => "0010010101101100000100",
			3397 => "0000001011010110001001",
			3398 => "0000000011010110001001",
			3399 => "0001000011000100010100",
			3400 => "0001010001111100010000",
			3401 => "0011101001011100001000",
			3402 => "0001111100000000000100",
			3403 => "0000000011010110001001",
			3404 => "1111111011010110001001",
			3405 => "0010010110000000000100",
			3406 => "0000000011010110001001",
			3407 => "0000000011010110001001",
			3408 => "0000001011010110001001",
			3409 => "1111111011010110001001",
			3410 => "0011011011101100001000",
			3411 => "0000010111110000000100",
			3412 => "0000001011010110001001",
			3413 => "0000000011010110001001",
			3414 => "0010101001010100000100",
			3415 => "1111111011010110001001",
			3416 => "0001011011111000000100",
			3417 => "0000000011010110001001",
			3418 => "0000000011010110001001",
			3419 => "0010011001001000001100",
			3420 => "0000000101010000001000",
			3421 => "0010101111101000000100",
			3422 => "1111111011010110001001",
			3423 => "0000000011010110001001",
			3424 => "0000000011010110001001",
			3425 => "1111111011010110001001",
			3426 => "0001011101001000101000",
			3427 => "0000111000000000011000",
			3428 => "0001001001000100001100",
			3429 => "0000111111011000001000",
			3430 => "0000110011000000000100",
			3431 => "0000000011011000111101",
			3432 => "0000000011011000111101",
			3433 => "1111111011011000111101",
			3434 => "0011010110001100000100",
			3435 => "0000000011011000111101",
			3436 => "0001111001010000000100",
			3437 => "1111111011011000111101",
			3438 => "0000000011011000111101",
			3439 => "0001001001001000001000",
			3440 => "0000000110111100000100",
			3441 => "0000000011011000111101",
			3442 => "0000000011011000111101",
			3443 => "0001011100110000000100",
			3444 => "0000000011011000111101",
			3445 => "0000000011011000111101",
			3446 => "0011001010100100001000",
			3447 => "0001001100000000000100",
			3448 => "0000001011011000111101",
			3449 => "0000000011011000111101",
			3450 => "0010001001001100001100",
			3451 => "0011111001011100000100",
			3452 => "0000000011011000111101",
			3453 => "0010101110111000000100",
			3454 => "0000000011011000111101",
			3455 => "0000000011011000111101",
			3456 => "0010101100001100011000",
			3457 => "0001001001010000010000",
			3458 => "0010101001011000001000",
			3459 => "0010010101101100000100",
			3460 => "0000000011011000111101",
			3461 => "0000000011011000111101",
			3462 => "0010011101101000000100",
			3463 => "0000000011011000111101",
			3464 => "0000000011011000111101",
			3465 => "0011100010001100000100",
			3466 => "0000000011011000111101",
			3467 => "1111111011011000111101",
			3468 => "0001011001101100000100",
			3469 => "0000000011011000111101",
			3470 => "0000000011011000111101",
			3471 => "0001011000000000001000",
			3472 => "0000111101001000000100",
			3473 => "0000000011011011000001",
			3474 => "0000000011011011000001",
			3475 => "0010000101101100101000",
			3476 => "0000101101110000100000",
			3477 => "0001110110101100010000",
			3478 => "0011101010110100000100",
			3479 => "0000000011011011000001",
			3480 => "0010101001010100000100",
			3481 => "0000000011011011000001",
			3482 => "0001001001010000000100",
			3483 => "0000000011011011000001",
			3484 => "0000000011011011000001",
			3485 => "0001101000110100001000",
			3486 => "0000001011111100000100",
			3487 => "0000000011011011000001",
			3488 => "0000000011011011000001",
			3489 => "0011101100011000000100",
			3490 => "0000000011011011000001",
			3491 => "0000000011011011000001",
			3492 => "0000001010111000000100",
			3493 => "0000000011011011000001",
			3494 => "0000000011011011000001",
			3495 => "0010101001011000000100",
			3496 => "0000000011011011000001",
			3497 => "0011000101011100000100",
			3498 => "0000000011011011000001",
			3499 => "0010101100110100000100",
			3500 => "0000000011011011000001",
			3501 => "0000111010011100000100",
			3502 => "0000000011011011000001",
			3503 => "0000000011011011000001",
			3504 => "0011001110011000011000",
			3505 => "0001100101001100001100",
			3506 => "0010001010100100000100",
			3507 => "0000000011011101101101",
			3508 => "0011011011101100000100",
			3509 => "1111111011011101101101",
			3510 => "0000000011011101101101",
			3511 => "0010010101011100001000",
			3512 => "0010001111111100000100",
			3513 => "0000001011011101101101",
			3514 => "0000000011011101101101",
			3515 => "0000000011011101101101",
			3516 => "0011100110110000110100",
			3517 => "0000010110010000011100",
			3518 => "0011101111110000001100",
			3519 => "0001001100001100000100",
			3520 => "1111111011011101101101",
			3521 => "0010001111111100000100",
			3522 => "0000000011011101101101",
			3523 => "0000000011011101101101",
			3524 => "0011111000001000001100",
			3525 => "0001011000000000000100",
			3526 => "0000000011011101101101",
			3527 => "0000101011010000000100",
			3528 => "0000000011011101101101",
			3529 => "0000001011011101101101",
			3530 => "0000000011011101101101",
			3531 => "0001011111101000001000",
			3532 => "0011111011110100000100",
			3533 => "1111111011011101101101",
			3534 => "0000000011011101101101",
			3535 => "0011010011010000001100",
			3536 => "0001000011000100001000",
			3537 => "0000000100110000000100",
			3538 => "0000000011011101101101",
			3539 => "0000001011011101101101",
			3540 => "0000000011011101101101",
			3541 => "0000000011011101101101",
			3542 => "0000010110010000000100",
			3543 => "1111111011011101101101",
			3544 => "0010011001001000000100",
			3545 => "0000000011011101101101",
			3546 => "0000000011011101101101",
			3547 => "0011001110011000011100",
			3548 => "0011101101100000010000",
			3549 => "0001001010000100001100",
			3550 => "0010001010100100000100",
			3551 => "0000000011100000101001",
			3552 => "0000010111100100000100",
			3553 => "0000000011100000101001",
			3554 => "0000000011100000101001",
			3555 => "0000000011100000101001",
			3556 => "0000001110101000001000",
			3557 => "0010001111111100000100",
			3558 => "0000000011100000101001",
			3559 => "0000000011100000101001",
			3560 => "0000000011100000101001",
			3561 => "0000011000011000110000",
			3562 => "0000001101110100010100",
			3563 => "0000110011000100000100",
			3564 => "0000000011100000101001",
			3565 => "0001110110101100001100",
			3566 => "0010011101101000000100",
			3567 => "0000000011100000101001",
			3568 => "0010110101010100000100",
			3569 => "0000000011100000101001",
			3570 => "0000000011100000101001",
			3571 => "0000000011100000101001",
			3572 => "0001100101001100001100",
			3573 => "0010000101101100001000",
			3574 => "0001111101001000000100",
			3575 => "0000000011100000101001",
			3576 => "0000000011100000101001",
			3577 => "0000000011100000101001",
			3578 => "0000001110110000001000",
			3579 => "0000001011001100000100",
			3580 => "0000000011100000101001",
			3581 => "0000000011100000101001",
			3582 => "0011101101100100000100",
			3583 => "0000000011100000101001",
			3584 => "0000000011100000101001",
			3585 => "0010101100110100001100",
			3586 => "0001111111101000000100",
			3587 => "0000000011100000101001",
			3588 => "0001110100101100000100",
			3589 => "0000000011100000101001",
			3590 => "0000000011100000101001",
			3591 => "0001111111101000000100",
			3592 => "0000000011100000101001",
			3593 => "0000000011100000101001",
			3594 => "0001011101001000100100",
			3595 => "0000100111111000011100",
			3596 => "0011010011110000000100",
			3597 => "0000000011100011100101",
			3598 => "0000111000000000001100",
			3599 => "0000111111011000001000",
			3600 => "0000110011000000000100",
			3601 => "0000000011100011100101",
			3602 => "0000000011100011100101",
			3603 => "0000000011100011100101",
			3604 => "0001001100101000000100",
			3605 => "0000000011100011100101",
			3606 => "0011100011101100000100",
			3607 => "0000000011100011100101",
			3608 => "0000000011100011100101",
			3609 => "0011110100110100000100",
			3610 => "0000000011100011100101",
			3611 => "0000000011100011100101",
			3612 => "0001011011000000010100",
			3613 => "0011100110110000001100",
			3614 => "0010011001000100001000",
			3615 => "0000000111101100000100",
			3616 => "0000000011100011100101",
			3617 => "0000000011100011100101",
			3618 => "0000000011100011100101",
			3619 => "0000000101010000000100",
			3620 => "0000000011100011100101",
			3621 => "0000000011100011100101",
			3622 => "0000110000111100011100",
			3623 => "0000100111000100001100",
			3624 => "0011100010001100001000",
			3625 => "0001101010100000000100",
			3626 => "0000000011100011100101",
			3627 => "0000000011100011100101",
			3628 => "0000000011100011100101",
			3629 => "0010000101101100000100",
			3630 => "0000000011100011100101",
			3631 => "0010100000111100000100",
			3632 => "0000000011100011100101",
			3633 => "0000111100101100000100",
			3634 => "0000000011100011100101",
			3635 => "0000000011100011100101",
			3636 => "0001011001101100001000",
			3637 => "0011111001011100000100",
			3638 => "0000000011100011100101",
			3639 => "0000000011100011100101",
			3640 => "0000000011100011100101",
			3641 => "0011001100101000110100",
			3642 => "0001100101001000010000",
			3643 => "0010000101101100000100",
			3644 => "1111111011100101010001",
			3645 => "0011011011101100001000",
			3646 => "0001000101010100000100",
			3647 => "1111111011100101010001",
			3648 => "0000010011100101010001",
			3649 => "1111111011100101010001",
			3650 => "0011100001000000100000",
			3651 => "0000110011001000001100",
			3652 => "0011010110110100001000",
			3653 => "0001111100110000000100",
			3654 => "1111111011100101010001",
			3655 => "0000001011100101010001",
			3656 => "1111111011100101010001",
			3657 => "0000010001100100010000",
			3658 => "0010101011111000001000",
			3659 => "0000000101101000000100",
			3660 => "0000000011100101010001",
			3661 => "0000001011100101010001",
			3662 => "0001011001101100000100",
			3663 => "0000001011100101010001",
			3664 => "1111111011100101010001",
			3665 => "1111111011100101010001",
			3666 => "1111111011100101010001",
			3667 => "1111111011100101010001",
			3668 => "0000011000011000110100",
			3669 => "0000011000111100001000",
			3670 => "0011010110110100000100",
			3671 => "1111111011100111001101",
			3672 => "0000000011100111001101",
			3673 => "0001011000000100000100",
			3674 => "1111111011100111001101",
			3675 => "0010111110011000001100",
			3676 => "0001100100011100000100",
			3677 => "1111111011100111001101",
			3678 => "0010001111111100000100",
			3679 => "0000001011100111001101",
			3680 => "0000000011100111001101",
			3681 => "0011101111110100010000",
			3682 => "0000100111110100001000",
			3683 => "0011100100100100000100",
			3684 => "0000000011100111001101",
			3685 => "1111111011100111001101",
			3686 => "0001101000101100000100",
			3687 => "0000001011100111001101",
			3688 => "0000001011100111001101",
			3689 => "0011101101100000000100",
			3690 => "1111111011100111001101",
			3691 => "0011100110110000000100",
			3692 => "0000000011100111001101",
			3693 => "0000000011100111001101",
			3694 => "0001111111101000000100",
			3695 => "1111111011100111001101",
			3696 => "0001110100101100000100",
			3697 => "0000001011100111001101",
			3698 => "1111111011100111001101",
			3699 => "0000110011100100011100",
			3700 => "0001100000001100010100",
			3701 => "0001011001010100010000",
			3702 => "0000111111011000001100",
			3703 => "0011100001101100001000",
			3704 => "0000110011000000000100",
			3705 => "0000000011101010000001",
			3706 => "0000000011101010000001",
			3707 => "0000000011101010000001",
			3708 => "0000000011101010000001",
			3709 => "0000000011101010000001",
			3710 => "0001000101010100000100",
			3711 => "0000000011101010000001",
			3712 => "0000000011101010000001",
			3713 => "0010010101101100100000",
			3714 => "0011001110011000001100",
			3715 => "0011101101100000000100",
			3716 => "0000000011101010000001",
			3717 => "0010001111111100000100",
			3718 => "0000000011101010000001",
			3719 => "0000000011101010000001",
			3720 => "0000011000011000010000",
			3721 => "0011101111110000000100",
			3722 => "0000000011101010000001",
			3723 => "0011101111010100000100",
			3724 => "0000000011101010000001",
			3725 => "0001101101010000000100",
			3726 => "0000000011101010000001",
			3727 => "0000000011101010000001",
			3728 => "0000000011101010000001",
			3729 => "0010101001011000000100",
			3730 => "0000000011101010000001",
			3731 => "0010110101010100010000",
			3732 => "0001001100101100000100",
			3733 => "0000000011101010000001",
			3734 => "0000110000111100000100",
			3735 => "0000000011101010000001",
			3736 => "0001011001101100000100",
			3737 => "0000000011101010000001",
			3738 => "0000000011101010000001",
			3739 => "0010101100110100000100",
			3740 => "0000000011101010000001",
			3741 => "0001011001101100000100",
			3742 => "0000000011101010000001",
			3743 => "0000000011101010000001",
			3744 => "0011001110011000010100",
			3745 => "0001100101001100001100",
			3746 => "0010001010100100000100",
			3747 => "0000000011101100100101",
			3748 => "0011011011101100000100",
			3749 => "1111111011101100100101",
			3750 => "0000000011101100100101",
			3751 => "0000010111110000000100",
			3752 => "0000001011101100100101",
			3753 => "0000000011101100100101",
			3754 => "0010000011010000001000",
			3755 => "0011100010011000000100",
			3756 => "0000000011101100100101",
			3757 => "0000001011101100100101",
			3758 => "0000110011100100010000",
			3759 => "0011100001101100001000",
			3760 => "0010101100010000000100",
			3761 => "0000000011101100100101",
			3762 => "0000000011101100100101",
			3763 => "0000001001101000000100",
			3764 => "1111111011101100100101",
			3765 => "0000000011101100100101",
			3766 => "0010010101101100010000",
			3767 => "0000011000011000001100",
			3768 => "0010000101101100001000",
			3769 => "0000001011111100000100",
			3770 => "0000000011101100100101",
			3771 => "0000001011101100100101",
			3772 => "0000000011101100100101",
			3773 => "0000000011101100100101",
			3774 => "0010101001011000001100",
			3775 => "0000000101010000000100",
			3776 => "1111111011101100100101",
			3777 => "0000001001101000000100",
			3778 => "0000000011101100100101",
			3779 => "0000000011101100100101",
			3780 => "0011010110001100000100",
			3781 => "0000000011101100100101",
			3782 => "0010010011000000000100",
			3783 => "0000000011101100100101",
			3784 => "0000000011101100100101",
			3785 => "0011100110110001001000",
			3786 => "0011011011101100101000",
			3787 => "0011101101100000100000",
			3788 => "0001011101001000010000",
			3789 => "0010101101001000001100",
			3790 => "0001100001100000001000",
			3791 => "0010010101011100000100",
			3792 => "0000000011101111011001",
			3793 => "0000000011101111011001",
			3794 => "0000000011101111011001",
			3795 => "0000000011101111011001",
			3796 => "0000001011100100001100",
			3797 => "0010001111111100001000",
			3798 => "0000110000111100000100",
			3799 => "0000000011101111011001",
			3800 => "0000000011101111011001",
			3801 => "0000000011101111011001",
			3802 => "0000000011101111011001",
			3803 => "0000010110010000000100",
			3804 => "0000000011101111011001",
			3805 => "0000000011101111011001",
			3806 => "0010001001001100001000",
			3807 => "0001100101001000000100",
			3808 => "0000000011101111011001",
			3809 => "0000000011101111011001",
			3810 => "0000111101001000000100",
			3811 => "0000000011101111011001",
			3812 => "0001011011000000001000",
			3813 => "0000001011111100000100",
			3814 => "0000000011101111011001",
			3815 => "0000000011101111011001",
			3816 => "0010101100110100000100",
			3817 => "0000000011101111011001",
			3818 => "0000111010011100000100",
			3819 => "0000000011101111011001",
			3820 => "0000000011101111011001",
			3821 => "0010111011101100001000",
			3822 => "0011110011111100000100",
			3823 => "0000000011101111011001",
			3824 => "0000000011101111011001",
			3825 => "0000010110010000000100",
			3826 => "0000000011101111011001",
			3827 => "0000011000011000000100",
			3828 => "0000000011101111011001",
			3829 => "0000000011101111011001",
			3830 => "0011100001000000110000",
			3831 => "0000100111111000101000",
			3832 => "0000100110100100100100",
			3833 => "0000001101110000011100",
			3834 => "0011100010110000010000",
			3835 => "0010101001000000001000",
			3836 => "0001000101011100000100",
			3837 => "0000000011110000111101",
			3838 => "0000000011110000111101",
			3839 => "0001000011000100000100",
			3840 => "0000000011110000111101",
			3841 => "0000000011110000111101",
			3842 => "0000100110101000001000",
			3843 => "0000010001100100000100",
			3844 => "0000000011110000111101",
			3845 => "0000000011110000111101",
			3846 => "0000000011110000111101",
			3847 => "0000010110010000000100",
			3848 => "0000000011110000111101",
			3849 => "0000000011110000111101",
			3850 => "0000000011110000111101",
			3851 => "0010000101101100000100",
			3852 => "0000000011110000111101",
			3853 => "0000000011110000111101",
			3854 => "0000000011110000111101",
			3855 => "0011010011010001000000",
			3856 => "0000110011001000001100",
			3857 => "0011010110110100001000",
			3858 => "0001000101010100000100",
			3859 => "1111111011110011000001",
			3860 => "0000001011110011000001",
			3861 => "1111111011110011000001",
			3862 => "0011100110110000100100",
			3863 => "0011111001011100001100",
			3864 => "0011100010001100001000",
			3865 => "0000001110010000000100",
			3866 => "1111111011110011000001",
			3867 => "0000001011110011000001",
			3868 => "1111111011110011000001",
			3869 => "0010101001011000001100",
			3870 => "0010000101101100001000",
			3871 => "0000000101101000000100",
			3872 => "0000000011110011000001",
			3873 => "0000001011110011000001",
			3874 => "1111111011110011000001",
			3875 => "0001011001101100001000",
			3876 => "0011010110001100000100",
			3877 => "0000000011110011000001",
			3878 => "0000001011110011000001",
			3879 => "1111111011110011000001",
			3880 => "0010111110011000001000",
			3881 => "0000001111001100000100",
			3882 => "1111111011110011000001",
			3883 => "0000001011110011000001",
			3884 => "0000001010111000000100",
			3885 => "1111111011110011000001",
			3886 => "0000000011110011000001",
			3887 => "1111111011110011000001",
			3888 => "0001011101001000101000",
			3889 => "0000110011100100011000",
			3890 => "0000100111111000010100",
			3891 => "0000111111011000010000",
			3892 => "0011010110110100001100",
			3893 => "0011011101000000000100",
			3894 => "0000000011110110000101",
			3895 => "0001001011101100000100",
			3896 => "0000000011110110000101",
			3897 => "0000000011110110000101",
			3898 => "0000000011110110000101",
			3899 => "1111111011110110000101",
			3900 => "0000000011110110000101",
			3901 => "0000000110111100000100",
			3902 => "1111111011110110000101",
			3903 => "0001111101001000000100",
			3904 => "0000001011110110000101",
			3905 => "0000010110010000000100",
			3906 => "0000000011110110000101",
			3907 => "0000000011110110000101",
			3908 => "0011100110110000110000",
			3909 => "0011101010011000010000",
			3910 => "0000001101010000001100",
			3911 => "0000110011000100000100",
			3912 => "0000000011110110000101",
			3913 => "0010101110111000000100",
			3914 => "0000001011110110000101",
			3915 => "0000000011110110000101",
			3916 => "1111111011110110000101",
			3917 => "0010000101101100010000",
			3918 => "0011011010100100001100",
			3919 => "0001011001101100001000",
			3920 => "0001111100110000000100",
			3921 => "0000000011110110000101",
			3922 => "0000001011110110000101",
			3923 => "0000000011110110000101",
			3924 => "0000000011110110000101",
			3925 => "0010101001011000000100",
			3926 => "1111111011110110000101",
			3927 => "0010001111001000001000",
			3928 => "0001001100001100000100",
			3929 => "0000001011110110000101",
			3930 => "0000000011110110000101",
			3931 => "0000000011110110000101",
			3932 => "0000101111001100000100",
			3933 => "1111111011110110000101",
			3934 => "0000100101101000000100",
			3935 => "0000000011110110000101",
			3936 => "0000000011110110000101",
			3937 => "0000110000111100111100",
			3938 => "0010010110000000111000",
			3939 => "0011001110011000010100",
			3940 => "0001100101001100001100",
			3941 => "0001001010000100001000",
			3942 => "0010001010100100000100",
			3943 => "0000000011111000011001",
			3944 => "1111111011111000011001",
			3945 => "0000001011111000011001",
			3946 => "0000010111110000000100",
			3947 => "0000001011111000011001",
			3948 => "0000000011111000011001",
			3949 => "0011100110110000010100",
			3950 => "0000001011111100000100",
			3951 => "1111111011111000011001",
			3952 => "0000110011100100001000",
			3953 => "0011010110001100000100",
			3954 => "0000000011111000011001",
			3955 => "1111111011111000011001",
			3956 => "0010000101101100000100",
			3957 => "0000001011111000011001",
			3958 => "0000000011111000011001",
			3959 => "0000010110010000000100",
			3960 => "1111111011111000011001",
			3961 => "0001101010110000001000",
			3962 => "0010101001010100000100",
			3963 => "0000000011111000011001",
			3964 => "0000000011111000011001",
			3965 => "0000000011111000011001",
			3966 => "1111111011111000011001",
			3967 => "0001011001101100001100",
			3968 => "0011111001011100000100",
			3969 => "0000000011111000011001",
			3970 => "0010011000000100000100",
			3971 => "0000001011111000011001",
			3972 => "0000000011111000011001",
			3973 => "0000000011111000011001",
			3974 => "0000001101110001000000",
			3975 => "0001010001010000011000",
			3976 => "0011000111011100001100",
			3977 => "0011100111001000000100",
			3978 => "1111111011111011110101",
			3979 => "0000111101001000000100",
			3980 => "0000000011111011110101",
			3981 => "0000000011111011110101",
			3982 => "0001111100110000001000",
			3983 => "0001111100010000000100",
			3984 => "0000000011111011110101",
			3985 => "0000000011111011110101",
			3986 => "0000000011111011110101",
			3987 => "0001011011000000001100",
			3988 => "0010101000101000000100",
			3989 => "0000000011111011110101",
			3990 => "0000010001100100000100",
			3991 => "0000000011111011110101",
			3992 => "0000000011111011110101",
			3993 => "0010101100001100010100",
			3994 => "0011100010001100001000",
			3995 => "0011111101101100000100",
			3996 => "0000000011111011110101",
			3997 => "0000000011111011110101",
			3998 => "0010001001001100000100",
			3999 => "0000000011111011110101",
			4000 => "0000000010101100000100",
			4001 => "1111111011111011110101",
			4002 => "0000000011111011110101",
			4003 => "0001011001101100000100",
			4004 => "0000000011111011110101",
			4005 => "0000000011111011110101",
			4006 => "0011100011011000000100",
			4007 => "0000000011111011110101",
			4008 => "0000111100010000010000",
			4009 => "0001100100100000001000",
			4010 => "0000100111111000000100",
			4011 => "1111111011111011110101",
			4012 => "0000000011111011110101",
			4013 => "0001101010110000000100",
			4014 => "0000000011111011110101",
			4015 => "0000000011111011110101",
			4016 => "0010001111111100001000",
			4017 => "0010001001001100000100",
			4018 => "0000000011111011110101",
			4019 => "0000000011111011110101",
			4020 => "0001011000100000001100",
			4021 => "0000101111001100000100",
			4022 => "0000000011111011110101",
			4023 => "0000001000001100000100",
			4024 => "0000000011111011110101",
			4025 => "0000000011111011110101",
			4026 => "0011001001001000000100",
			4027 => "0000000011111011110101",
			4028 => "0000000011111011110101",
			4029 => "0001110110101100110000",
			4030 => "0000111000000000010000",
			4031 => "0001001001000100000100",
			4032 => "1111111011111111000001",
			4033 => "0000010001110000000100",
			4034 => "0000000011111111000001",
			4035 => "0001000110000000000100",
			4036 => "0000000011111111000001",
			4037 => "0000000011111111000001",
			4038 => "0000011000011000011100",
			4039 => "0001111100010000010000",
			4040 => "0001111100000000001000",
			4041 => "0000000100110000000100",
			4042 => "0000000011111111000001",
			4043 => "0000000011111111000001",
			4044 => "0001001001010000000100",
			4045 => "0000000011111111000001",
			4046 => "0000000011111111000001",
			4047 => "0001100101001000000100",
			4048 => "0000000011111111000001",
			4049 => "0000001101110100000100",
			4050 => "0000000011111111000001",
			4051 => "0000001011111111000001",
			4052 => "0000000011111111000001",
			4053 => "0000101101110000101100",
			4054 => "0010010101011100001000",
			4055 => "0011111010110000000100",
			4056 => "0000000011111111000001",
			4057 => "1111111011111111000001",
			4058 => "0010001001001100001000",
			4059 => "0000001000010000000100",
			4060 => "0000000011111111000001",
			4061 => "0000000011111111000001",
			4062 => "0010101001010100001100",
			4063 => "0011100011010100001000",
			4064 => "0001111101001000000100",
			4065 => "0000000011111111000001",
			4066 => "0000000011111111000001",
			4067 => "1111111011111111000001",
			4068 => "0010011001000100001000",
			4069 => "0000000011001100000100",
			4070 => "0000000011111111000001",
			4071 => "0000000011111111000001",
			4072 => "0010101100110100000100",
			4073 => "0000000011111111000001",
			4074 => "0000000011111111000001",
			4075 => "0011100001000000001000",
			4076 => "0010000101101100000100",
			4077 => "0000000011111111000001",
			4078 => "0000000011111111000001",
			4079 => "0000000011111111000001",
			4080 => "0001010001111101001000",
			4081 => "0000011001100100010100",
			4082 => "0011001110011000000100",
			4083 => "1111111100000001011101",
			4084 => "0010011001001000001000",
			4085 => "0000111111011000000100",
			4086 => "0000000100000001011101",
			4087 => "0000001100000001011101",
			4088 => "0011011011101100000100",
			4089 => "1111111100000001011101",
			4090 => "0000000100000001011101",
			4091 => "0011011010100100100100",
			4092 => "0000011000011000100000",
			4093 => "0010101101001000010000",
			4094 => "0011001110011000001000",
			4095 => "0011001011101100000100",
			4096 => "0000000100000001011101",
			4097 => "1111111100000001011101",
			4098 => "0000000110111100000100",
			4099 => "0000000100000001011101",
			4100 => "0000000100000001011101",
			4101 => "0011001010100100001000",
			4102 => "0001011000000000000100",
			4103 => "0000000100000001011101",
			4104 => "0000001100000001011101",
			4105 => "0011100110110000000100",
			4106 => "0000000100000001011101",
			4107 => "1111111100000001011101",
			4108 => "1111111100000001011101",
			4109 => "0011101111010100001000",
			4110 => "0010111010100100000100",
			4111 => "0000000100000001011101",
			4112 => "1111111100000001011101",
			4113 => "0011111110000100000100",
			4114 => "0000000100000001011101",
			4115 => "0000000100000001011101",
			4116 => "0001011001101100000100",
			4117 => "0000001100000001011101",
			4118 => "0000000100000001011101",
			4119 => "0000011000011001001100",
			4120 => "0011011010100101000100",
			4121 => "0000011001100100011000",
			4122 => "0010001111111100010000",
			4123 => "0011011011101100001100",
			4124 => "0011110101111100001000",
			4125 => "0010101001011000000100",
			4126 => "0000000100000100011001",
			4127 => "0000000100000100011001",
			4128 => "0000000100000100011001",
			4129 => "0000000100000100011001",
			4130 => "0001111100010000000100",
			4131 => "0000000100000100011001",
			4132 => "0000000100000100011001",
			4133 => "0010000101011100010100",
			4134 => "0001011000000000001000",
			4135 => "0001111001010000000100",
			4136 => "0000000100000100011001",
			4137 => "0000000100000100011001",
			4138 => "0001000110011100001000",
			4139 => "0011101010110100000100",
			4140 => "0000000100000100011001",
			4141 => "0000000100000100011001",
			4142 => "0000000100000100011001",
			4143 => "0001011111101000001100",
			4144 => "0000001110110000001000",
			4145 => "0001100000010000000100",
			4146 => "0000000100000100011001",
			4147 => "0000000100000100011001",
			4148 => "0000000100000100011001",
			4149 => "0001001100101100001000",
			4150 => "0010000101101100000100",
			4151 => "0000000100000100011001",
			4152 => "0000000100000100011001",
			4153 => "0000000100000100011001",
			4154 => "0011000111011100000100",
			4155 => "0000000100000100011001",
			4156 => "0000000100000100011001",
			4157 => "0001001001011000001100",
			4158 => "0001111111101000000100",
			4159 => "0000000100000100011001",
			4160 => "0001110100101100000100",
			4161 => "0000000100000100011001",
			4162 => "0000000100000100011001",
			4163 => "0001010001011100000100",
			4164 => "0000000100000100011001",
			4165 => "0000000100000100011001",
			4166 => "0000010001100100110000",
			4167 => "0001011000000100000100",
			4168 => "1111111100000101111101",
			4169 => "0010001010100100000100",
			4170 => "0000001100000101111101",
			4171 => "0010101001011000010100",
			4172 => "0010000101101100010000",
			4173 => "0000101101110000001000",
			4174 => "0011111101001100000100",
			4175 => "0000000100000101111101",
			4176 => "1111111100000101111101",
			4177 => "0001100000001100000100",
			4178 => "0000001100000101111101",
			4179 => "0000000100000101111101",
			4180 => "1111111100000101111101",
			4181 => "0000100111000100001100",
			4182 => "0011110001101100001000",
			4183 => "0010011101101000000100",
			4184 => "1111111100000101111101",
			4185 => "0000001100000101111101",
			4186 => "1111111100000101111101",
			4187 => "0001100111101000000100",
			4188 => "0000001100000101111101",
			4189 => "0000000100000101111101",
			4190 => "1111111100000101111101",
			4191 => "0011100110110001001100",
			4192 => "0001100000010001001000",
			4193 => "0001010110101100011000",
			4194 => "0000111000000000010000",
			4195 => "0011010110110100001100",
			4196 => "0011011111011100000100",
			4197 => "0000000100001000111001",
			4198 => "0011101001011100000100",
			4199 => "0000000100001000111001",
			4200 => "0000000100001000111001",
			4201 => "0000000100001000111001",
			4202 => "0010001111111100000100",
			4203 => "0000000100001000111001",
			4204 => "0000000100001000111001",
			4205 => "0000010111100100011000",
			4206 => "0011110101111100010000",
			4207 => "0011010110001100001000",
			4208 => "0011010110110100000100",
			4209 => "0000000100001000111001",
			4210 => "0000000100001000111001",
			4211 => "0011011010100100000100",
			4212 => "0000000100001000111001",
			4213 => "0000000100001000111001",
			4214 => "0000010001110000000100",
			4215 => "0000000100001000111001",
			4216 => "0000000100001000111001",
			4217 => "0000111011111000001100",
			4218 => "0001011001010000000100",
			4219 => "0000000100001000111001",
			4220 => "0001011000100000000100",
			4221 => "0000000100001000111001",
			4222 => "0000000100001000111001",
			4223 => "0011100101001000000100",
			4224 => "0000000100001000111001",
			4225 => "0011010011010000000100",
			4226 => "0000000100001000111001",
			4227 => "0000000100001000111001",
			4228 => "0000000100001000111001",
			4229 => "0010111011101100001000",
			4230 => "0011110111001100000100",
			4231 => "0000000100001000111001",
			4232 => "0000000100001000111001",
			4233 => "0000010110010000000100",
			4234 => "0000000100001000111001",
			4235 => "0000011000011000000100",
			4236 => "0000000100001000111001",
			4237 => "0000000100001000111001",
			4238 => "0000011001100100011100",
			4239 => "0011001110011000000100",
			4240 => "1111111100001100110111",
			4241 => "0010011001001000001000",
			4242 => "0001010110101100000100",
			4243 => "0000000100001100110111",
			4244 => "0000001100001100110111",
			4245 => "0011011011101100001000",
			4246 => "0010001001001100000100",
			4247 => "0000000100001100110111",
			4248 => "1111111100001100110111",
			4249 => "0001001001010000000100",
			4250 => "0000000100001100110111",
			4251 => "0000000100001100110111",
			4252 => "0010000101011100101000",
			4253 => "0000011000011000100100",
			4254 => "0001001001000100010000",
			4255 => "0001001100101000001100",
			4256 => "0001000101010100001000",
			4257 => "0011011011101100000100",
			4258 => "0000000100001100110111",
			4259 => "0000000100001100110111",
			4260 => "0000001100001100110111",
			4261 => "0000000100001100110111",
			4262 => "0001000110011100010000",
			4263 => "0000101011100100001000",
			4264 => "0000001001110100000100",
			4265 => "0000000100001100110111",
			4266 => "0000001100001100110111",
			4267 => "0001101010101100000100",
			4268 => "0000001100001100110111",
			4269 => "0000000100001100110111",
			4270 => "0000000100001100110111",
			4271 => "1111111100001100110111",
			4272 => "0000111101001000010000",
			4273 => "0000001001101000001000",
			4274 => "0010100100101100000100",
			4275 => "1111111100001100110111",
			4276 => "0000000100001100110111",
			4277 => "0000001101011000000100",
			4278 => "0000001100001100110111",
			4279 => "1111111100001100110111",
			4280 => "0001011011000000010000",
			4281 => "0010101000101000000100",
			4282 => "0000000100001100110111",
			4283 => "0010011001000100001000",
			4284 => "0001101101010100000100",
			4285 => "0000001100001100110111",
			4286 => "0000000100001100110111",
			4287 => "0000000100001100110111",
			4288 => "0010101001000000001100",
			4289 => "0001001111011000000100",
			4290 => "0000000100001100110111",
			4291 => "0001111001010100000100",
			4292 => "1111111100001100110111",
			4293 => "0000000100001100110111",
			4294 => "0001011110010100001000",
			4295 => "0001011100110100000100",
			4296 => "0000000100001100110111",
			4297 => "0000001100001100110111",
			4298 => "0010101100110100000100",
			4299 => "1111111100001100110111",
			4300 => "0000001100001100110111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1489, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2851, initial_addr_3'length));
	end generate gen_rom_2;

	gen_rom_3: if SELECT_ROM = 3 generate
		bank <= (
			0 => "0011011100101000100000",
			1 => "0010011110011000000100",
			2 => "0000001000000001010101",
			3 => "0010101111011000001000",
			4 => "0010001010100100000100",
			5 => "0000000000000001010101",
			6 => "1111111000000001010101",
			7 => "0010100011001000000100",
			8 => "0000001000000001010101",
			9 => "0001001011111000001100",
			10 => "0001001001010000001000",
			11 => "0010110101010100000100",
			12 => "0000000000000001010101",
			13 => "0000000000000001010101",
			14 => "0000001000000001010101",
			15 => "1111111000000001010101",
			16 => "0000010001100100001000",
			17 => "0000000111101100000100",
			18 => "0000000000000001010101",
			19 => "0000001000000001010101",
			20 => "1111111000000001010101",
			21 => "0011111101100100010100",
			22 => "0001000111110000001000",
			23 => "0001101011000000000100",
			24 => "1111111000000010111001",
			25 => "0000100000000010111001",
			26 => "0011000111011100001000",
			27 => "0010110011010000000100",
			28 => "1111111000000010111001",
			29 => "0000001000000010111001",
			30 => "1111111000000010111001",
			31 => "0010011111011000011100",
			32 => "0000111011000000011000",
			33 => "0011101001011100000100",
			34 => "0000001000000010111001",
			35 => "0000110011000000001000",
			36 => "0000001101011100000100",
			37 => "1111111000000010111001",
			38 => "0000000000000010111001",
			39 => "0000101011101000000100",
			40 => "1111111000000010111001",
			41 => "0011100100011100000100",
			42 => "0000000000000010111001",
			43 => "1111111000000010111001",
			44 => "0000000000000010111001",
			45 => "1111111000000010111001",
			46 => "0000100111110100011000",
			47 => "0011111101100100010000",
			48 => "0010011010100100000100",
			49 => "0000000000000100101101",
			50 => "0011000111011100001000",
			51 => "0010110111011100000100",
			52 => "1111111000000100101101",
			53 => "0000001000000100101101",
			54 => "1111111000000100101101",
			55 => "0001110110101100000100",
			56 => "0000001000000100101101",
			57 => "1111111000000100101101",
			58 => "0010011111011000100000",
			59 => "0011100100011100011100",
			60 => "0011000101011100010100",
			61 => "0011010101010100010000",
			62 => "0001111101001000001000",
			63 => "0001011101001000000100",
			64 => "0000001000000100101101",
			65 => "1111111000000100101101",
			66 => "0000010001110000000100",
			67 => "0000010000000100101101",
			68 => "0000001000000100101101",
			69 => "0000000000000100101101",
			70 => "0010101011111000000100",
			71 => "0000001000000100101101",
			72 => "0000010000000100101101",
			73 => "1111111000000100101101",
			74 => "1111111000000100101101",
			75 => "0001001100000000101100",
			76 => "0001001000000100101000",
			77 => "0010000000110000011000",
			78 => "0010101011000000010100",
			79 => "0001010100101100010000",
			80 => "0011000101010100001000",
			81 => "0001000011010000000100",
			82 => "0000000000000110111001",
			83 => "0000000000000110111001",
			84 => "0001001100101000000100",
			85 => "1111111000000110111001",
			86 => "0000000000000110111001",
			87 => "0000000000000110111001",
			88 => "0000001000000110111001",
			89 => "0001001001001000001100",
			90 => "0001111111101000000100",
			91 => "0000000000000110111001",
			92 => "0001111011111000000100",
			93 => "0000000000000110111001",
			94 => "0000000000000110111001",
			95 => "1111111000000110111001",
			96 => "0000001000000110111001",
			97 => "0001001001010000001100",
			98 => "0010110101010100000100",
			99 => "1111111000000110111001",
			100 => "0010111100101000000100",
			101 => "0000000000000110111001",
			102 => "1111111000000110111001",
			103 => "0001000100101100001100",
			104 => "0011110001100000000100",
			105 => "0000000000000110111001",
			106 => "0000111011000000000100",
			107 => "0000001000000110111001",
			108 => "0000000000000110111001",
			109 => "0000000000000110111001",
			110 => "0000001001110100011100",
			111 => "0011010111011100010000",
			112 => "0010011101101000000100",
			113 => "0000000000001001011101",
			114 => "0000111001010100000100",
			115 => "0000000000001001011101",
			116 => "0001011100110100000100",
			117 => "0000000000001001011101",
			118 => "0000000000001001011101",
			119 => "0001011000111000001000",
			120 => "0010010110000000000100",
			121 => "0000000000001001011101",
			122 => "0000000000001001011101",
			123 => "0000000000001001011101",
			124 => "0001100101000000001000",
			125 => "0000011000011000000100",
			126 => "0000000000001001011101",
			127 => "0000000000001001011101",
			128 => "0000100110010100001100",
			129 => "0000100011111000000100",
			130 => "0000000000001001011101",
			131 => "0011001110011000000100",
			132 => "0000000000001001011101",
			133 => "0000000000001001011101",
			134 => "0001101010111100010000",
			135 => "0000000101101000001100",
			136 => "0001110110101100000100",
			137 => "0000000000001001011101",
			138 => "0001010011000100000100",
			139 => "0000000000001001011101",
			140 => "0000000000001001011101",
			141 => "0000000000001001011101",
			142 => "0000010001110000000100",
			143 => "0000000000001001011101",
			144 => "0000001010111000001000",
			145 => "0001011100101100000100",
			146 => "0000000000001001011101",
			147 => "0000000000001001011101",
			148 => "0001110100101100000100",
			149 => "0000000000001001011101",
			150 => "0000000000001001011101",
			151 => "0001000111110000001000",
			152 => "0011101011111000000100",
			153 => "0000000000001010111001",
			154 => "0000011000001010111001",
			155 => "0011100010001100000100",
			156 => "1111111000001010111001",
			157 => "0000000100111000000100",
			158 => "0000001000001010111001",
			159 => "0011111101100100000100",
			160 => "1111111000001010111001",
			161 => "0011111100111100010000",
			162 => "0011011011101100001000",
			163 => "0000010110010000000100",
			164 => "0000000000001010111001",
			165 => "0000001000001010111001",
			166 => "0011000011010000000100",
			167 => "1111111000001010111001",
			168 => "0000000000001010111001",
			169 => "0000001010010100000100",
			170 => "1111111000001010111001",
			171 => "0011010101010100000100",
			172 => "0000000000001010111001",
			173 => "0000000000001010111001",
			174 => "0001001100000000110000",
			175 => "0001001000000100101100",
			176 => "0001001111011000100100",
			177 => "0000011000111100010000",
			178 => "0001110110101100001100",
			179 => "0011010110110100001000",
			180 => "0010010111011100000100",
			181 => "0000000000001101010101",
			182 => "0000000000001101010101",
			183 => "0000000000001101010101",
			184 => "0000000000001101010101",
			185 => "0010101011000000010000",
			186 => "0010100100101100001000",
			187 => "0000001010111000000100",
			188 => "0000000000001101010101",
			189 => "0000000000001101010101",
			190 => "0011010111011100000100",
			191 => "1111111000001101010101",
			192 => "0000000000001101010101",
			193 => "0000000000001101010101",
			194 => "0010011101101000000100",
			195 => "0000000000001101010101",
			196 => "1111111000001101010101",
			197 => "0000001000001101010101",
			198 => "0001000110101100001100",
			199 => "0001011000100000000100",
			200 => "0000000000001101010101",
			201 => "0001010001001000000100",
			202 => "0000000000001101010101",
			203 => "0000000000001101010101",
			204 => "0001000100101100010000",
			205 => "0011000101010100000100",
			206 => "0000000000001101010101",
			207 => "0000101000011100000100",
			208 => "0000000000001101010101",
			209 => "0001110001001000000100",
			210 => "0000000000001101010101",
			211 => "0000000000001101010101",
			212 => "0000000000001101010101",
			213 => "0000001011111100011100",
			214 => "0011111101100100010000",
			215 => "0010011010100100000100",
			216 => "1101000000001111111001",
			217 => "0011000111011100001000",
			218 => "0011000011010000000100",
			219 => "1100111000001111111001",
			220 => "1100111000001111111001",
			221 => "1100111000001111111001",
			222 => "0001110110101100000100",
			223 => "1101011000001111111001",
			224 => "0000100111110100000100",
			225 => "1100111000001111111001",
			226 => "1101000000001111111001",
			227 => "0010010101111000110000",
			228 => "0011100110000100101100",
			229 => "0010011001000100011100",
			230 => "0010101000101000001100",
			231 => "0011100010001000000100",
			232 => "1110100000001111111001",
			233 => "0000110011000000000100",
			234 => "1100111000001111111001",
			235 => "1101101000001111111001",
			236 => "0001010001010000001000",
			237 => "0011110110011000000100",
			238 => "1101100000001111111001",
			239 => "1101000000001111111001",
			240 => "0000001001101000000100",
			241 => "1100111000001111111001",
			242 => "1101000000001111111001",
			243 => "0001110100101100001000",
			244 => "0011110111000000000100",
			245 => "1101110000001111111001",
			246 => "1110100000001111111001",
			247 => "0010101011000000000100",
			248 => "1101011000001111111001",
			249 => "1110001000001111111001",
			250 => "1100111000001111111001",
			251 => "0011010101011100000100",
			252 => "1101001000001111111001",
			253 => "1100111000001111111001",
			254 => "0011111101100100001100",
			255 => "0011000111011100001000",
			256 => "0010110111011100000100",
			257 => "1111111000010010000101",
			258 => "0000001000010010000101",
			259 => "1111111000010010000101",
			260 => "0010011111011000111000",
			261 => "0001100000001100100000",
			262 => "0011111000001000010100",
			263 => "0001101010111100010000",
			264 => "0000010110010000001000",
			265 => "0010010101011100000100",
			266 => "0000001000010010000101",
			267 => "1111111000010010000101",
			268 => "0000000110111100000100",
			269 => "0000000000010010000101",
			270 => "0000001000010010000101",
			271 => "1111111000010010000101",
			272 => "0011001010100100000100",
			273 => "1111111000010010000101",
			274 => "0000001110110000000100",
			275 => "0000010000010010000101",
			276 => "0000001000010010000101",
			277 => "0010111010100100001100",
			278 => "0001101110000100000100",
			279 => "1111111000010010000101",
			280 => "0011010110001100000100",
			281 => "0000001000010010000101",
			282 => "1111111000010010000101",
			283 => "0001111100101100000100",
			284 => "0000001000010010000101",
			285 => "0001011011111000000100",
			286 => "1111111000010010000101",
			287 => "0000000000010010000101",
			288 => "1111111000010010000101",
			289 => "0001101010101101001000",
			290 => "0011100011101100110000",
			291 => "0011100010110000101100",
			292 => "0000001011010000011100",
			293 => "0011001010100100001100",
			294 => "0000111101000000000100",
			295 => "0000000000010101010001",
			296 => "0001001010000100000100",
			297 => "0000000000010101010001",
			298 => "0000000000010101010001",
			299 => "0000011000011000001000",
			300 => "0000100100111100000100",
			301 => "0000000000010101010001",
			302 => "0000000000010101010001",
			303 => "0001011000000100000100",
			304 => "0000000000010101010001",
			305 => "0000000000010101010001",
			306 => "0001011100110000001000",
			307 => "0001100100000100000100",
			308 => "0000000000010101010001",
			309 => "0000000000010101010001",
			310 => "0000010110010000000100",
			311 => "0000000000010101010001",
			312 => "0000000000010101010001",
			313 => "0000000000010101010001",
			314 => "0000100110010100001100",
			315 => "0000000010100100001000",
			316 => "0000001010101000000100",
			317 => "0000000000010101010001",
			318 => "0000000000010101010001",
			319 => "0000000000010101010001",
			320 => "0000101100100100000100",
			321 => "0000000000010101010001",
			322 => "0010110111011100000100",
			323 => "0000000000010101010001",
			324 => "0000000000010101010001",
			325 => "0000001010111000010100",
			326 => "0000010001110000000100",
			327 => "0000000000010101010001",
			328 => "0010111001001000001000",
			329 => "0001001100000000000100",
			330 => "0000000000010101010001",
			331 => "0000000000010101010001",
			332 => "0001001111011000000100",
			333 => "0000000000010101010001",
			334 => "0000000000010101010001",
			335 => "0011100010110100001000",
			336 => "0010011001001000000100",
			337 => "0000000000010101010001",
			338 => "0000000000010101010001",
			339 => "0000000000010101010001",
			340 => "0011010101010101010100",
			341 => "0011000011010000101000",
			342 => "0010010101011100011000",
			343 => "0000001110110000010100",
			344 => "0010110110001100001000",
			345 => "0001001010100100000100",
			346 => "0000000000011000101101",
			347 => "0000000000011000101101",
			348 => "0001001010000100001000",
			349 => "0010010101010100000100",
			350 => "0000000000011000101101",
			351 => "0000000000011000101101",
			352 => "0000000000011000101101",
			353 => "0000000000011000101101",
			354 => "0011100001000000001000",
			355 => "0010111010100100000100",
			356 => "0000000000011000101101",
			357 => "0000000000011000101101",
			358 => "0011100110000100000100",
			359 => "0000000000011000101101",
			360 => "0000000000011000101101",
			361 => "0000010111110000010100",
			362 => "0001000101101100001000",
			363 => "0001110110101100000100",
			364 => "0000000000011000101101",
			365 => "0000000000011000101101",
			366 => "0001010110101100000100",
			367 => "0000000000011000101101",
			368 => "0000011000111100000100",
			369 => "0000000000011000101101",
			370 => "0000000000011000101101",
			371 => "0011110100111100010100",
			372 => "0000100110111100010000",
			373 => "0001101100000100001000",
			374 => "0010101011000000000100",
			375 => "0000000000011000101101",
			376 => "0000000000011000101101",
			377 => "0010110111011100000100",
			378 => "0000000000011000101101",
			379 => "0000000000011000101101",
			380 => "0000000000011000101101",
			381 => "0000000000011000101101",
			382 => "0010010011000000001100",
			383 => "0011000101011100001000",
			384 => "0011000101010100000100",
			385 => "0000000000011000101101",
			386 => "0000000000011000101101",
			387 => "0000000000011000101101",
			388 => "0001001111011000001100",
			389 => "0010001111011000001000",
			390 => "0010001010000100000100",
			391 => "0000000000011000101101",
			392 => "0000000000011000101101",
			393 => "0000000000011000101101",
			394 => "0000000000011000101101",
			395 => "0010011110011000000100",
			396 => "0000001000011010100001",
			397 => "0011011100101000101100",
			398 => "0010101111011000001000",
			399 => "0010001010100100000100",
			400 => "0000000000011010100001",
			401 => "1111111000011010100001",
			402 => "0010100011001000000100",
			403 => "0000001000011010100001",
			404 => "0001001100101000010000",
			405 => "0001000011010000001000",
			406 => "0000011001100000000100",
			407 => "0000000000011010100001",
			408 => "1111111000011010100001",
			409 => "0010010101011100000100",
			410 => "0000000000011010100001",
			411 => "1111111000011010100001",
			412 => "0000111000000000001000",
			413 => "0000010011110000000100",
			414 => "0000000000011010100001",
			415 => "1111111000011010100001",
			416 => "0000100110010100000100",
			417 => "0000000000011010100001",
			418 => "0000000000011010100001",
			419 => "0000010001100100001000",
			420 => "0000000111101100000100",
			421 => "0000000000011010100001",
			422 => "0000001000011010100001",
			423 => "1111111000011010100001",
			424 => "0001001100000000110100",
			425 => "0001001000000100110000",
			426 => "0010001111011000101100",
			427 => "0001100000001100011100",
			428 => "0000010001100100010000",
			429 => "0011000111011100001000",
			430 => "0001011101001000000100",
			431 => "0000000000011101001101",
			432 => "0000000000011101001101",
			433 => "0000010111100100000100",
			434 => "1111111000011101001101",
			435 => "0000001000011101001101",
			436 => "0001100101100000001000",
			437 => "0001111101101000000100",
			438 => "0000000000011101001101",
			439 => "1111111000011101001101",
			440 => "0000000000011101001101",
			441 => "0000001111001100000100",
			442 => "1111111000011101001101",
			443 => "0010011001000100001000",
			444 => "0011110111001100000100",
			445 => "0000000000011101001101",
			446 => "0000000000011101001101",
			447 => "0000000000011101001101",
			448 => "1111111000011101001101",
			449 => "0000001000011101001101",
			450 => "0001000110101100010000",
			451 => "0000001001101000001000",
			452 => "0000111100101100000100",
			453 => "1111111000011101001101",
			454 => "0000000000011101001101",
			455 => "0001100000000100000100",
			456 => "0000000000011101001101",
			457 => "1111111000011101001101",
			458 => "0011110001100000000100",
			459 => "1111111000011101001101",
			460 => "0000010111100100000100",
			461 => "0000001000011101001101",
			462 => "0000000000000000000100",
			463 => "1111111000011101001101",
			464 => "0000001101111000000100",
			465 => "0000001000011101001101",
			466 => "0000000000011101001101",
			467 => "0001001111011001010000",
			468 => "0000001010101000100000",
			469 => "0010001111111100010000",
			470 => "0010001001001100000100",
			471 => "0000000000100000110001",
			472 => "0011110001010100000100",
			473 => "0000000000100000110001",
			474 => "0001110110101100000100",
			475 => "0000000000100000110001",
			476 => "0000000000100000110001",
			477 => "0011010110001100000100",
			478 => "0000000000100000110001",
			479 => "0011100001101100000100",
			480 => "0000000000100000110001",
			481 => "0011100001000000000100",
			482 => "0000000000100000110001",
			483 => "0000000000100000110001",
			484 => "0011111100111100010000",
			485 => "0001111100110000001000",
			486 => "0011100010001000000100",
			487 => "0000000000100000110001",
			488 => "0000000000100000110001",
			489 => "0001011011111000000100",
			490 => "0000000000100000110001",
			491 => "0000000000100000110001",
			492 => "0001111101001000001100",
			493 => "0000110011100100001000",
			494 => "0000001110110000000100",
			495 => "0000000000100000110001",
			496 => "0000000000100000110001",
			497 => "0000000000100000110001",
			498 => "0001111001010000000100",
			499 => "0000000000100000110001",
			500 => "0001011101001000001000",
			501 => "0000010110010000000100",
			502 => "0000000000100000110001",
			503 => "0000000000100000110001",
			504 => "0000111001010000000100",
			505 => "0000000000100000110001",
			506 => "0000000000100000110001",
			507 => "0001001000000100001000",
			508 => "0001110100101100000100",
			509 => "0000000000100000110001",
			510 => "0000000000100000110001",
			511 => "0001001100000000000100",
			512 => "0000000000100000110001",
			513 => "0001000110101100001000",
			514 => "0000111100101100000100",
			515 => "0000000000100000110001",
			516 => "0000000000100000110001",
			517 => "0001000100101100001100",
			518 => "0011000101010100000100",
			519 => "0000000000100000110001",
			520 => "0000101000011100000100",
			521 => "0000000000100000110001",
			522 => "0000000000100000110001",
			523 => "0000000000100000110001",
			524 => "0001101010111101000100",
			525 => "0000100110101000110100",
			526 => "0001011100000000011000",
			527 => "0000110011000000001000",
			528 => "0010011010100100000100",
			529 => "0000000000100011111101",
			530 => "0000000000100011111101",
			531 => "0000010011110000001100",
			532 => "0000000101000100000100",
			533 => "0000000000100011111101",
			534 => "0001111001010000000100",
			535 => "0000000000100011111101",
			536 => "0000000000100011111101",
			537 => "0000000000100011111101",
			538 => "0000011000011000010100",
			539 => "0000010110010000001000",
			540 => "0011001110011000000100",
			541 => "0000000000100011111101",
			542 => "0000000000100011111101",
			543 => "0010101001000000001000",
			544 => "0001001010000100000100",
			545 => "0000000000100011111101",
			546 => "0000000000100011111101",
			547 => "0000000000100011111101",
			548 => "0011100110110000000100",
			549 => "0000000000100011111101",
			550 => "0000000000100011111101",
			551 => "0011100100001100000100",
			552 => "0000000000100011111101",
			553 => "0000000101101000001000",
			554 => "0010100011000100000100",
			555 => "0000000000100011111101",
			556 => "0000000000100011111101",
			557 => "0000000000100011111101",
			558 => "0000010001110000000100",
			559 => "0000000000100011111101",
			560 => "0011000101010100001000",
			561 => "0000001111010000000100",
			562 => "0000000000100011111101",
			563 => "0000000000100011111101",
			564 => "0010011010000100000100",
			565 => "0000000000100011111101",
			566 => "0011100110000100001100",
			567 => "0010111001001000000100",
			568 => "0000000000100011111101",
			569 => "0010111001000100000100",
			570 => "0000000000100011111101",
			571 => "0000000000100011111101",
			572 => "0011101000101100000100",
			573 => "0000000000100011111101",
			574 => "0000000000100011111101",
			575 => "0001101010111101010000",
			576 => "0011100011101100111000",
			577 => "0010010101011100010100",
			578 => "0000001001110100001100",
			579 => "0010001001001100000100",
			580 => "0000000000100111101001",
			581 => "0010110110001100000100",
			582 => "0000000000100111101001",
			583 => "0000000000100111101001",
			584 => "0001100001100000000100",
			585 => "0000001000100111101001",
			586 => "0000000000100111101001",
			587 => "0011000011010000010000",
			588 => "0010111010100100001100",
			589 => "0011100000110100001000",
			590 => "0001000101101100000100",
			591 => "0000000000100111101001",
			592 => "0000000000100111101001",
			593 => "1111111000100111101001",
			594 => "0000000000100111101001",
			595 => "0011100010110000010000",
			596 => "0010101000101000001000",
			597 => "0001001100101000000100",
			598 => "0000000000100111101001",
			599 => "0000000000100111101001",
			600 => "0000010111100100000100",
			601 => "0000000000100111101001",
			602 => "0000000000100111101001",
			603 => "0000000000100111101001",
			604 => "0000100110010100001100",
			605 => "0000000010100100001000",
			606 => "0000100111000100000100",
			607 => "0000000000100111101001",
			608 => "0000000000100111101001",
			609 => "0000000000100111101001",
			610 => "0000101100100100000100",
			611 => "0000001000100111101001",
			612 => "0000010111100100000100",
			613 => "1111111000100111101001",
			614 => "0000000000100111101001",
			615 => "0000101100100100000100",
			616 => "1111111000100111101001",
			617 => "0010000000110000010100",
			618 => "0010011001001000001000",
			619 => "0000010111110000000100",
			620 => "0000000000100111101001",
			621 => "1111111000100111101001",
			622 => "0001001111011000001000",
			623 => "0001100010000100000100",
			624 => "0000000000100111101001",
			625 => "0000000000100111101001",
			626 => "0000000000100111101001",
			627 => "0001001000111000001000",
			628 => "0000111100010000000100",
			629 => "0000000000100111101001",
			630 => "1111111000100111101001",
			631 => "0001001100010000000100",
			632 => "0000000000100111101001",
			633 => "0000000000100111101001",
			634 => "0011010101010101011000",
			635 => "0011000011010000101100",
			636 => "0001001010000100100100",
			637 => "0001101010111100011000",
			638 => "0000001011010000010000",
			639 => "0011001010100100001000",
			640 => "0001010110001100000100",
			641 => "0000000000101011101101",
			642 => "0000000000101011101101",
			643 => "0011101100100000000100",
			644 => "0000000000101011101101",
			645 => "0000000000101011101101",
			646 => "0010010101011100000100",
			647 => "0000000000101011101101",
			648 => "0000000000101011101101",
			649 => "0001000101011100001000",
			650 => "0001001010100100000100",
			651 => "0000000000101011101101",
			652 => "0000000000101011101101",
			653 => "0000000000101011101101",
			654 => "0010111010100100000100",
			655 => "0000000000101011101101",
			656 => "0000000000101011101101",
			657 => "0010101111101000010100",
			658 => "0000110011000000000100",
			659 => "0000000000101011101101",
			660 => "0000010001100100001100",
			661 => "0001111100000000000100",
			662 => "0000000000101011101101",
			663 => "0000111100010000000100",
			664 => "0000000000101011101101",
			665 => "0000000000101011101101",
			666 => "0000000000101011101101",
			667 => "0010001001000100001100",
			668 => "0011011010100100000100",
			669 => "0000000000101011101101",
			670 => "0010110101010100000100",
			671 => "0000000000101011101101",
			672 => "0000000000101011101101",
			673 => "0001010110011100000100",
			674 => "0000000000101011101101",
			675 => "0001001111101000000100",
			676 => "0000000000101011101101",
			677 => "0000000000101011101101",
			678 => "0001011100101100010100",
			679 => "0000001000001100010000",
			680 => "0010111100101000001000",
			681 => "0010001010000100000100",
			682 => "0000000000101011101101",
			683 => "0000000000101011101101",
			684 => "0010111001001000000100",
			685 => "0000000000101011101101",
			686 => "0000000000101011101101",
			687 => "0000000000101011101101",
			688 => "0001011001011000001100",
			689 => "0000000000000000000100",
			690 => "0000000000101011101101",
			691 => "0000101011001100000100",
			692 => "0000000000101011101101",
			693 => "0000000000101011101101",
			694 => "0000000010100100001000",
			695 => "0000001001110100000100",
			696 => "0000000000101011101101",
			697 => "0000000000101011101101",
			698 => "0000000000101011101101",
			699 => "0000000011111000100100",
			700 => "0010010101101100011000",
			701 => "0010001001001100000100",
			702 => "0000000000101111010001",
			703 => "0010001111111100001100",
			704 => "0001101110001100000100",
			705 => "0000000000101111010001",
			706 => "0011100010010100000100",
			707 => "0000000000101111010001",
			708 => "0000000000101111010001",
			709 => "0001100111100000000100",
			710 => "0000000000101111010001",
			711 => "0000000000101111010001",
			712 => "0011010110001100001000",
			713 => "0001000110000000000100",
			714 => "0000000000101111010001",
			715 => "0000000000101111010001",
			716 => "1111111000101111010001",
			717 => "0001101010111100110000",
			718 => "0000010111100100011000",
			719 => "0010010101011100001000",
			720 => "0001001101101000000100",
			721 => "0000000000101111010001",
			722 => "0000000000101111010001",
			723 => "0000110011001000000100",
			724 => "1111111000101111010001",
			725 => "0001100101100000001000",
			726 => "0011111011011100000100",
			727 => "0000000000101111010001",
			728 => "0000000000101111010001",
			729 => "0000000000101111010001",
			730 => "0000001011100100010000",
			731 => "0010101000101000000100",
			732 => "0000000000101111010001",
			733 => "0010110101010100000100",
			734 => "0000000000101111010001",
			735 => "0000001111101100000100",
			736 => "0000000000101111010001",
			737 => "0000000000101111010001",
			738 => "0001010011000100000100",
			739 => "0000001000101111010001",
			740 => "0000000000101111010001",
			741 => "0000101100100100000100",
			742 => "1111111000101111010001",
			743 => "0001111101001000000100",
			744 => "0000000000101111010001",
			745 => "0001001111011000001100",
			746 => "0000111001010000001000",
			747 => "0010011001000100000100",
			748 => "0000000000101111010001",
			749 => "0000001000101111010001",
			750 => "0000000000101111010001",
			751 => "0010010101111000000100",
			752 => "0000000000101111010001",
			753 => "0000111011111000000100",
			754 => "0000000000101111010001",
			755 => "0000000000101111010001",
			756 => "0001101010101101011100",
			757 => "0011100011101101000000",
			758 => "0001011100000000010100",
			759 => "0000110011000000001000",
			760 => "0010011010100100000100",
			761 => "0000000000110011000101",
			762 => "0000000000110011000101",
			763 => "0000010011110000001000",
			764 => "0000000101000100000100",
			765 => "0000000000110011000101",
			766 => "0000000000110011000101",
			767 => "0000000000110011000101",
			768 => "0001000011000000010000",
			769 => "0010010101011100000100",
			770 => "0000000000110011000101",
			771 => "0001111000101000001000",
			772 => "0001101100011000000100",
			773 => "0000000000110011000101",
			774 => "0000000000110011000101",
			775 => "0000000000110011000101",
			776 => "0010101011000000001100",
			777 => "0011010011010000001000",
			778 => "0011010110001100000100",
			779 => "0000000000110011000101",
			780 => "0000000000110011000101",
			781 => "0000000000110011000101",
			782 => "0011010101010100001000",
			783 => "0010001001000100000100",
			784 => "0000000000110011000101",
			785 => "0000000000110011000101",
			786 => "0010001001000100000100",
			787 => "0000000000110011000101",
			788 => "0000000000110011000101",
			789 => "0000100110010100001100",
			790 => "0000000010100100001000",
			791 => "0000001010101000000100",
			792 => "0000000000110011000101",
			793 => "0000000000110011000101",
			794 => "0000000000110011000101",
			795 => "0000001110110000001100",
			796 => "0010100011000100001000",
			797 => "0000100110111100000100",
			798 => "0000000000110011000101",
			799 => "0000000000110011000101",
			800 => "0000000000110011000101",
			801 => "0000000000110011000101",
			802 => "0000001010111000010100",
			803 => "0000010001110000000100",
			804 => "0000000000110011000101",
			805 => "0010111001001000001000",
			806 => "0001001100000000000100",
			807 => "0000000000110011000101",
			808 => "0000000000110011000101",
			809 => "0001001111011000000100",
			810 => "0000000000110011000101",
			811 => "0000000000110011000101",
			812 => "0001111100101100001000",
			813 => "0010011001001000000100",
			814 => "0000000000110011000101",
			815 => "0000000000110011000101",
			816 => "0000000000110011000101",
			817 => "0000100110010100111000",
			818 => "0000010001100100101000",
			819 => "0010101111101000011000",
			820 => "0001100100110000010100",
			821 => "0000001011111100001100",
			822 => "0001111100010000001000",
			823 => "0010001001001100000100",
			824 => "0000000000110110110001",
			825 => "0000000000110110110001",
			826 => "1111111000110110110001",
			827 => "0010101000111000000100",
			828 => "0000000000110110110001",
			829 => "0000001000110110110001",
			830 => "0000000000110110110001",
			831 => "0010011101101000000100",
			832 => "1111111000110110110001",
			833 => "0010001111001000000100",
			834 => "0000000000110110110001",
			835 => "0000100111001100000100",
			836 => "0000000000110110110001",
			837 => "0000000000110110110001",
			838 => "0000011111001000001100",
			839 => "0010101001000000000100",
			840 => "1111111000110110110001",
			841 => "0001100110000100000100",
			842 => "0000000000110110110001",
			843 => "0000000000110110110001",
			844 => "0000000000110110110001",
			845 => "0001111001011000110100",
			846 => "0000000101101000011100",
			847 => "0010111010100100010000",
			848 => "0011011011101100001100",
			849 => "0000001101110000000100",
			850 => "0000000000110110110001",
			851 => "0011110110011000000100",
			852 => "0000000000110110110001",
			853 => "0000000000110110110001",
			854 => "0000000000110110110001",
			855 => "0010001111001000000100",
			856 => "0000001000110110110001",
			857 => "0000001101111000000100",
			858 => "0000000000110110110001",
			859 => "0000000000110110110001",
			860 => "0011110011111100010100",
			861 => "0001101110101100010000",
			862 => "0010000101011100001000",
			863 => "0001010110101100000100",
			864 => "0000000000110110110001",
			865 => "1111111000110110110001",
			866 => "0010010101101100000100",
			867 => "0000000000110110110001",
			868 => "0000000000110110110001",
			869 => "0000000000110110110001",
			870 => "0000000000110110110001",
			871 => "0000100101101000000100",
			872 => "1111111000110110110001",
			873 => "0001100111010000000100",
			874 => "0000000000110110110001",
			875 => "0000000000110110110001",
			876 => "0000100101011000010100",
			877 => "0001000111110000001000",
			878 => "0001000001110000000100",
			879 => "0000000000111001010101",
			880 => "0000000000111001010101",
			881 => "0001010110011100000100",
			882 => "0000000000111001010101",
			883 => "0000001110100000000100",
			884 => "0000000000111001010101",
			885 => "0000000000111001010101",
			886 => "0000010110110100111000",
			887 => "0000110011000000000100",
			888 => "0000000000111001010101",
			889 => "0001101101010000100000",
			890 => "0000010110010000010000",
			891 => "0001001001000100001000",
			892 => "0010010101011100000100",
			893 => "0000000000111001010101",
			894 => "0000000000111001010101",
			895 => "0011001110011000000100",
			896 => "0000000000111001010101",
			897 => "0000000000111001010101",
			898 => "0000100110010100001000",
			899 => "0000010001100100000100",
			900 => "0000000000111001010101",
			901 => "0000000000111001010101",
			902 => "0001011001010100000100",
			903 => "0000000000111001010101",
			904 => "0000000000111001010101",
			905 => "0000010110010000000100",
			906 => "0000000000111001010101",
			907 => "0011110011111100001000",
			908 => "0001001111011000000100",
			909 => "0000000000111001010101",
			910 => "0000000000111001010101",
			911 => "0011110111001100000100",
			912 => "0000000000111001010101",
			913 => "0000000000111001010101",
			914 => "0000010011000000000100",
			915 => "0000000000111001010101",
			916 => "0000000000111001010101",
			917 => "0000000011111000011100",
			918 => "0001110110101100011000",
			919 => "0010001001001100000100",
			920 => "0000000000111100011001",
			921 => "0011111101100100010000",
			922 => "0001000111110000000100",
			923 => "0000000000111100011001",
			924 => "0010011101101000000100",
			925 => "0000000000111100011001",
			926 => "0010011010000100000100",
			927 => "0000000000111100011001",
			928 => "0000000000111100011001",
			929 => "0000000000111100011001",
			930 => "0000000000111100011001",
			931 => "0011010011010000110000",
			932 => "0001110110101100010000",
			933 => "0011100010001000000100",
			934 => "0000000000111100011001",
			935 => "0001000101010100000100",
			936 => "0000000000111100011001",
			937 => "0001100100000100000100",
			938 => "0000000000111100011001",
			939 => "0000000000111100011001",
			940 => "0010100100101100010100",
			941 => "0011101000101100010000",
			942 => "0001001001000100001000",
			943 => "0010111110011000000100",
			944 => "0000000000111100011001",
			945 => "0000000000111100011001",
			946 => "0010000101101100000100",
			947 => "0000000000111100011001",
			948 => "0000000000111100011001",
			949 => "0000000000111100011001",
			950 => "0001001000000000001000",
			951 => "0011101100011000000100",
			952 => "0000000000111100011001",
			953 => "0000000000111100011001",
			954 => "0000000000111100011001",
			955 => "0000000010100100000100",
			956 => "0000000000111100011001",
			957 => "0001011101001000000100",
			958 => "0000000000111100011001",
			959 => "0001010011000100001100",
			960 => "0000101000010000000100",
			961 => "0000000000111100011001",
			962 => "0001001111011000000100",
			963 => "0000000000111100011001",
			964 => "0000000000111100011001",
			965 => "0000000000111100011001",
			966 => "0011100100011100101100",
			967 => "0010101110111000101000",
			968 => "0010011010100100000100",
			969 => "0000001000111101110101",
			970 => "0000110011000000000100",
			971 => "1111111000111101110101",
			972 => "0011000101011100010000",
			973 => "0010001010000100001000",
			974 => "0010101011000000000100",
			975 => "0000000000111101110101",
			976 => "0000000000111101110101",
			977 => "0000010011110000000100",
			978 => "0000000000111101110101",
			979 => "1111111000111101110101",
			980 => "0011011010100100001000",
			981 => "0000010111100100000100",
			982 => "1111111000111101110101",
			983 => "0000001000111101110101",
			984 => "0010011010000100000100",
			985 => "0000001000111101110101",
			986 => "0000000000111101110101",
			987 => "1111111000111101110101",
			988 => "1111111000111101110101",
			989 => "0010111010100100101000",
			990 => "0001100000001100011100",
			991 => "0001011111101000011000",
			992 => "0000101101110000010100",
			993 => "0001101110001000010000",
			994 => "0010010101011100001000",
			995 => "0010110110001100000100",
			996 => "0000000001000001011001",
			997 => "0000000001000001011001",
			998 => "0001111001010000000100",
			999 => "0000000001000001011001",
			1000 => "0000001001000001011001",
			1001 => "0000001001000001011001",
			1002 => "0000000001000001011001",
			1003 => "1111111001000001011001",
			1004 => "0001101110000100000100",
			1005 => "1111111001000001011001",
			1006 => "0010000101101100000100",
			1007 => "0000000001000001011001",
			1008 => "1111111001000001011001",
			1009 => "0000000000101000101000",
			1010 => "0000010001100100011100",
			1011 => "0000010110010000001000",
			1012 => "0010011001001000000100",
			1013 => "0000000001000001011001",
			1014 => "1111111001000001011001",
			1015 => "0001111001010100001000",
			1016 => "0000100100111100000100",
			1017 => "0000000001000001011001",
			1018 => "0000001001000001011001",
			1019 => "0001111000101000000100",
			1020 => "1111111001000001011001",
			1021 => "0000001101110100000100",
			1022 => "0000000001000001011001",
			1023 => "0000001001000001011001",
			1024 => "0010101001000000000100",
			1025 => "1111111001000001011001",
			1026 => "0001100100000100000100",
			1027 => "0000000001000001011001",
			1028 => "0000000001000001011001",
			1029 => "0000110011100100000100",
			1030 => "0000000001000001011001",
			1031 => "0011100110110000001000",
			1032 => "0000010111100100000100",
			1033 => "0000000001000001011001",
			1034 => "0000001001000001011001",
			1035 => "0000111001010000001000",
			1036 => "0011100010110100000100",
			1037 => "0000001001000001011001",
			1038 => "0000000001000001011001",
			1039 => "0010101011000000001000",
			1040 => "0001011100101100000100",
			1041 => "0000000001000001011001",
			1042 => "1111111001000001011001",
			1043 => "0000011110011000000100",
			1044 => "0000000001000001011001",
			1045 => "0000000001000001011001",
			1046 => "0000000011111000100100",
			1047 => "0001111100010000011100",
			1048 => "0010111010100100010000",
			1049 => "0001000111110000000100",
			1050 => "0000000001000101011101",
			1051 => "0000011001100100001000",
			1052 => "0001010011001000000100",
			1053 => "0000000001000101011101",
			1054 => "0000000001000101011101",
			1055 => "0000000001000101011101",
			1056 => "0001111100000000000100",
			1057 => "0000000001000101011101",
			1058 => "0011000111011100000100",
			1059 => "0000000001000101011101",
			1060 => "0000000001000101011101",
			1061 => "0010011100101000000100",
			1062 => "0000000001000101011101",
			1063 => "0000000001000101011101",
			1064 => "0011111100111100101000",
			1065 => "0010010101011100001000",
			1066 => "0001111100010000000100",
			1067 => "0000000001000101011101",
			1068 => "0000000001000101011101",
			1069 => "0000010111100100001000",
			1070 => "0011111110101100000100",
			1071 => "0000000001000101011101",
			1072 => "0000000001000101011101",
			1073 => "0001001100000000001100",
			1074 => "0000010001100100000100",
			1075 => "0000000001000101011101",
			1076 => "0011110111000000000100",
			1077 => "0000000001000101011101",
			1078 => "0000000001000101011101",
			1079 => "0000111100101100000100",
			1080 => "0000000001000101011101",
			1081 => "0000110011000100000100",
			1082 => "0000000001000101011101",
			1083 => "0000000001000101011101",
			1084 => "0011111101001100010100",
			1085 => "0001001111011000001100",
			1086 => "0011010110110100000100",
			1087 => "0000000001000101011101",
			1088 => "0010110111011100000100",
			1089 => "0000000001000101011101",
			1090 => "0000000001000101011101",
			1091 => "0000111111101000000100",
			1092 => "0000000001000101011101",
			1093 => "0000000001000101011101",
			1094 => "0011100011101000010100",
			1095 => "0001011100110000001000",
			1096 => "0000010111100100000100",
			1097 => "0000000001000101011101",
			1098 => "0000000001000101011101",
			1099 => "0001101101010000001000",
			1100 => "0011011011101100000100",
			1101 => "0000000001000101011101",
			1102 => "0000000001000101011101",
			1103 => "0000000001000101011101",
			1104 => "0001110001010000000100",
			1105 => "0000000001000101011101",
			1106 => "0010010101111000000100",
			1107 => "0000000001000101011101",
			1108 => "0001101110101100000100",
			1109 => "0000000001000101011101",
			1110 => "0000000001000101011101",
			1111 => "0000101011101000010100",
			1112 => "0011011110011000000100",
			1113 => "1111111001001000010001",
			1114 => "0011000111011100001100",
			1115 => "0010001111001000001000",
			1116 => "0001111100000000000100",
			1117 => "0000000001001000010001",
			1118 => "0000001001001000010001",
			1119 => "1111111001001000010001",
			1120 => "1111111001001000010001",
			1121 => "0001110011000101000100",
			1122 => "0010111010100100101000",
			1123 => "0000010001110000010000",
			1124 => "0011001110011000001000",
			1125 => "0000000111111000000100",
			1126 => "0000001001001000010001",
			1127 => "0000000001001000010001",
			1128 => "0011101101100000000100",
			1129 => "0000000001001000010001",
			1130 => "0000001001001000010001",
			1131 => "0001101010111100001100",
			1132 => "0001001010000100001000",
			1133 => "0000110011001000000100",
			1134 => "0000000001001000010001",
			1135 => "0000000001001000010001",
			1136 => "1111111001001000010001",
			1137 => "0001001100101000001000",
			1138 => "0000001010111000000100",
			1139 => "1111111001001000010001",
			1140 => "0000000001001000010001",
			1141 => "1111111001001000010001",
			1142 => "0011011110011000001000",
			1143 => "0010000101011100000100",
			1144 => "0000000001001000010001",
			1145 => "0000001001001000010001",
			1146 => "0000010110010000000100",
			1147 => "1111111001001000010001",
			1148 => "0000000110111100001000",
			1149 => "0000011000011000000100",
			1150 => "0000001001001000010001",
			1151 => "0000000001001000010001",
			1152 => "0011100001000000000100",
			1153 => "0000000001001000010001",
			1154 => "0000000001001000010001",
			1155 => "1111111001001000010001",
			1156 => "0011010110001100110000",
			1157 => "0010111110011000011100",
			1158 => "0000110011001000010000",
			1159 => "0010100011000000001100",
			1160 => "0000110110110100000100",
			1161 => "0000000001001100110101",
			1162 => "0001001110011000000100",
			1163 => "0000000001001100110101",
			1164 => "0000000001001100110101",
			1165 => "0000000001001100110101",
			1166 => "0011110111010000000100",
			1167 => "0000000001001100110101",
			1168 => "0010101111101000000100",
			1169 => "0000000001001100110101",
			1170 => "0000000001001100110101",
			1171 => "0011011101000000000100",
			1172 => "0000000001001100110101",
			1173 => "0001101000110100001100",
			1174 => "0010101100010000001000",
			1175 => "0000110011000000000100",
			1176 => "0000000001001100110101",
			1177 => "0000000001001100110101",
			1178 => "0000000001001100110101",
			1179 => "0000001001001100110101",
			1180 => "0001000110000000101100",
			1181 => "0011101100011000011100",
			1182 => "0011100000110100010100",
			1183 => "0010000101011100001000",
			1184 => "0010111010100100000100",
			1185 => "0000000001001100110101",
			1186 => "0000000001001100110101",
			1187 => "0001011111011000001000",
			1188 => "0001111000111000000100",
			1189 => "0000000001001100110101",
			1190 => "0000000001001100110101",
			1191 => "0000000001001100110101",
			1192 => "0001011111011000000100",
			1193 => "0000000001001100110101",
			1194 => "1111111001001100110101",
			1195 => "0010011001000100001100",
			1196 => "0001100000001100000100",
			1197 => "0000000001001100110101",
			1198 => "0011110111001100000100",
			1199 => "1111111001001100110101",
			1200 => "0000000001001100110101",
			1201 => "0000000001001100110101",
			1202 => "0010101000101000010100",
			1203 => "0000010011110000001100",
			1204 => "0000010110010000000100",
			1205 => "0000000001001100110101",
			1206 => "0001111100000000000100",
			1207 => "0000000001001100110101",
			1208 => "0000001001001100110101",
			1209 => "0011001100101000000100",
			1210 => "0000000001001100110101",
			1211 => "0000000001001100110101",
			1212 => "0011000101010100001100",
			1213 => "0010001001001100000100",
			1214 => "0000000001001100110101",
			1215 => "0000001101111000000100",
			1216 => "1111111001001100110101",
			1217 => "0000000001001100110101",
			1218 => "0001010100101100001000",
			1219 => "0011100001000000000100",
			1220 => "0000000001001100110101",
			1221 => "0000000001001100110101",
			1222 => "0010101011111000001000",
			1223 => "0010100100101100000100",
			1224 => "0000000001001100110101",
			1225 => "0000000001001100110101",
			1226 => "0011101110100000000100",
			1227 => "0000000001001100110101",
			1228 => "0000000001001100110101",
			1229 => "0000001001110100101100",
			1230 => "0011001010100100000100",
			1231 => "0000000001010000000001",
			1232 => "0001010110101100010100",
			1233 => "0011111101100100000100",
			1234 => "0000000001010000000001",
			1235 => "0010011001000100001100",
			1236 => "0001010101111000000100",
			1237 => "0000000001010000000001",
			1238 => "0011100001000100000100",
			1239 => "0000000001010000000001",
			1240 => "0000000001010000000001",
			1241 => "0000000001010000000001",
			1242 => "0011101001011100010000",
			1243 => "0011011010100100001100",
			1244 => "0001001000101000001000",
			1245 => "0000111100010000000100",
			1246 => "0000000001010000000001",
			1247 => "0000000001010000000001",
			1248 => "0000000001010000000001",
			1249 => "0000000001010000000001",
			1250 => "0000000001010000000001",
			1251 => "0001100101000000001000",
			1252 => "0000011000011000000100",
			1253 => "0000000001010000000001",
			1254 => "0000000001010000000001",
			1255 => "0000100110010100001100",
			1256 => "0000100011111000000100",
			1257 => "0000000001010000000001",
			1258 => "0011001110011000000100",
			1259 => "0000000001010000000001",
			1260 => "0000000001010000000001",
			1261 => "0001101010111100010100",
			1262 => "0000010110010000001100",
			1263 => "0011001110011000000100",
			1264 => "0000000001010000000001",
			1265 => "0000100110100100000100",
			1266 => "0000000001010000000001",
			1267 => "0000000001010000000001",
			1268 => "0001010011000100000100",
			1269 => "0000000001010000000001",
			1270 => "0000000001010000000001",
			1271 => "0000010001110000000100",
			1272 => "0000000001010000000001",
			1273 => "0000001010111000001000",
			1274 => "0001011100101100000100",
			1275 => "0000000001010000000001",
			1276 => "0000000001010000000001",
			1277 => "0001110100101100000100",
			1278 => "0000000001010000000001",
			1279 => "0000000001010000000001",
			1280 => "0001001100000001000100",
			1281 => "0001001000000101000000",
			1282 => "0010011101101000101100",
			1283 => "0000010001100100100000",
			1284 => "0010011001001000010000",
			1285 => "0001101010101100001000",
			1286 => "0011011110011000000100",
			1287 => "0000000001010010111101",
			1288 => "0000000001010010111101",
			1289 => "0000010111110000000100",
			1290 => "0000000001010010111101",
			1291 => "1111111001010010111101",
			1292 => "0011100001101100001000",
			1293 => "0010101101001000000100",
			1294 => "0000000001010010111101",
			1295 => "0000000001010010111101",
			1296 => "0010100100101100000100",
			1297 => "0000000001010010111101",
			1298 => "0000000001010010111101",
			1299 => "0000100100010100001000",
			1300 => "0000111001000100000100",
			1301 => "0000000001010010111101",
			1302 => "1111111001010010111101",
			1303 => "0000000001010010111101",
			1304 => "0010101011000000010000",
			1305 => "0001100001111000001100",
			1306 => "0001111111101000000100",
			1307 => "0000000001010010111101",
			1308 => "0011111010101100000100",
			1309 => "0000000001010010111101",
			1310 => "0000000001010010111101",
			1311 => "1111111001010010111101",
			1312 => "0000000001010010111101",
			1313 => "0000001001010010111101",
			1314 => "0001001000111000000100",
			1315 => "1111111001010010111101",
			1316 => "0000000000000000001100",
			1317 => "0000010111100100001000",
			1318 => "0000010110010000000100",
			1319 => "0000000001010010111101",
			1320 => "0000000001010010111101",
			1321 => "1111111001010010111101",
			1322 => "0001010000111100001000",
			1323 => "0011100011101000000100",
			1324 => "0000000001010010111101",
			1325 => "0000000001010010111101",
			1326 => "0000000001010010111101",
			1327 => "0011111100111101011000",
			1328 => "0000000011111000110100",
			1329 => "0001000101101100011100",
			1330 => "0001001100101000010000",
			1331 => "0001000111110000001000",
			1332 => "0001000001110000000100",
			1333 => "0000000001010111100001",
			1334 => "0000000001010111100001",
			1335 => "0011111000010100000100",
			1336 => "0000000001010111100001",
			1337 => "0000000001010111100001",
			1338 => "0001111000000000000100",
			1339 => "0000000001010111100001",
			1340 => "0001111001010000000100",
			1341 => "0000000001010111100001",
			1342 => "0000000001010111100001",
			1343 => "0010011101101000001000",
			1344 => "0011100101110100000100",
			1345 => "0000000001010111100001",
			1346 => "0000000001010111100001",
			1347 => "0010110101010100001100",
			1348 => "0010110111011100000100",
			1349 => "0000000001010111100001",
			1350 => "0010011010000100000100",
			1351 => "0000000001010111100001",
			1352 => "0000000001010111100001",
			1353 => "0000000001010111100001",
			1354 => "0001001100000000010100",
			1355 => "0010101000111000000100",
			1356 => "0000000001010111100001",
			1357 => "0000010000011000000100",
			1358 => "0000000001010111100001",
			1359 => "0000010001100100000100",
			1360 => "0000000001010111100001",
			1361 => "0011011100101000000100",
			1362 => "0000000001010111100001",
			1363 => "0000000001010111100001",
			1364 => "0000111100101100001000",
			1365 => "0011100110110000000100",
			1366 => "0000000001010111100001",
			1367 => "0000000001010111100001",
			1368 => "0000110011000100000100",
			1369 => "0000000001010111100001",
			1370 => "0000000001010111100001",
			1371 => "0011111101001100010100",
			1372 => "0011010110001100001000",
			1373 => "0010101001010100000100",
			1374 => "0000000001010111100001",
			1375 => "0000000001010111100001",
			1376 => "0001010110011100000100",
			1377 => "0000000001010111100001",
			1378 => "0001010000111100000100",
			1379 => "0000000001010111100001",
			1380 => "0000000001010111100001",
			1381 => "0000010001110000000100",
			1382 => "0000000001010111100001",
			1383 => "0011000101010100010000",
			1384 => "0000001000110000001100",
			1385 => "0001100000001100000100",
			1386 => "0000000001010111100001",
			1387 => "0001000011010000000100",
			1388 => "0000000001010111100001",
			1389 => "0000000001010111100001",
			1390 => "0000000001010111100001",
			1391 => "0000001101011000001100",
			1392 => "0001010011000100001000",
			1393 => "0001101110101100000100",
			1394 => "0000000001010111100001",
			1395 => "0000000001010111100001",
			1396 => "0000000001010111100001",
			1397 => "0000111001010100000100",
			1398 => "0000000001010111100001",
			1399 => "0000000001010111100001",
			1400 => "0001111001011001001100",
			1401 => "0011100110000101001000",
			1402 => "0011100011101100101000",
			1403 => "0010010101011100010100",
			1404 => "0001001001001000001100",
			1405 => "0010101000000100001000",
			1406 => "0001010110110100000100",
			1407 => "0000001001011010001101",
			1408 => "0000000001011010001101",
			1409 => "0000001001011010001101",
			1410 => "0000110011100100000100",
			1411 => "0000000001011010001101",
			1412 => "0000000001011010001101",
			1413 => "0000010000011000000100",
			1414 => "1111111001011010001101",
			1415 => "0001000011000000001000",
			1416 => "0001011100000000000100",
			1417 => "0000000001011010001101",
			1418 => "0000000001011010001101",
			1419 => "0010101011000000000100",
			1420 => "0000001001011010001101",
			1421 => "0000000001011010001101",
			1422 => "0000000110111100001100",
			1423 => "0000000010100100001000",
			1424 => "0011110010010000000100",
			1425 => "0000000001011010001101",
			1426 => "0000000001011010001101",
			1427 => "1111111001011010001101",
			1428 => "0001101010111100001000",
			1429 => "0000100110111100000100",
			1430 => "0000001001011010001101",
			1431 => "0000000001011010001101",
			1432 => "0000010001110000000100",
			1433 => "0000001001011010001101",
			1434 => "0001011101001000000100",
			1435 => "0000000001011010001101",
			1436 => "0000000001011010001101",
			1437 => "1111111001011010001101",
			1438 => "0000100101101000000100",
			1439 => "1111111001011010001101",
			1440 => "0000100101101000000100",
			1441 => "0000000001011010001101",
			1442 => "0000000001011010001101",
			1443 => "0011111101100100010000",
			1444 => "0010011010100100000100",
			1445 => "0000000001011101000001",
			1446 => "0011000111011100001000",
			1447 => "0010010110000000000100",
			1448 => "1111111001011101000001",
			1449 => "0000000001011101000001",
			1450 => "1111111001011101000001",
			1451 => "0010011111011001001000",
			1452 => "0001101010111100110000",
			1453 => "0000010110010000011000",
			1454 => "0011001110011000001000",
			1455 => "0000001101011100000100",
			1456 => "0000000001011101000001",
			1457 => "0000001001011101000001",
			1458 => "0000111000000000001000",
			1459 => "0001011111011000000100",
			1460 => "1111111001011101000001",
			1461 => "0000001001011101000001",
			1462 => "0000000010101100000100",
			1463 => "0000000001011101000001",
			1464 => "1111111001011101000001",
			1465 => "0000000110111100010000",
			1466 => "0000010001100100001000",
			1467 => "0011000011010000000100",
			1468 => "0000000001011101000001",
			1469 => "0000001001011101000001",
			1470 => "0010101101001000000100",
			1471 => "0000000001011101000001",
			1472 => "1111111001011101000001",
			1473 => "0011010111011100000100",
			1474 => "0000001001011101000001",
			1475 => "0000001001011101000001",
			1476 => "0011111101001100001000",
			1477 => "0001111100101100000100",
			1478 => "1111111001011101000001",
			1479 => "0000000001011101000001",
			1480 => "0010111011101100000100",
			1481 => "1111111001011101000001",
			1482 => "0000010001110000000100",
			1483 => "0000001001011101000001",
			1484 => "0000101010010100000100",
			1485 => "1111111001011101000001",
			1486 => "0000001001011101000001",
			1487 => "1111111001011101000001",
			1488 => "0011010110001100110000",
			1489 => "0010111110011000011100",
			1490 => "0000110011001000010000",
			1491 => "0010100011000000001100",
			1492 => "0000110110110100000100",
			1493 => "0000000001100010000101",
			1494 => "0001001110011000000100",
			1495 => "0000000001100010000101",
			1496 => "0000000001100010000101",
			1497 => "0000000001100010000101",
			1498 => "0011110111010000000100",
			1499 => "0000000001100010000101",
			1500 => "0010101111101000000100",
			1501 => "0000000001100010000101",
			1502 => "0000000001100010000101",
			1503 => "0001000011000000010000",
			1504 => "0000110011001000001000",
			1505 => "0010010101011100000100",
			1506 => "0000000001100010000101",
			1507 => "0000000001100010000101",
			1508 => "0001011101001000000100",
			1509 => "0000001001100010000101",
			1510 => "0000000001100010000101",
			1511 => "0000000001100010000101",
			1512 => "0001000110000000101100",
			1513 => "0011101100011000011100",
			1514 => "0011100000110100010100",
			1515 => "0010000101011100001000",
			1516 => "0010111010100100000100",
			1517 => "0000000001100010000101",
			1518 => "0000000001100010000101",
			1519 => "0001011111011000001000",
			1520 => "0010101000000100000100",
			1521 => "0000000001100010000101",
			1522 => "0000000001100010000101",
			1523 => "0000000001100010000101",
			1524 => "0001011111011000000100",
			1525 => "0000000001100010000101",
			1526 => "1111111001100010000101",
			1527 => "0010011001000100001100",
			1528 => "0001100000001100000100",
			1529 => "0000000001100010000101",
			1530 => "0011110111001100000100",
			1531 => "1111111001100010000101",
			1532 => "0000000001100010000101",
			1533 => "0000000001100010000101",
			1534 => "0001010100101100100000",
			1535 => "0001100011101000001100",
			1536 => "0001111000111000001000",
			1537 => "0000010111100100000100",
			1538 => "0000000001100010000101",
			1539 => "0000000001100010000101",
			1540 => "0000000001100010000101",
			1541 => "0001110100101100001100",
			1542 => "0010000101011100000100",
			1543 => "0000000001100010000101",
			1544 => "0011111101010100000100",
			1545 => "0000000001100010000101",
			1546 => "0000001001100010000101",
			1547 => "0000111101001000000100",
			1548 => "0000000001100010000101",
			1549 => "0000000001100010000101",
			1550 => "0001010110011100010000",
			1551 => "0011111011000100001000",
			1552 => "0000011101000000000100",
			1553 => "1111111001100010000101",
			1554 => "0000000001100010000101",
			1555 => "0011100110000100000100",
			1556 => "0000000001100010000101",
			1557 => "0000000001100010000101",
			1558 => "0001011001011000001000",
			1559 => "0010000011001000000100",
			1560 => "0000000001100010000101",
			1561 => "0000000001100010000101",
			1562 => "0000000010100100001000",
			1563 => "0011110001100000000100",
			1564 => "0000000001100010000101",
			1565 => "0000000001100010000101",
			1566 => "0010110101010100000100",
			1567 => "0000000001100010000101",
			1568 => "0000000001100010000101",
			1569 => "0010110110001100001000",
			1570 => "0011001101000000000100",
			1571 => "0000000001100100111001",
			1572 => "1111111001100100111001",
			1573 => "0001000011010000011000",
			1574 => "0000011001100100000100",
			1575 => "1111111001100100111001",
			1576 => "0011000111011100010000",
			1577 => "0011100110000100001100",
			1578 => "0001101110001100000100",
			1579 => "0000000001100100111001",
			1580 => "0000010111100100000100",
			1581 => "0000001001100100111001",
			1582 => "0000000001100100111001",
			1583 => "0000000001100100111001",
			1584 => "1111111001100100111001",
			1585 => "0010100000111100110100",
			1586 => "0001100010000100011100",
			1587 => "0011111101001100010000",
			1588 => "0001101010111100001000",
			1589 => "0000110011001000000100",
			1590 => "0000000001100100111001",
			1591 => "0000000001100100111001",
			1592 => "0001010110011100000100",
			1593 => "1111111001100100111001",
			1594 => "0000000001100100111001",
			1595 => "0011001010100100000100",
			1596 => "1111111001100100111001",
			1597 => "0000001001101000000100",
			1598 => "0000001001100100111001",
			1599 => "0000000001100100111001",
			1600 => "0011110011111100001100",
			1601 => "0011101010001000000100",
			1602 => "1111111001100100111001",
			1603 => "0000100101101000000100",
			1604 => "1111111001100100111001",
			1605 => "0000001001100100111001",
			1606 => "0000001000110000001000",
			1607 => "0001101001111000000100",
			1608 => "0000001001100100111001",
			1609 => "0000000001100100111001",
			1610 => "0000000001100100111001",
			1611 => "0001011001000000000100",
			1612 => "0000000001100100111001",
			1613 => "1111111001100100111001",
			1614 => "0010111010100101001100",
			1615 => "0010010101011100100100",
			1616 => "0001101010111100011100",
			1617 => "0001001010000100011000",
			1618 => "0000001011010000010000",
			1619 => "0010001001001100001000",
			1620 => "0011101001011100000100",
			1621 => "1111111001101001110101",
			1622 => "0000000001101001110101",
			1623 => "0000010111110000000100",
			1624 => "0000001001101001110101",
			1625 => "0000000001101001110101",
			1626 => "0001100100000100000100",
			1627 => "0000001001101001110101",
			1628 => "0000000001101001110101",
			1629 => "0000000001101001110101",
			1630 => "0010000101011100000100",
			1631 => "0000000001101001110101",
			1632 => "1111111001101001110101",
			1633 => "0000100000101000011100",
			1634 => "0011100000110100001100",
			1635 => "0001011100000000001000",
			1636 => "0001010101111000000100",
			1637 => "0000000001101001110101",
			1638 => "0000000001101001110101",
			1639 => "0000000001101001110101",
			1640 => "0011100011101100000100",
			1641 => "1111111001101001110101",
			1642 => "0001100101100000000100",
			1643 => "0000000001101001110101",
			1644 => "0010101111101000000100",
			1645 => "1111111001101001110101",
			1646 => "0000000001101001110101",
			1647 => "0000111100010000000100",
			1648 => "0000000001101001110101",
			1649 => "0001011001010000000100",
			1650 => "1111111001101001110101",
			1651 => "0000000001101001110101",
			1652 => "0011110111010000101100",
			1653 => "0000010001100100100000",
			1654 => "0000010110010000000100",
			1655 => "1111111001101001110101",
			1656 => "0001010110011100010000",
			1657 => "0001111101001000001000",
			1658 => "0011011010100100000100",
			1659 => "0000001001101001110101",
			1660 => "0000000001101001110101",
			1661 => "0010110101010100000100",
			1662 => "0000000001101001110101",
			1663 => "0000000001101001110101",
			1664 => "0010101001000000001000",
			1665 => "0001001011111000000100",
			1666 => "0000001001101001110101",
			1667 => "0000000001101001110101",
			1668 => "0000000001101001110101",
			1669 => "0000111100101100000100",
			1670 => "1111111001101001110101",
			1671 => "0000110011000100000100",
			1672 => "0000000001101001110101",
			1673 => "0000000001101001110101",
			1674 => "0001101110101100010100",
			1675 => "0010110011010000000100",
			1676 => "0000001001101001110101",
			1677 => "0000011001100000000100",
			1678 => "0000000001101001110101",
			1679 => "0011010101010100000100",
			1680 => "0000001001101001110101",
			1681 => "0001011100101100000100",
			1682 => "0000000001101001110101",
			1683 => "0000000001101001110101",
			1684 => "0011110011111100001100",
			1685 => "0010101011000000000100",
			1686 => "1111111001101001110101",
			1687 => "0001101110000100000100",
			1688 => "0000000001101001110101",
			1689 => "0000000001101001110101",
			1690 => "0001000011000000000100",
			1691 => "0000001001101001110101",
			1692 => "0000000001101001110101",
			1693 => "0001111011111001111000",
			1694 => "0010111010100100111100",
			1695 => "0010010101011100100000",
			1696 => "0010111110011000011000",
			1697 => "0001100001100000001100",
			1698 => "0001101110001100000100",
			1699 => "0000000001101110011001",
			1700 => "0000001001110100000100",
			1701 => "0000000001101110011001",
			1702 => "0000000001101110011001",
			1703 => "0001111001010100001000",
			1704 => "0000110011001000000100",
			1705 => "0000000001101110011001",
			1706 => "0000000001101110011001",
			1707 => "0000000001101110011001",
			1708 => "0000000011001100000100",
			1709 => "0000000001101110011001",
			1710 => "0000000001101110011001",
			1711 => "0000100000101000010100",
			1712 => "0001111001010000001100",
			1713 => "0011100000110100001000",
			1714 => "0001100101110100000100",
			1715 => "0000000001101110011001",
			1716 => "0000000001101110011001",
			1717 => "0000000001101110011001",
			1718 => "0001001100101000000100",
			1719 => "0000000001101110011001",
			1720 => "0000000001101110011001",
			1721 => "0000111100010000000100",
			1722 => "0000000001101110011001",
			1723 => "0000000001101110011001",
			1724 => "0010101111101000100000",
			1725 => "0000010001100100011000",
			1726 => "0010101000111000001100",
			1727 => "0011010110001100000100",
			1728 => "0000000001101110011001",
			1729 => "0010110111011100000100",
			1730 => "0000000001101110011001",
			1731 => "0000000001101110011001",
			1732 => "0010110101011100001000",
			1733 => "0000001011001000000100",
			1734 => "0000000001101110011001",
			1735 => "0000001001101110011001",
			1736 => "0000000001101110011001",
			1737 => "0001011101001000000100",
			1738 => "0000000001101110011001",
			1739 => "0000000001101110011001",
			1740 => "0010001001000100001100",
			1741 => "0001001001010000000100",
			1742 => "0000000001101110011001",
			1743 => "0001010010111000000100",
			1744 => "0000000001101110011001",
			1745 => "0000000001101110011001",
			1746 => "0011110111000000001100",
			1747 => "0000011000011000000100",
			1748 => "0000000001101110011001",
			1749 => "0000111100101100000100",
			1750 => "0000000001101110011001",
			1751 => "0000000001101110011001",
			1752 => "0000000001101110011001",
			1753 => "0010101011000000000100",
			1754 => "0000000001101110011001",
			1755 => "0000001111001100001100",
			1756 => "0001010001001000000100",
			1757 => "0000000001101110011001",
			1758 => "0011100100010000000100",
			1759 => "0000000001101110011001",
			1760 => "0000000001101110011001",
			1761 => "0000100101101000000100",
			1762 => "0000000001101110011001",
			1763 => "0000100101010000000100",
			1764 => "0000000001101110011001",
			1765 => "0000000001101110011001",
			1766 => "0001000111110000001100",
			1767 => "0001000001110000000100",
			1768 => "0000000001110001010101",
			1769 => "0000111101000000000100",
			1770 => "0000110001110001010101",
			1771 => "0000000001110001010101",
			1772 => "0010011111011001010000",
			1773 => "0000111000000000100000",
			1774 => "0010001001000100011000",
			1775 => "0001100000001100010000",
			1776 => "0011100011101100001000",
			1777 => "0001100100110000000100",
			1778 => "0000000001110001010101",
			1779 => "0000000001110001010101",
			1780 => "0001111001010000000100",
			1781 => "0000001001110001010101",
			1782 => "0000000001110001010101",
			1783 => "0001000111011100000100",
			1784 => "0000000001110001010101",
			1785 => "1111111001110001010101",
			1786 => "0000110011100100000100",
			1787 => "1111111001110001010101",
			1788 => "0000000001110001010101",
			1789 => "0000101111101100011100",
			1790 => "0011100100001100010000",
			1791 => "0000011000011000001000",
			1792 => "0010001001000100000100",
			1793 => "0000000001110001010101",
			1794 => "0000001001110001010101",
			1795 => "0010101001010100000100",
			1796 => "0000000001110001010101",
			1797 => "1111111001110001010101",
			1798 => "0010101001011000001000",
			1799 => "0001111000101000000100",
			1800 => "1111111001110001010101",
			1801 => "0000000001110001010101",
			1802 => "0000000001110001010101",
			1803 => "0001110110101100000100",
			1804 => "1111111001110001010101",
			1805 => "0001101010111100001000",
			1806 => "0000101011100100000100",
			1807 => "0000001001110001010101",
			1808 => "0000000001110001010101",
			1809 => "0000111000101000000100",
			1810 => "0000000001110001010101",
			1811 => "0000000001110001010101",
			1812 => "1111111001110001010101",
			1813 => "0000100110101001011000",
			1814 => "0000010001100101001100",
			1815 => "0010101000101000110000",
			1816 => "0010101000111000011100",
			1817 => "0011010110001100010000",
			1818 => "0010001001001100001000",
			1819 => "0001111100010000000100",
			1820 => "0000000001110101011001",
			1821 => "0000000001110101011001",
			1822 => "0011110001010100000100",
			1823 => "0000000001110101011001",
			1824 => "0000000001110101011001",
			1825 => "0010001111111100000100",
			1826 => "1111111001110101011001",
			1827 => "0010011100101000000100",
			1828 => "0000000001110101011001",
			1829 => "0000000001110101011001",
			1830 => "0011101111110100001100",
			1831 => "0011011010100100001000",
			1832 => "0011000101010100000100",
			1833 => "0000001001110101011001",
			1834 => "0000000001110101011001",
			1835 => "0000000001110101011001",
			1836 => "0011110000000100000100",
			1837 => "0000000001110101011001",
			1838 => "1111111001110101011001",
			1839 => "0010001111001000010100",
			1840 => "0011111010110000001100",
			1841 => "0011010101010100000100",
			1842 => "1111111001110101011001",
			1843 => "0001011001111100000100",
			1844 => "0000000001110101011001",
			1845 => "0000000001110101011001",
			1846 => "0000000110101000000100",
			1847 => "0000000001110101011001",
			1848 => "0000000001110101011001",
			1849 => "0000101000011100000100",
			1850 => "0000000001110101011001",
			1851 => "0000000001110101011001",
			1852 => "0010101001000000000100",
			1853 => "1111111001110101011001",
			1854 => "0011101110100100000100",
			1855 => "0000000001110101011001",
			1856 => "0000000001110101011001",
			1857 => "0011110101111100000100",
			1858 => "0000001001110101011001",
			1859 => "0011101111110100000100",
			1860 => "0000000001110101011001",
			1861 => "0011010101010100010100",
			1862 => "0001100101001100000100",
			1863 => "0000000001110101011001",
			1864 => "0011001110011000001000",
			1865 => "0001111000101000000100",
			1866 => "1111111001110101011001",
			1867 => "0000000001110101011001",
			1868 => "0001111001010000000100",
			1869 => "0000000001110101011001",
			1870 => "0000000001110101011001",
			1871 => "0000111000000000000100",
			1872 => "1111111001110101011001",
			1873 => "0010000000110000000100",
			1874 => "0000000001110101011001",
			1875 => "0011111100111100000100",
			1876 => "0000000001110101011001",
			1877 => "1111111001110101011001",
			1878 => "0011100100011110000000",
			1879 => "0000001010010101010100",
			1880 => "0001100100000100111100",
			1881 => "0010101000101000100000",
			1882 => "0010101000111000010000",
			1883 => "0001111001010100001000",
			1884 => "0011100010011000000100",
			1885 => "0000000001111001011111",
			1886 => "1111111001111001011111",
			1887 => "0010001001000100000100",
			1888 => "0000001001111001011111",
			1889 => "0000000001111001011111",
			1890 => "0001011100110000001000",
			1891 => "0001111101001000000100",
			1892 => "0000001001111001011111",
			1893 => "0000000001111001011111",
			1894 => "0011011010100100000100",
			1895 => "0000000001111001011111",
			1896 => "0000000001111001011111",
			1897 => "0000011000011000010000",
			1898 => "0010001001000100001000",
			1899 => "0011111010101100000100",
			1900 => "0000000001111001011111",
			1901 => "0000000001111001011111",
			1902 => "0001100111001000000100",
			1903 => "0000000001111001011111",
			1904 => "0000000001111001011111",
			1905 => "0001111000101000000100",
			1906 => "1111111001111001011111",
			1907 => "0000111111101000000100",
			1908 => "0000000001111001011111",
			1909 => "0000000001111001011111",
			1910 => "0010110111011100000100",
			1911 => "1111111001111001011111",
			1912 => "0001001100000000001000",
			1913 => "0001101110001000000100",
			1914 => "0000000001111001011111",
			1915 => "0000000001111001011111",
			1916 => "0011100110110000000100",
			1917 => "0000000001111001011111",
			1918 => "0001001001010100000100",
			1919 => "0000000001111001011111",
			1920 => "0000000001111001011111",
			1921 => "0001101010101100010000",
			1922 => "0000000101101000001100",
			1923 => "0000010111100100001000",
			1924 => "0000100110111100000100",
			1925 => "0000000001111001011111",
			1926 => "0000000001111001011111",
			1927 => "0000001001111001011111",
			1928 => "0000000001111001011111",
			1929 => "0000010001110000000100",
			1930 => "0000000001111001011111",
			1931 => "0001011101001000001000",
			1932 => "0000110011001000000100",
			1933 => "0000000001111001011111",
			1934 => "1111111001111001011111",
			1935 => "0010000000110000001000",
			1936 => "0000011001100000000100",
			1937 => "0000000001111001011111",
			1938 => "0000000001111001011111",
			1939 => "0001001000111000000100",
			1940 => "0000000001111001011111",
			1941 => "0000000001111001011111",
			1942 => "0000000001111001011111",
			1943 => "0011100100011100011100",
			1944 => "0011110001010100000100",
			1945 => "1111111001111010011001",
			1946 => "0010010111011100000100",
			1947 => "0000001001111010011001",
			1948 => "0000110011000000000100",
			1949 => "1111111001111010011001",
			1950 => "0010001010100100000100",
			1951 => "1111111001111010011001",
			1952 => "0001111100000000000100",
			1953 => "1111111001111010011001",
			1954 => "0011111100111100000100",
			1955 => "0000000001111010011001",
			1956 => "0000000001111010011001",
			1957 => "1111111001111010011001",
			1958 => "0011111101100100010000",
			1959 => "0010011010100100000100",
			1960 => "0000000001111011110101",
			1961 => "0011000111011100001000",
			1962 => "0010010110000000000100",
			1963 => "1111111001111011110101",
			1964 => "0000000001111011110101",
			1965 => "1111111001111011110101",
			1966 => "0010011111011000011100",
			1967 => "0011100100011100011000",
			1968 => "0011011111011100000100",
			1969 => "0000001001111011110101",
			1970 => "0001001010100100000100",
			1971 => "1111111001111011110101",
			1972 => "0010111011101100001000",
			1973 => "0001100100000100000100",
			1974 => "0000001001111011110101",
			1975 => "1111111001111011110101",
			1976 => "0000000110111100000100",
			1977 => "0000000001111011110101",
			1978 => "0000001001111011110101",
			1979 => "1111111001111011110101",
			1980 => "1111111001111011110101",
			1981 => "0011100100011100100000",
			1982 => "0011110001010100000100",
			1983 => "0000000001111100111001",
			1984 => "0010010111011100000100",
			1985 => "0000000001111100111001",
			1986 => "0000110011000000000100",
			1987 => "0000000001111100111001",
			1988 => "0010001010100100000100",
			1989 => "0000000001111100111001",
			1990 => "0010101111101000001000",
			1991 => "0000010001100100000100",
			1992 => "0000000001111100111001",
			1993 => "0000000001111100111001",
			1994 => "0000010111110000000100",
			1995 => "1111111001111100111001",
			1996 => "0000000001111100111001",
			1997 => "0000000001111100111001",
			1998 => "0001001100000000101100",
			1999 => "0001001000000100101000",
			2000 => "0010000000110000011000",
			2001 => "0010101011000000010100",
			2002 => "0001010100101100010000",
			2003 => "0011000101010100001000",
			2004 => "0000010001100100000100",
			2005 => "0000000001111111000101",
			2006 => "0000000001111111000101",
			2007 => "0001001100101000000100",
			2008 => "0000000001111111000101",
			2009 => "0000000001111111000101",
			2010 => "0000000001111111000101",
			2011 => "0000001001111111000101",
			2012 => "0001001001001000001100",
			2013 => "0001111111101000000100",
			2014 => "0000000001111111000101",
			2015 => "0001111011111000000100",
			2016 => "0000000001111111000101",
			2017 => "0000000001111111000101",
			2018 => "1111111001111111000101",
			2019 => "0000001001111111000101",
			2020 => "0001001001010000001100",
			2021 => "0010110101010100000100",
			2022 => "1111111001111111000101",
			2023 => "0010111100101000000100",
			2024 => "0000000001111111000101",
			2025 => "1111111001111111000101",
			2026 => "0001000100101100001100",
			2027 => "0011110001100000000100",
			2028 => "0000000001111111000101",
			2029 => "0000111011000000000100",
			2030 => "0000001001111111000101",
			2031 => "0000000001111111000101",
			2032 => "0000000001111111000101",
			2033 => "0000101010000000011000",
			2034 => "0011111101100100010000",
			2035 => "0010011010100100000100",
			2036 => "0000000010000001001001",
			2037 => "0011000111011100001000",
			2038 => "0011000011010000000100",
			2039 => "1111111010000001001001",
			2040 => "1111111010000001001001",
			2041 => "1111111010000001001001",
			2042 => "0001110110101100000100",
			2043 => "0000001010000001001001",
			2044 => "1111111010000001001001",
			2045 => "0010011111011000101000",
			2046 => "0001100111010000100100",
			2047 => "0001101010111100010100",
			2048 => "0010110101010100010000",
			2049 => "0010010101011100001000",
			2050 => "0011111100111100000100",
			2051 => "0000010010000001001001",
			2052 => "0000001010000001001001",
			2053 => "0000100110010100000100",
			2054 => "0000000010000001001001",
			2055 => "0000001010000001001001",
			2056 => "0000010010000001001001",
			2057 => "0000101100100100000100",
			2058 => "1111111010000001001001",
			2059 => "0000010001110000000100",
			2060 => "0000010010000001001001",
			2061 => "0010010101101100000100",
			2062 => "0000000010000001001001",
			2063 => "0000001010000001001001",
			2064 => "1111111010000001001001",
			2065 => "1111111010000001001001",
			2066 => "0000100101011000010100",
			2067 => "0000010111100100000100",
			2068 => "1111111010000011101101",
			2069 => "0011000111011100001100",
			2070 => "0000010011110000001000",
			2071 => "0001111100000000000100",
			2072 => "1111111010000011101101",
			2073 => "0000001010000011101101",
			2074 => "1111111010000011101101",
			2075 => "1111111010000011101101",
			2076 => "0011010101010100110100",
			2077 => "0001101101010000100000",
			2078 => "0011111000001000010100",
			2079 => "0011111011110100010000",
			2080 => "0010010101011100001000",
			2081 => "0010101000000100000100",
			2082 => "0000000010000011101101",
			2083 => "0000001010000011101101",
			2084 => "0000010000011000000100",
			2085 => "1111111010000011101101",
			2086 => "0000000010000011101101",
			2087 => "1111111010000011101101",
			2088 => "0011001010100100000100",
			2089 => "1111111010000011101101",
			2090 => "0011011011101100000100",
			2091 => "0000001010000011101101",
			2092 => "0000001010000011101101",
			2093 => "0000101011001100001100",
			2094 => "0001110100101100000100",
			2095 => "1111111010000011101101",
			2096 => "0011011110011000000100",
			2097 => "0000000010000011101101",
			2098 => "0000000010000011101101",
			2099 => "0011110011111100000100",
			2100 => "0000000010000011101101",
			2101 => "0000001010000011101101",
			2102 => "0011000101011100000100",
			2103 => "1111111010000011101101",
			2104 => "0010010101111000000100",
			2105 => "0000001010000011101101",
			2106 => "1111111010000011101101",
			2107 => "0000100101011000010100",
			2108 => "0000010111100100000100",
			2109 => "1111111010000110000001",
			2110 => "0011000111011100001100",
			2111 => "0000010011110000001000",
			2112 => "0001111100000000000100",
			2113 => "1111111010000110000001",
			2114 => "0000001010000110000001",
			2115 => "1111111010000110000001",
			2116 => "1111111010000110000001",
			2117 => "0011010101010100101100",
			2118 => "0011101111110000000100",
			2119 => "0000001010000110000001",
			2120 => "0000100110010100010000",
			2121 => "0010101111101000001100",
			2122 => "0001101000110100001000",
			2123 => "0001101110010000000100",
			2124 => "0000000010000110000001",
			2125 => "0000000010000110000001",
			2126 => "1111111010000110000001",
			2127 => "1111111010000110000001",
			2128 => "0001110110101100001000",
			2129 => "0011001110011000000100",
			2130 => "0000000010000110000001",
			2131 => "1111111010000110000001",
			2132 => "0001101101010000001000",
			2133 => "0011101110100100000100",
			2134 => "0000000010000110000001",
			2135 => "0000001010000110000001",
			2136 => "0000001110101000000100",
			2137 => "1111111010000110000001",
			2138 => "0000000010000110000001",
			2139 => "0011000101011100000100",
			2140 => "1111111010000110000001",
			2141 => "0010010101111000000100",
			2142 => "0000001010000110000001",
			2143 => "1111111010000110000001",
			2144 => "0001000111110000001100",
			2145 => "0001000001110000000100",
			2146 => "0000000010000111110101",
			2147 => "0010011001000100000100",
			2148 => "0000001010000111110101",
			2149 => "0000000010000111110101",
			2150 => "0010101110111000101100",
			2151 => "0011100010001100000100",
			2152 => "1111111010000111110101",
			2153 => "0011100010000000010000",
			2154 => "0000001001110100001100",
			2155 => "0011001010100100000100",
			2156 => "1111111010000111110101",
			2157 => "0011011010100100000100",
			2158 => "0000001010000111110101",
			2159 => "0000000010000111110101",
			2160 => "0000001010000111110101",
			2161 => "0011100001101100001000",
			2162 => "0011001010100100000100",
			2163 => "0000000010000111110101",
			2164 => "1111111010000111110101",
			2165 => "0010111110011000001000",
			2166 => "0000110011100100000100",
			2167 => "0000000010000111110101",
			2168 => "1111111010000111110101",
			2169 => "0001111001010100000100",
			2170 => "0000000010000111110101",
			2171 => "0000000010000111110101",
			2172 => "1111111010000111110101",
			2173 => "0000101011101000010100",
			2174 => "0011011110011000000100",
			2175 => "1111111010001010000001",
			2176 => "0011000111011100001100",
			2177 => "0010001111001000001000",
			2178 => "0001111100000000000100",
			2179 => "0000000010001010000001",
			2180 => "0000001010001010000001",
			2181 => "1111111010001010000001",
			2182 => "1111111010001010000001",
			2183 => "0001110011000100110000",
			2184 => "0010110101010100100000",
			2185 => "0010000000110000011100",
			2186 => "0011111011011100001100",
			2187 => "0000010111100100001000",
			2188 => "0011001010100100000100",
			2189 => "0000000010001010000001",
			2190 => "0000001010001010000001",
			2191 => "0000000010001010000001",
			2192 => "0000100110010100001000",
			2193 => "0000111000000000000100",
			2194 => "0000000010001010000001",
			2195 => "1111111010001010000001",
			2196 => "0001011001010000000100",
			2197 => "0000000010001010000001",
			2198 => "0000000010001010000001",
			2199 => "1111111010001010000001",
			2200 => "0000011110011000001100",
			2201 => "0001011100101100000100",
			2202 => "0000000010001010000001",
			2203 => "0001001001010100000100",
			2204 => "0000001010001010000001",
			2205 => "1111111010001010000001",
			2206 => "1111111010001010000001",
			2207 => "1111111010001010000001",
			2208 => "0010011010100100000100",
			2209 => "0000001010001011010101",
			2210 => "0000110011000000000100",
			2211 => "1111111010001011010101",
			2212 => "0001000100101100100000",
			2213 => "0000011011101100011100",
			2214 => "0001100000001100010000",
			2215 => "0010010101011100001000",
			2216 => "0000001110110000000100",
			2217 => "0000001010001011010101",
			2218 => "1111111010001011010101",
			2219 => "0000010110010000000100",
			2220 => "0000000010001011010101",
			2221 => "0000000010001011010101",
			2222 => "0000001111001100000100",
			2223 => "1111111010001011010101",
			2224 => "0011110011111100000100",
			2225 => "0000000010001011010101",
			2226 => "0000001010001011010101",
			2227 => "1111111010001011010101",
			2228 => "1111111010001011010101",
			2229 => "0000001011111100011000",
			2230 => "0011111101100100010000",
			2231 => "0010011010100100000100",
			2232 => "0000000010001101101001",
			2233 => "0011000111011100001000",
			2234 => "0011000011010000000100",
			2235 => "1111111010001101101001",
			2236 => "1111111010001101101001",
			2237 => "1111111010001101101001",
			2238 => "0001111101001000000100",
			2239 => "0000010010001101101001",
			2240 => "1111111010001101101001",
			2241 => "0010011111011000110000",
			2242 => "0011100100011100101100",
			2243 => "0011000101010100011100",
			2244 => "0000111101001000010000",
			2245 => "0000101101110000001000",
			2246 => "0010101111011000000100",
			2247 => "0000000010001101101001",
			2248 => "0000011010001101101001",
			2249 => "0011101101100100000100",
			2250 => "0000000010001101101001",
			2251 => "0000011010001101101001",
			2252 => "0001001100000000001000",
			2253 => "0011101101100000000100",
			2254 => "0000011010001101101001",
			2255 => "0000000010001101101001",
			2256 => "1111111010001101101001",
			2257 => "0010001111011000001100",
			2258 => "0000100011001100000100",
			2259 => "0000010010001101101001",
			2260 => "0000011001100000000100",
			2261 => "0000011010001101101001",
			2262 => "0000101010001101101001",
			2263 => "0000001010001101101001",
			2264 => "1111111010001101101001",
			2265 => "1111111010001101101001",
			2266 => "0000000011111000000100",
			2267 => "0000000010010000001101",
			2268 => "0010101111101000101000",
			2269 => "0011010101010100100000",
			2270 => "0001111101001000010100",
			2271 => "0001100100000100001000",
			2272 => "0010101000111000000100",
			2273 => "0000000010010000001101",
			2274 => "0000000010010000001101",
			2275 => "0000110011100100001000",
			2276 => "0011111011010100000100",
			2277 => "0000000010010000001101",
			2278 => "0000000010010000001101",
			2279 => "0000000010010000001101",
			2280 => "0011110100110100000100",
			2281 => "0000000010010000001101",
			2282 => "0011110011111100000100",
			2283 => "0000000010010000001101",
			2284 => "0000000010010000001101",
			2285 => "0000001011001100000100",
			2286 => "0000000010010000001101",
			2287 => "0000000010010000001101",
			2288 => "0010110101010100010100",
			2289 => "0011111011000100001100",
			2290 => "0011101101100000001000",
			2291 => "0011100011011000000100",
			2292 => "0000000010010000001101",
			2293 => "0000000010010000001101",
			2294 => "0000000010010000001101",
			2295 => "0011100011101000000100",
			2296 => "0000000010010000001101",
			2297 => "0000000010010000001101",
			2298 => "0011011100101000001000",
			2299 => "0011100100101000000100",
			2300 => "0000000010010000001101",
			2301 => "0000000010010000001101",
			2302 => "0001001111011000001000",
			2303 => "0000000101101000000100",
			2304 => "0000000010010000001101",
			2305 => "0000000010010000001101",
			2306 => "0000000010010000001101",
			2307 => "0000101000011100010000",
			2308 => "0011000111011100001100",
			2309 => "0011000011010000000100",
			2310 => "1111111010010010100001",
			2311 => "0000010111100100000100",
			2312 => "1111111010010010100001",
			2313 => "0000001010010010100001",
			2314 => "1111111010010010100001",
			2315 => "0011011001001000110100",
			2316 => "0010101110111000110000",
			2317 => "0011111100111100010100",
			2318 => "0000100110101000001100",
			2319 => "0000010001100100001000",
			2320 => "0010001111111100000100",
			2321 => "0000000010010010100001",
			2322 => "0000001010010010100001",
			2323 => "1111111010010010100001",
			2324 => "0000010110010000000100",
			2325 => "0000000010010010100001",
			2326 => "0000001010010010100001",
			2327 => "0000100000101000010000",
			2328 => "0010111010100100001000",
			2329 => "0000110011100100000100",
			2330 => "0000000010010010100001",
			2331 => "1111111010010010100001",
			2332 => "0010001111001000000100",
			2333 => "0000001010010010100001",
			2334 => "1111111010010010100001",
			2335 => "0000000101101000000100",
			2336 => "0000001010010010100001",
			2337 => "0011111011000100000100",
			2338 => "1111111010010010100001",
			2339 => "0000000010010010100001",
			2340 => "1111111010010010100001",
			2341 => "0000010110001100000100",
			2342 => "0000000010010010100001",
			2343 => "1111111010010010100001",
			2344 => "0011111101100100010100",
			2345 => "0010011010100100000100",
			2346 => "0000001010010101000101",
			2347 => "0011000111011100001100",
			2348 => "0010001001000100000100",
			2349 => "1111111010010101000101",
			2350 => "0011011010100100000100",
			2351 => "0000010010010101000101",
			2352 => "1111111010010101000101",
			2353 => "1111111010010101000101",
			2354 => "0010001111011000111000",
			2355 => "0000111011000000110000",
			2356 => "0011000101010100011100",
			2357 => "0010101000101000010000",
			2358 => "0001100100000100001000",
			2359 => "0010100011000000000100",
			2360 => "0000000010010101000101",
			2361 => "0000001010010101000101",
			2362 => "0000001010010100000100",
			2363 => "1111111010010101000101",
			2364 => "0000000010010101000101",
			2365 => "0000101111101100000100",
			2366 => "1111111010010101000101",
			2367 => "0010101011111000000100",
			2368 => "0000000010010101000101",
			2369 => "1111111010010101000101",
			2370 => "0000000110111100001000",
			2371 => "0001011000101000000100",
			2372 => "1111111010010101000101",
			2373 => "0000000010010101000101",
			2374 => "0000011001100000000100",
			2375 => "0000000010010101000101",
			2376 => "0011110101100100000100",
			2377 => "0000001010010101000101",
			2378 => "0000001010010101000101",
			2379 => "0010001001000100000100",
			2380 => "1111111010010101000101",
			2381 => "0000000010010101000101",
			2382 => "0000010110001100000100",
			2383 => "0000000010010101000101",
			2384 => "1111111010010101000101",
			2385 => "0001001100000000110000",
			2386 => "0001001000000100101100",
			2387 => "0010001111011000101000",
			2388 => "0001101101010000011000",
			2389 => "0010001010100100001000",
			2390 => "0010010111011100000100",
			2391 => "0000000010010111111001",
			2392 => "1111111010010111111001",
			2393 => "0011111101001100001000",
			2394 => "0000010001100100000100",
			2395 => "0000000010010111111001",
			2396 => "0000000010010111111001",
			2397 => "0011001010100100000100",
			2398 => "1111111010010111111001",
			2399 => "0000001010010111111001",
			2400 => "0000010110010000000100",
			2401 => "0000000010010111111001",
			2402 => "0000001010111000000100",
			2403 => "1111111010010111111001",
			2404 => "0001011100110000000100",
			2405 => "0000000010010111111001",
			2406 => "0000000010010111111001",
			2407 => "1111111010010111111001",
			2408 => "0000001010010111111001",
			2409 => "0001000110101100010100",
			2410 => "0010110101010100001000",
			2411 => "0001011100101100000100",
			2412 => "0000000010010111111001",
			2413 => "1111111010010111111001",
			2414 => "0001011000100000000100",
			2415 => "1111111010010111111001",
			2416 => "0001010001001000000100",
			2417 => "0000001010010111111001",
			2418 => "0000000010010111111001",
			2419 => "0011110001100000000100",
			2420 => "1111111010010111111001",
			2421 => "0010101001000000010000",
			2422 => "0001011010011100001100",
			2423 => "0000000000000000000100",
			2424 => "1111111010010111111001",
			2425 => "0001001000101000000100",
			2426 => "0000001010010111111001",
			2427 => "0000000010010111111001",
			2428 => "0000001010010111111001",
			2429 => "1111111010010111111001",
			2430 => "0000001001110100011100",
			2431 => "0001000111110000001000",
			2432 => "0001101011111000000100",
			2433 => "0000000010011010100101",
			2434 => "0000000010011010100101",
			2435 => "0001100001100000001100",
			2436 => "0001011010011100000100",
			2437 => "0000000010011010100101",
			2438 => "0001011110001100000100",
			2439 => "0000000010011010100101",
			2440 => "0000000010011010100101",
			2441 => "0000001010000000000100",
			2442 => "0000000010011010100101",
			2443 => "0000000010011010100101",
			2444 => "0011100010000000000100",
			2445 => "0000000010011010100101",
			2446 => "0001110110101100001000",
			2447 => "0000010110010000000100",
			2448 => "0000000010011010100101",
			2449 => "0000000010011010100101",
			2450 => "0011010011010000011100",
			2451 => "0010101111101000010000",
			2452 => "0010111010100100001000",
			2453 => "0000001111001100000100",
			2454 => "0000000010011010100101",
			2455 => "0000000010011010100101",
			2456 => "0000000101101000000100",
			2457 => "0000000010011010100101",
			2458 => "0000000010011010100101",
			2459 => "0000010111110000000100",
			2460 => "0000000010011010100101",
			2461 => "0000100011001100000100",
			2462 => "0000000010011010100101",
			2463 => "0000000010011010100101",
			2464 => "0010101000101000000100",
			2465 => "0000000010011010100101",
			2466 => "0010001111011000001000",
			2467 => "0001001100000000000100",
			2468 => "0000000010011010100101",
			2469 => "0000000010011010100101",
			2470 => "0000111011000000000100",
			2471 => "0000000010011010100101",
			2472 => "0000000010011010100101",
			2473 => "0000111011000000110100",
			2474 => "0010011010100100001000",
			2475 => "0000001010011000000100",
			2476 => "1111111010011100010001",
			2477 => "0000010010011100010001",
			2478 => "0000110011000000000100",
			2479 => "1111111010011100010001",
			2480 => "0010001111011000100000",
			2481 => "0010110111011100010000",
			2482 => "0010010110000000001000",
			2483 => "0011000101010100000100",
			2484 => "0000000010011100010001",
			2485 => "0000001010011100010001",
			2486 => "0000011001100000000100",
			2487 => "0000000010011100010001",
			2488 => "1111111010011100010001",
			2489 => "0000010110010000001000",
			2490 => "0001010110101100000100",
			2491 => "0000001010011100010001",
			2492 => "1111111010011100010001",
			2493 => "0001011101001000000100",
			2494 => "0000000010011100010001",
			2495 => "0000001010011100010001",
			2496 => "0001110100101100000100",
			2497 => "0000000010011100010001",
			2498 => "1111111010011100010001",
			2499 => "1111111010011100010001",
			2500 => "0000100101011000010100",
			2501 => "0010011010100100000100",
			2502 => "0000000010011110101101",
			2503 => "0011000111011100001100",
			2504 => "0010110111011100001000",
			2505 => "0000100100111100000100",
			2506 => "1111111010011110101101",
			2507 => "0000000010011110101101",
			2508 => "0000001010011110101101",
			2509 => "1111111010011110101101",
			2510 => "0010011111011000111000",
			2511 => "0011100010110100110000",
			2512 => "0000100110010100011000",
			2513 => "0001100100110000010000",
			2514 => "0010101111101000001000",
			2515 => "0011001010100100000100",
			2516 => "0000001010011110101101",
			2517 => "0000010010011110101101",
			2518 => "0001000110101100000100",
			2519 => "1111111010011110101101",
			2520 => "0000001010011110101101",
			2521 => "0001111000101000000100",
			2522 => "1111111010011110101101",
			2523 => "0000000010011110101101",
			2524 => "0001110110101100001000",
			2525 => "0010001001001100000100",
			2526 => "0000001010011110101101",
			2527 => "1111111010011110101101",
			2528 => "0000000101101000001000",
			2529 => "0000110011100100000100",
			2530 => "0000001010011110101101",
			2531 => "0000010010011110101101",
			2532 => "0011111101001100000100",
			2533 => "0000000010011110101101",
			2534 => "0000001010011110101101",
			2535 => "0011110101100100000100",
			2536 => "0000000010011110101101",
			2537 => "1111111010011110101101",
			2538 => "1111111010011110101101",
			2539 => "0001000111110000001000",
			2540 => "0001101011000000000100",
			2541 => "1111111010100001011001",
			2542 => "0000100010100001011001",
			2543 => "0000101011101000011000",
			2544 => "0000010111100100000100",
			2545 => "1111111010100001011001",
			2546 => "0011000111011100010000",
			2547 => "0000011000011000000100",
			2548 => "0000001010100001011001",
			2549 => "0010000101101100001000",
			2550 => "0001011111011000000100",
			2551 => "1111111010100001011001",
			2552 => "0000001010100001011001",
			2553 => "1111111010100001011001",
			2554 => "1111111010100001011001",
			2555 => "0010010101011100010100",
			2556 => "0001100111101000001000",
			2557 => "0000111111011000000100",
			2558 => "0000000010100001011001",
			2559 => "0000001010100001011001",
			2560 => "0011001010100100001000",
			2561 => "0001000101010100000100",
			2562 => "0000000010100001011001",
			2563 => "1111111010100001011001",
			2564 => "0000000010100001011001",
			2565 => "0010000101011100010000",
			2566 => "0001111101001000001000",
			2567 => "0011110000001000000100",
			2568 => "0000000010100001011001",
			2569 => "1111111010100001011001",
			2570 => "0001011100110000000100",
			2571 => "0000000010100001011001",
			2572 => "0000000010100001011001",
			2573 => "0000011110011000010000",
			2574 => "0000000110111100001000",
			2575 => "0000100011111000000100",
			2576 => "0000000010100001011001",
			2577 => "1111111010100001011001",
			2578 => "0000110011100100000100",
			2579 => "0000000010100001011001",
			2580 => "0000000010100001011001",
			2581 => "1111111010100001011001",
			2582 => "0001001100000001010100",
			2583 => "0001011001010000111100",
			2584 => "0000010001100100110000",
			2585 => "0001000101101100011100",
			2586 => "0011000011010000010000",
			2587 => "0011010110001100001000",
			2588 => "0000010111110000000100",
			2589 => "0000000010100101000101",
			2590 => "0000000010100101000101",
			2591 => "0011100000110100000100",
			2592 => "0000000010100101000101",
			2593 => "1111111010100101000101",
			2594 => "0001001100101000001000",
			2595 => "0001011000000100000100",
			2596 => "0000000010100101000101",
			2597 => "0000000010100101000101",
			2598 => "0000001010100101000101",
			2599 => "0000011000011000010000",
			2600 => "0001000110000000001000",
			2601 => "0010111010100100000100",
			2602 => "1111111010100101000101",
			2603 => "0000000010100101000101",
			2604 => "0010000101011100000100",
			2605 => "0000000010100101000101",
			2606 => "0000000010100101000101",
			2607 => "0000000010100101000101",
			2608 => "0000111000000000000100",
			2609 => "1111111010100101000101",
			2610 => "0011110000001000000100",
			2611 => "0000000010100101000101",
			2612 => "0000000010100101000101",
			2613 => "0010001111011000010100",
			2614 => "0010000101101100001000",
			2615 => "0011110101111100000100",
			2616 => "0000000010100101000101",
			2617 => "1111111010100101000101",
			2618 => "0000000010101100000100",
			2619 => "0000000010100101000101",
			2620 => "0001111011111000000100",
			2621 => "0000001010100101000101",
			2622 => "0000000010100101000101",
			2623 => "0000000010100101000101",
			2624 => "0001000110101100001100",
			2625 => "0001011000100000000100",
			2626 => "0000000010100101000101",
			2627 => "0001010001001000000100",
			2628 => "0000000010100101000101",
			2629 => "0000000010100101000101",
			2630 => "0000000000000000001100",
			2631 => "0000010111100100001000",
			2632 => "0000010110010000000100",
			2633 => "0000000010100101000101",
			2634 => "0000000010100101000101",
			2635 => "0000000010100101000101",
			2636 => "0001001000101000001000",
			2637 => "0001100010000100000100",
			2638 => "0000000010100101000101",
			2639 => "0000000010100101000101",
			2640 => "0000000010100101000101",
			2641 => "0010001111011001011000",
			2642 => "0010111010100100100000",
			2643 => "0001100000001100010100",
			2644 => "0001011111101000010000",
			2645 => "0000101101110000001100",
			2646 => "0001101110001000001000",
			2647 => "0011001110011000000100",
			2648 => "0000000010101000001001",
			2649 => "0000000010101000001001",
			2650 => "0000000010101000001001",
			2651 => "0000000010101000001001",
			2652 => "1111111010101000001001",
			2653 => "0001101110000100000100",
			2654 => "1111111010101000001001",
			2655 => "0011010110001100000100",
			2656 => "0000000010101000001001",
			2657 => "1111111010101000001001",
			2658 => "0000100011001100100100",
			2659 => "0000010001100100011000",
			2660 => "0000010110010000001000",
			2661 => "0010011001001000000100",
			2662 => "0000000010101000001001",
			2663 => "1111111010101000001001",
			2664 => "0001111001010100001000",
			2665 => "0000100100111100000100",
			2666 => "0000000010101000001001",
			2667 => "0000001010101000001001",
			2668 => "0001111000101000000100",
			2669 => "1111111010101000001001",
			2670 => "0000000010101000001001",
			2671 => "0010101001000000000100",
			2672 => "1111111010101000001001",
			2673 => "0011011001001000000100",
			2674 => "0000000010101000001001",
			2675 => "0000000010101000001001",
			2676 => "0000111000000000000100",
			2677 => "0000000010101000001001",
			2678 => "0010101111101000000100",
			2679 => "0000001010101000001001",
			2680 => "0000011001100000000100",
			2681 => "0000000010101000001001",
			2682 => "0010001010000100000100",
			2683 => "0000001010101000001001",
			2684 => "0000000010101000001001",
			2685 => "0011000101101100000100",
			2686 => "1111111010101000001001",
			2687 => "0011011001001000000100",
			2688 => "0000001010101000001001",
			2689 => "0000000010101000001001",
			2690 => "0000100110010100111000",
			2691 => "0000010001100100101000",
			2692 => "0010101111101000011000",
			2693 => "0001100100110000010100",
			2694 => "0000001011111100001100",
			2695 => "0001111100010000001000",
			2696 => "0010001001001100000100",
			2697 => "1111111010101011101101",
			2698 => "0000000010101011101101",
			2699 => "1111111010101011101101",
			2700 => "0010101000111000000100",
			2701 => "0000000010101011101101",
			2702 => "0000001010101011101101",
			2703 => "0000000010101011101101",
			2704 => "0010011101101000000100",
			2705 => "1111111010101011101101",
			2706 => "0010001111001000000100",
			2707 => "0000000010101011101101",
			2708 => "0000100111001100000100",
			2709 => "0000000010101011101101",
			2710 => "0000000010101011101101",
			2711 => "0000011111001000001100",
			2712 => "0010101001000000000100",
			2713 => "1111111010101011101101",
			2714 => "0001100110000100000100",
			2715 => "0000000010101011101101",
			2716 => "0000000010101011101101",
			2717 => "0000000010101011101101",
			2718 => "0001111001011000110000",
			2719 => "0000000101101000011000",
			2720 => "0000110011001000000100",
			2721 => "0000000010101011101101",
			2722 => "0001110110101100000100",
			2723 => "0000000010101011101101",
			2724 => "0001101010111100001000",
			2725 => "0001010011000100000100",
			2726 => "0000001010101011101101",
			2727 => "0000000010101011101101",
			2728 => "0001011100010000000100",
			2729 => "0000000010101011101101",
			2730 => "0000000010101011101101",
			2731 => "0011110011111100010100",
			2732 => "0001101110101100010000",
			2733 => "0011111101001100001000",
			2734 => "0001111101001000000100",
			2735 => "0000000010101011101101",
			2736 => "1111111010101011101101",
			2737 => "0011010110001100000100",
			2738 => "1111111010101011101101",
			2739 => "0000000010101011101101",
			2740 => "0000000010101011101101",
			2741 => "0000000010101011101101",
			2742 => "0000100101101000000100",
			2743 => "1111111010101011101101",
			2744 => "0000001010010000000100",
			2745 => "0000000010101011101101",
			2746 => "0000000010101011101101",
			2747 => "0000010001110000100000",
			2748 => "0011100011101100011000",
			2749 => "0011001110011000001000",
			2750 => "0000001001110100000100",
			2751 => "0000000010101111011001",
			2752 => "0000000010101111011001",
			2753 => "0000010000011000001100",
			2754 => "0001111000111000001000",
			2755 => "0000101101010000000100",
			2756 => "0000000010101111011001",
			2757 => "0000000010101111011001",
			2758 => "1111111010101111011001",
			2759 => "0000000010101111011001",
			2760 => "0001011001010100000100",
			2761 => "0000000010101111011001",
			2762 => "0000000010101111011001",
			2763 => "0001101101010001000000",
			2764 => "0000010111100100011100",
			2765 => "0001111001010100011000",
			2766 => "0001011100000000001000",
			2767 => "0011110001010100000100",
			2768 => "0000000010101111011001",
			2769 => "0000000010101111011001",
			2770 => "0010000101011100001000",
			2771 => "0001111100010000000100",
			2772 => "0000000010101111011001",
			2773 => "0000000010101111011001",
			2774 => "0010000101101100000100",
			2775 => "0000000010101111011001",
			2776 => "0000000010101111011001",
			2777 => "1111111010101111011001",
			2778 => "0000001011100100011000",
			2779 => "0000010001100100001100",
			2780 => "0001001100000000001000",
			2781 => "0011000011010000000100",
			2782 => "0000000010101111011001",
			2783 => "0000000010101111011001",
			2784 => "0000000010101111011001",
			2785 => "0000011001000100001000",
			2786 => "0011100110110000000100",
			2787 => "0000000010101111011001",
			2788 => "0000000010101111011001",
			2789 => "0000000010101111011001",
			2790 => "0000011110011000001000",
			2791 => "0001011001010000000100",
			2792 => "0000000010101111011001",
			2793 => "0000000010101111011001",
			2794 => "0000000010101111011001",
			2795 => "0010101011000000010000",
			2796 => "0011010110001100000100",
			2797 => "0000000010101111011001",
			2798 => "0000010110001100000100",
			2799 => "1111111010101111011001",
			2800 => "0000011010100100000100",
			2801 => "0000000010101111011001",
			2802 => "0000000010101111011001",
			2803 => "0001010011000100000100",
			2804 => "0000000010101111011001",
			2805 => "0000000010101111011001",
			2806 => "0001001111011001001000",
			2807 => "0000010001100100110000",
			2808 => "0000110011000000001000",
			2809 => "0010011010100100000100",
			2810 => "0000000010110010111101",
			2811 => "0000000010110010111101",
			2812 => "0001000101010100010000",
			2813 => "0001001010100100001000",
			2814 => "0011100100111000000100",
			2815 => "0000000010110010111101",
			2816 => "0000000010110010111101",
			2817 => "0000001010101000000100",
			2818 => "0000000010110010111101",
			2819 => "0000000010110010111101",
			2820 => "0001001100101000001000",
			2821 => "0001011100000000000100",
			2822 => "0000000010110010111101",
			2823 => "0000000010110010111101",
			2824 => "0000011000011000001000",
			2825 => "0000010001110000000100",
			2826 => "0000000010110010111101",
			2827 => "0000000010110010111101",
			2828 => "0001100001100000000100",
			2829 => "0000000010110010111101",
			2830 => "0000000010110010111101",
			2831 => "0001011001010100001000",
			2832 => "0001111101101000000100",
			2833 => "0000000010110010111101",
			2834 => "0000000010110010111101",
			2835 => "0000001101111000000100",
			2836 => "0000000010110010111101",
			2837 => "0000001101011000001000",
			2838 => "0011100001000000000100",
			2839 => "0000000010110010111101",
			2840 => "0000000010110010111101",
			2841 => "0000000010110010111101",
			2842 => "0001001000000100001000",
			2843 => "0001110100101100000100",
			2844 => "0000000010110010111101",
			2845 => "0000000010110010111101",
			2846 => "0001001100000000000100",
			2847 => "0000000010110010111101",
			2848 => "0001000110101100010000",
			2849 => "0000111100101100001100",
			2850 => "0011110000100100000100",
			2851 => "0000000010110010111101",
			2852 => "0011110000101100000100",
			2853 => "0000000010110010111101",
			2854 => "0000000010110010111101",
			2855 => "0000000010110010111101",
			2856 => "0001000100101100001100",
			2857 => "0011000101010100000100",
			2858 => "0000000010110010111101",
			2859 => "0000101000011100000100",
			2860 => "0000000010110010111101",
			2861 => "0000000010110010111101",
			2862 => "0000000010110010111101",
			2863 => "0010010101011100011100",
			2864 => "0011111001111000010100",
			2865 => "0000001011010000001100",
			2866 => "0010101000000100001000",
			2867 => "0001000111110000000100",
			2868 => "0000000010110110110001",
			2869 => "0000000010110110110001",
			2870 => "0000000010110110110001",
			2871 => "0001001101101000000100",
			2872 => "0000000010110110110001",
			2873 => "0000000010110110110001",
			2874 => "0011001110011000000100",
			2875 => "0000000010110110110001",
			2876 => "0000000010110110110001",
			2877 => "0000001010010100110000",
			2878 => "0000100011111000100100",
			2879 => "0011110010010000011100",
			2880 => "0011101001011100001100",
			2881 => "0011111101100100001000",
			2882 => "0000001111010100000100",
			2883 => "0000000010110110110001",
			2884 => "0000000010110110110001",
			2885 => "0000000010110110110001",
			2886 => "0001000101111000001000",
			2887 => "0001000101010100000100",
			2888 => "0000000010110110110001",
			2889 => "0000000010110110110001",
			2890 => "0011100000110100000100",
			2891 => "0000000010110110110001",
			2892 => "0000000010110110110001",
			2893 => "0000000011111000000100",
			2894 => "0000000010110110110001",
			2895 => "0000000010110110110001",
			2896 => "0010110101010100000100",
			2897 => "0000000010110110110001",
			2898 => "0011110101111100000100",
			2899 => "0000000010110110110001",
			2900 => "0000000010110110110001",
			2901 => "0001101010101100001100",
			2902 => "0010000101011100000100",
			2903 => "0000000010110110110001",
			2904 => "0001011001011000000100",
			2905 => "0000000010110110110001",
			2906 => "0000000010110110110001",
			2907 => "0000111000000000001000",
			2908 => "0001110001010000000100",
			2909 => "0000000010110110110001",
			2910 => "0000000010110110110001",
			2911 => "0000111001010100001100",
			2912 => "0010110101011100000100",
			2913 => "0000000010110110110001",
			2914 => "0001011100101100000100",
			2915 => "0000000010110110110001",
			2916 => "0000000010110110110001",
			2917 => "0000001111001100001000",
			2918 => "0010100011000100000100",
			2919 => "0000000010110110110001",
			2920 => "0000000010110110110001",
			2921 => "0000101101111000000100",
			2922 => "0000000010110110110001",
			2923 => "0000000010110110110001",
			2924 => "0011100011101001001000",
			2925 => "0000001010010001000100",
			2926 => "0001101010111100110000",
			2927 => "0011101100011000011100",
			2928 => "0010010101011100001100",
			2929 => "0001101110001100000100",
			2930 => "0000000010111001100101",
			2931 => "0001001010000100000100",
			2932 => "0000000010111001100101",
			2933 => "0000000010111001100101",
			2934 => "0000110011001000001000",
			2935 => "0011010110110100000100",
			2936 => "0000000010111001100101",
			2937 => "1111111010111001100101",
			2938 => "0000010000011000000100",
			2939 => "1111111010111001100101",
			2940 => "0000000010111001100101",
			2941 => "0011110111010000001100",
			2942 => "0001111001011000000100",
			2943 => "0000000010111001100101",
			2944 => "0010101000100000000100",
			2945 => "0000000010111001100101",
			2946 => "0000000010111001100101",
			2947 => "0001011000100000000100",
			2948 => "0000001010111001100101",
			2949 => "0000000010111001100101",
			2950 => "0000101100100100000100",
			2951 => "1111111010111001100101",
			2952 => "0010011100101000000100",
			2953 => "0000000010111001100101",
			2954 => "0011111101001100000100",
			2955 => "0000000010111001100101",
			2956 => "0000001001101000000100",
			2957 => "0000000010111001100101",
			2958 => "0000000010111001100101",
			2959 => "0000000010111001100101",
			2960 => "0011001100101000001000",
			2961 => "0001010101111000000100",
			2962 => "0000000010111001100101",
			2963 => "1111111010111001100101",
			2964 => "0001001100000000001000",
			2965 => "0000100101101000000100",
			2966 => "0000000010111001100101",
			2967 => "0000000010111001100101",
			2968 => "0000000010111001100101",
			2969 => "0001101101010001010000",
			2970 => "0011111000001001000000",
			2971 => "0011111100111100101100",
			2972 => "0000101111101100100000",
			2973 => "0000010001100100010000",
			2974 => "0010101111101000001000",
			2975 => "0011110001010100000100",
			2976 => "1111111010111101000001",
			2977 => "0000000010111101000001",
			2978 => "0001011010011100000100",
			2979 => "1111111010111101000001",
			2980 => "0000000010111101000001",
			2981 => "0000111100101100001000",
			2982 => "0000011100101000000100",
			2983 => "1111111010111101000001",
			2984 => "0000000010111101000001",
			2985 => "0001011110111000000100",
			2986 => "0000000010111101000001",
			2987 => "0000000010111101000001",
			2988 => "0000010110010000000100",
			2989 => "0000000010111101000001",
			2990 => "0011011100101000000100",
			2991 => "0000001010111101000001",
			2992 => "0000000010111101000001",
			2993 => "0011010110110100000100",
			2994 => "0000000010111101000001",
			2995 => "0000010111100100000100",
			2996 => "1111111010111101000001",
			2997 => "0000100000101000001000",
			2998 => "0001001000000000000100",
			2999 => "1111111010111101000001",
			3000 => "0000000010111101000001",
			3001 => "0000001010111101000001",
			3002 => "0011001010100100000100",
			3003 => "1111111010111101000001",
			3004 => "0010011101101000001000",
			3005 => "0011011011101100000100",
			3006 => "0000000010111101000001",
			3007 => "0000001010111101000001",
			3008 => "0000000010111101000001",
			3009 => "0000010110010000000100",
			3010 => "0000000010111101000001",
			3011 => "0011000101010100001000",
			3012 => "0011110111001100000100",
			3013 => "1111111010111101000001",
			3014 => "0000000010111101000001",
			3015 => "0010100100101100001000",
			3016 => "0000001010111000000100",
			3017 => "0000000010111101000001",
			3018 => "0000000010111101000001",
			3019 => "0000111011111000000100",
			3020 => "1111111010111101000001",
			3021 => "0000111100101100000100",
			3022 => "0000000010111101000001",
			3023 => "0000000010111101000001",
			3024 => "0000001011001000100100",
			3025 => "0001000111110000001100",
			3026 => "0001000001110000000100",
			3027 => "0000000011000000110101",
			3028 => "0001100011001000000100",
			3029 => "0000000011000000110101",
			3030 => "0000000011000000110101",
			3031 => "0010011101101000001000",
			3032 => "0011010111011100000100",
			3033 => "0000000011000000110101",
			3034 => "0000000011000000110101",
			3035 => "0011011010100100001100",
			3036 => "0010011010000100001000",
			3037 => "0010110111011100000100",
			3038 => "0000000011000000110101",
			3039 => "0000000011000000110101",
			3040 => "0000000011000000110101",
			3041 => "0000000011000000110101",
			3042 => "0001101010101100111000",
			3043 => "0001110110101100010000",
			3044 => "0001100010110100000100",
			3045 => "0000000011000000110101",
			3046 => "0011001110011000001000",
			3047 => "0000010001110000000100",
			3048 => "0000000011000000110101",
			3049 => "0000000011000000110101",
			3050 => "0000000011000000110101",
			3051 => "0010001111001000010000",
			3052 => "0001001010000100000100",
			3053 => "0000000011000000110101",
			3054 => "0000100000101000001000",
			3055 => "0000000010100100000100",
			3056 => "0000000011000000110101",
			3057 => "0000000011000000110101",
			3058 => "0000000011000000110101",
			3059 => "0011100111001000001100",
			3060 => "0011101111110100001000",
			3061 => "0011100010000000000100",
			3062 => "0000000011000000110101",
			3063 => "0000000011000000110101",
			3064 => "0000000011000000110101",
			3065 => "0001100111101000000100",
			3066 => "0000000011000000110101",
			3067 => "0001001101001000000100",
			3068 => "0000000011000000110101",
			3069 => "0000000011000000110101",
			3070 => "0000101100100100000100",
			3071 => "0000000011000000110101",
			3072 => "0001111101001000000100",
			3073 => "0000000011000000110101",
			3074 => "0001111100101100001100",
			3075 => "0000111001010100001000",
			3076 => "0000010110010000000100",
			3077 => "0000000011000000110101",
			3078 => "0000000011000000110101",
			3079 => "0000000011000000110101",
			3080 => "0000001111001100000100",
			3081 => "0000000011000000110101",
			3082 => "0000111111101000000100",
			3083 => "0000000011000000110101",
			3084 => "0000000011000000110101",
			3085 => "0000110011000000001000",
			3086 => "0011010011110000000100",
			3087 => "0000000011000011110001",
			3088 => "0000000011000011110001",
			3089 => "0001011100000000010100",
			3090 => "0001111000101000010000",
			3091 => "0011001010100100001000",
			3092 => "0001010011001000000100",
			3093 => "0000000011000011110001",
			3094 => "0000000011000011110001",
			3095 => "0000000101000100000100",
			3096 => "0000000011000011110001",
			3097 => "0000000011000011110001",
			3098 => "0000000011000011110001",
			3099 => "0011111101001100101100",
			3100 => "0000010110010000010100",
			3101 => "0000011000111100000100",
			3102 => "0000000011000011110001",
			3103 => "0011011010100100001000",
			3104 => "0011001110011000000100",
			3105 => "0000000011000011110001",
			3106 => "0000000011000011110001",
			3107 => "0011001100101000000100",
			3108 => "0000000011000011110001",
			3109 => "0000000011000011110001",
			3110 => "0011011011101100001000",
			3111 => "0000000100111100000100",
			3112 => "0000000011000011110001",
			3113 => "0000000011000011110001",
			3114 => "0001010110011100001000",
			3115 => "0010001001000100000100",
			3116 => "0000000011000011110001",
			3117 => "0000000011000011110001",
			3118 => "0001001100000000000100",
			3119 => "0000000011000011110001",
			3120 => "0000000011000011110001",
			3121 => "0001111100101100001100",
			3122 => "0010010101101100001000",
			3123 => "0011110000100100000100",
			3124 => "0000000011000011110001",
			3125 => "0000000011000011110001",
			3126 => "0000000011000011110001",
			3127 => "0010101011000000000100",
			3128 => "0000000011000011110001",
			3129 => "0001010011000100000100",
			3130 => "0000000011000011110001",
			3131 => "0000000011000011110001",
			3132 => "0011111100111101000100",
			3133 => "0000101111101100111000",
			3134 => "0010101000101000100000",
			3135 => "0000001011001000010100",
			3136 => "0001000111110000001000",
			3137 => "0001000001110000000100",
			3138 => "0000000011000111111101",
			3139 => "0000000011000111111101",
			3140 => "0011000011010000000100",
			3141 => "0000000011000111111101",
			3142 => "0011000111011100000100",
			3143 => "0000000011000111111101",
			3144 => "0000000011000111111101",
			3145 => "0011111011011100001000",
			3146 => "0011001010100100000100",
			3147 => "0000000011000111111101",
			3148 => "0000000011000111111101",
			3149 => "0000000011000111111101",
			3150 => "0000100110010100010100",
			3151 => "0001011010011100001000",
			3152 => "0001111001011000000100",
			3153 => "0000000011000111111101",
			3154 => "0000000011000111111101",
			3155 => "0001010010111000001000",
			3156 => "0000010111100100000100",
			3157 => "0000000011000111111101",
			3158 => "0000000011000111111101",
			3159 => "0000000011000111111101",
			3160 => "0000000011000111111101",
			3161 => "0011011100101000001000",
			3162 => "0000010111100100000100",
			3163 => "0000000011000111111101",
			3164 => "0000000011000111111101",
			3165 => "0000000011000111111101",
			3166 => "0011111000001000010000",
			3167 => "0010101100010000000100",
			3168 => "0000000011000111111101",
			3169 => "0001001000000100000100",
			3170 => "0000000011000111111101",
			3171 => "0001010000111100000100",
			3172 => "0000000011000111111101",
			3173 => "0000000011000111111101",
			3174 => "0001100000001100001100",
			3175 => "0011001010100100000100",
			3176 => "0000000011000111111101",
			3177 => "0010110011010000000100",
			3178 => "0000000011000111111101",
			3179 => "0000000011000111111101",
			3180 => "0010011001000100010100",
			3181 => "0011110111001100001100",
			3182 => "0000111001010100001000",
			3183 => "0001000111011100000100",
			3184 => "0000000011000111111101",
			3185 => "0000000011000111111101",
			3186 => "0000000011000111111101",
			3187 => "0011110111111100000100",
			3188 => "0000000011000111111101",
			3189 => "0000000011000111111101",
			3190 => "0001001111011000001000",
			3191 => "0011001001001000000100",
			3192 => "0000000011000111111101",
			3193 => "0000000011000111111101",
			3194 => "0010101011000000000100",
			3195 => "0000000011000111111101",
			3196 => "0010101001011000000100",
			3197 => "0000000011000111111101",
			3198 => "0000000011000111111101",
			3199 => "0001001100000000101100",
			3200 => "0001001000000100101000",
			3201 => "0010001111011000100100",
			3202 => "0001110110011100100000",
			3203 => "0001011000101000010000",
			3204 => "0011010101010100001000",
			3205 => "0001001010000100000100",
			3206 => "0000000011001010101001",
			3207 => "0000000011001010101001",
			3208 => "0010101001010100000100",
			3209 => "1111111011001010101001",
			3210 => "0000000011001010101001",
			3211 => "0001010100101100001000",
			3212 => "0011100111001000000100",
			3213 => "0000001011001010101001",
			3214 => "0000000011001010101001",
			3215 => "0001111001010000000100",
			3216 => "1111111011001010101001",
			3217 => "0000000011001010101001",
			3218 => "1111111011001010101001",
			3219 => "1111111011001010101001",
			3220 => "0000001011001010101001",
			3221 => "0001001000111000000100",
			3222 => "1111111011001010101001",
			3223 => "0010001001000100010000",
			3224 => "0001110100101100001100",
			3225 => "0011000101011100000100",
			3226 => "1111111011001010101001",
			3227 => "0001010010111000000100",
			3228 => "0000000011001010101001",
			3229 => "0000000011001010101001",
			3230 => "0000000011001010101001",
			3231 => "0011100100010000010100",
			3232 => "0011010011010000001000",
			3233 => "0010101001000000000100",
			3234 => "0000001011001010101001",
			3235 => "0000000011001010101001",
			3236 => "0000111100101100000100",
			3237 => "1111111011001010101001",
			3238 => "0001010011110100000100",
			3239 => "0000001011001010101001",
			3240 => "0000000011001010101001",
			3241 => "1111111011001010101001",
			3242 => "0001110110011101011100",
			3243 => "0010110111011100100100",
			3244 => "0010001111001000100000",
			3245 => "0010110110001100001000",
			3246 => "0011001101000000000100",
			3247 => "0000000011001101110101",
			3248 => "0000000011001101110101",
			3249 => "0011100110110000001100",
			3250 => "0001100000010000001000",
			3251 => "0001011101001000000100",
			3252 => "0000000011001101110101",
			3253 => "0000000011001101110101",
			3254 => "0000000011001101110101",
			3255 => "0000010110010000000100",
			3256 => "0000000011001101110101",
			3257 => "0001000011010000000100",
			3258 => "0000000011001101110101",
			3259 => "0000000011001101110101",
			3260 => "0000000011001101110101",
			3261 => "0000010110010000010000",
			3262 => "0001010110101100001100",
			3263 => "0011011011101100000100",
			3264 => "0000000011001101110101",
			3265 => "0000010000011000000100",
			3266 => "0000000011001101110101",
			3267 => "0000000011001101110101",
			3268 => "0000000011001101110101",
			3269 => "0001011101001000001100",
			3270 => "0010000101101100001000",
			3271 => "0000111001000100000100",
			3272 => "0000000011001101110101",
			3273 => "0000000011001101110101",
			3274 => "0000000011001101110101",
			3275 => "0010010011000000001100",
			3276 => "0000000110111100001000",
			3277 => "0010011101101000000100",
			3278 => "0000000011001101110101",
			3279 => "0000000011001101110101",
			3280 => "0000000011001101110101",
			3281 => "0010111001001000001000",
			3282 => "0011010101010100000100",
			3283 => "0000000011001101110101",
			3284 => "0000000011001101110101",
			3285 => "0011001001000100000100",
			3286 => "0000000011001101110101",
			3287 => "0000000011001101110101",
			3288 => "0011101101100100001000",
			3289 => "0011011001001000000100",
			3290 => "0000000011001101110101",
			3291 => "0000000011001101110101",
			3292 => "0000000011001101110101",
			3293 => "0001111011111001111000",
			3294 => "0010111010100101000000",
			3295 => "0010010101011100100000",
			3296 => "0010111110011000011000",
			3297 => "0001100001100000001100",
			3298 => "0001101110001100000100",
			3299 => "0000000011010010100001",
			3300 => "0000001001110100000100",
			3301 => "0000000011010010100001",
			3302 => "0000000011010010100001",
			3303 => "0001111001010100001000",
			3304 => "0000110011001000000100",
			3305 => "0000000011010010100001",
			3306 => "0000000011010010100001",
			3307 => "0000000011010010100001",
			3308 => "0011100111001000000100",
			3309 => "0000000011010010100001",
			3310 => "0000000011010010100001",
			3311 => "0000100000101000010100",
			3312 => "0001111001010000001100",
			3313 => "0011100000110100001000",
			3314 => "0001100101110100000100",
			3315 => "0000000011010010100001",
			3316 => "0000000011010010100001",
			3317 => "0000000011010010100001",
			3318 => "0001001100101000000100",
			3319 => "0000000011010010100001",
			3320 => "0000000011010010100001",
			3321 => "0000010111100100001000",
			3322 => "0000111100010000000100",
			3323 => "0000000011010010100001",
			3324 => "0000000011010010100001",
			3325 => "0000000011010010100001",
			3326 => "0010101111101000011100",
			3327 => "0000010001100100010100",
			3328 => "0010101000111000001100",
			3329 => "0011010110001100000100",
			3330 => "0000000011010010100001",
			3331 => "0001010011001000000100",
			3332 => "0000000011010010100001",
			3333 => "0000000011010010100001",
			3334 => "0010110101011100000100",
			3335 => "0000000011010010100001",
			3336 => "0000000011010010100001",
			3337 => "0001011101001000000100",
			3338 => "0000000011010010100001",
			3339 => "0000000011010010100001",
			3340 => "0010001001000100001100",
			3341 => "0001001001010000000100",
			3342 => "0000000011010010100001",
			3343 => "0001010010111000000100",
			3344 => "0000000011010010100001",
			3345 => "0000000011010010100001",
			3346 => "0011110111000000001100",
			3347 => "0000011000011000000100",
			3348 => "0000000011010010100001",
			3349 => "0000111100101100000100",
			3350 => "0000000011010010100001",
			3351 => "0000000011010010100001",
			3352 => "0000000011010010100001",
			3353 => "0010101011000000001000",
			3354 => "0001001000111000000100",
			3355 => "0000000011010010100001",
			3356 => "0000000011010010100001",
			3357 => "0000001111001100001100",
			3358 => "0001010001001000000100",
			3359 => "0000000011010010100001",
			3360 => "0011100100010000000100",
			3361 => "0000000011010010100001",
			3362 => "0000000011010010100001",
			3363 => "0000100101101000000100",
			3364 => "0000000011010010100001",
			3365 => "0000100101010000000100",
			3366 => "0000000011010010100001",
			3367 => "0000000011010010100001",
			3368 => "0010110110001100001000",
			3369 => "0011001101000000000100",
			3370 => "0000000011010101010101",
			3371 => "1111111011010101010101",
			3372 => "0001000011010000011000",
			3373 => "0000011001100100000100",
			3374 => "1111111011010101010101",
			3375 => "0011000111011100010000",
			3376 => "0011100110000100001100",
			3377 => "0001101110001100000100",
			3378 => "0000000011010101010101",
			3379 => "0000010111100100000100",
			3380 => "0000001011010101010101",
			3381 => "0000000011010101010101",
			3382 => "0000000011010101010101",
			3383 => "0000000011010101010101",
			3384 => "0010100000111100110100",
			3385 => "0001100010000100011100",
			3386 => "0011111101001100010000",
			3387 => "0001101010111100001000",
			3388 => "0000110011001000000100",
			3389 => "0000000011010101010101",
			3390 => "0000000011010101010101",
			3391 => "0001010110011100000100",
			3392 => "1111111011010101010101",
			3393 => "0000000011010101010101",
			3394 => "0011001010100100000100",
			3395 => "1111111011010101010101",
			3396 => "0000001001101000000100",
			3397 => "0000001011010101010101",
			3398 => "0000000011010101010101",
			3399 => "0011110011111100001100",
			3400 => "0011101010001000000100",
			3401 => "1111111011010101010101",
			3402 => "0000100101101000000100",
			3403 => "1111111011010101010101",
			3404 => "0000000011010101010101",
			3405 => "0000001000110000001000",
			3406 => "0001101001111000000100",
			3407 => "0000001011010101010101",
			3408 => "0000000011010101010101",
			3409 => "0000000011010101010101",
			3410 => "0001011001000000000100",
			3411 => "0000000011010101010101",
			3412 => "1111111011010101010101",
			3413 => "0011000101010101011100",
			3414 => "0011000111011101001100",
			3415 => "0010111010100100110000",
			3416 => "0010001001001100011000",
			3417 => "0000001001110100001000",
			3418 => "0010011100101000000100",
			3419 => "0000000011011001111001",
			3420 => "0000000011011001111001",
			3421 => "0010010101011100001000",
			3422 => "0011001110011000000100",
			3423 => "0000000011011001111001",
			3424 => "0000000011011001111001",
			3425 => "0001011101001000000100",
			3426 => "0000000011011001111001",
			3427 => "0000000011011001111001",
			3428 => "0010010101101100010000",
			3429 => "0011100010000000001000",
			3430 => "0011010110110100000100",
			3431 => "0000000011011001111001",
			3432 => "0000000011011001111001",
			3433 => "0000000010100000000100",
			3434 => "0000000011011001111001",
			3435 => "0000000011011001111001",
			3436 => "0001111001010100000100",
			3437 => "0000000011011001111001",
			3438 => "0000000011011001111001",
			3439 => "0010101000101000010000",
			3440 => "0011011010100100001100",
			3441 => "0000010001110000000100",
			3442 => "0000000011011001111001",
			3443 => "0000110011000000000100",
			3444 => "0000000011011001111001",
			3445 => "0000000011011001111001",
			3446 => "0000000011011001111001",
			3447 => "0000111000101000000100",
			3448 => "0000000011011001111001",
			3449 => "0010011001000100000100",
			3450 => "0000000011011001111001",
			3451 => "0000000011011001111001",
			3452 => "0000010000011000000100",
			3453 => "0000000011011001111001",
			3454 => "0001011001010100000100",
			3455 => "0000000011011001111001",
			3456 => "0000111000101000000100",
			3457 => "0000000011011001111001",
			3458 => "0000000011011001111001",
			3459 => "0010111100101000101100",
			3460 => "0010000101101100011000",
			3461 => "0000010000011000001100",
			3462 => "0011011011101100000100",
			3463 => "0000000011011001111001",
			3464 => "0001011001010100000100",
			3465 => "0000000011011001111001",
			3466 => "0000000011011001111001",
			3467 => "0001010000111000000100",
			3468 => "0000000011011001111001",
			3469 => "0001111101001000000100",
			3470 => "0000000011011001111001",
			3471 => "0000000011011001111001",
			3472 => "0001011101001000000100",
			3473 => "0000000011011001111001",
			3474 => "0000011110011000001100",
			3475 => "0000001011100100001000",
			3476 => "0001010011000100000100",
			3477 => "0000000011011001111001",
			3478 => "0000000011011001111001",
			3479 => "0000000011011001111001",
			3480 => "0000000011011001111001",
			3481 => "0000111011000000000100",
			3482 => "0000000011011001111001",
			3483 => "0010100000111100000100",
			3484 => "0000000011011001111001",
			3485 => "0000000011011001111001",
			3486 => "0001101010111101000000",
			3487 => "0000000101101000111100",
			3488 => "0000001010010100110100",
			3489 => "0010010101011100010100",
			3490 => "0010110110001100001000",
			3491 => "0011000110110100000100",
			3492 => "0000000011011101010101",
			3493 => "0000000011011101010101",
			3494 => "0010001010100100000100",
			3495 => "0000000011011101010101",
			3496 => "0010101000000100000100",
			3497 => "0000000011011101010101",
			3498 => "0000000011011101010101",
			3499 => "0000010110010000010000",
			3500 => "0010001001000100001000",
			3501 => "0010100011001000000100",
			3502 => "0000000011011101010101",
			3503 => "0000000011011101010101",
			3504 => "0001111001010000000100",
			3505 => "0000000011011101010101",
			3506 => "0000000011011101010101",
			3507 => "0000010001100100001000",
			3508 => "0011001010100100000100",
			3509 => "0000000011011101010101",
			3510 => "0000000011011101010101",
			3511 => "0000000110111100000100",
			3512 => "0000000011011101010101",
			3513 => "0000000011011101010101",
			3514 => "0010001111001000000100",
			3515 => "0000000011011101010101",
			3516 => "0000000011011101010101",
			3517 => "0000000011011101010101",
			3518 => "0011111101001100001000",
			3519 => "0010101000101000000100",
			3520 => "0000000011011101010101",
			3521 => "0000000011011101010101",
			3522 => "0001100000001100001000",
			3523 => "0011011011101100000100",
			3524 => "0000000011011101010101",
			3525 => "0000000011011101010101",
			3526 => "0000101111001100010000",
			3527 => "0011000101010100000100",
			3528 => "0000000011011101010101",
			3529 => "0000111000101000001000",
			3530 => "0011110000101100000100",
			3531 => "0000000011011101010101",
			3532 => "0000000011011101010101",
			3533 => "0000000011011101010101",
			3534 => "0001011000111000000100",
			3535 => "0000000011011101010101",
			3536 => "0011110100110100000100",
			3537 => "0000000011011101010101",
			3538 => "0011111110011100000100",
			3539 => "0000000011011101010101",
			3540 => "0000000011011101010101",
			3541 => "0011111101100100000100",
			3542 => "1111111011011111100001",
			3543 => "0001110011000101000000",
			3544 => "0011010110001100011000",
			3545 => "0001000101111000010100",
			3546 => "0000011001100100000100",
			3547 => "0000001011011111100001",
			3548 => "0010111011101100001000",
			3549 => "0001100100000100000100",
			3550 => "0000001011011111100001",
			3551 => "1111111011011111100001",
			3552 => "0000111111011000000100",
			3553 => "0000000011011111100001",
			3554 => "0000001011011111100001",
			3555 => "1111111011011111100001",
			3556 => "0011001010100100001000",
			3557 => "0001011000000000000100",
			3558 => "1111111011011111100001",
			3559 => "0000000011011111100001",
			3560 => "0000010111110000010000",
			3561 => "0001010110101100001000",
			3562 => "0000000010101100000100",
			3563 => "1111111011011111100001",
			3564 => "0000000011011111100001",
			3565 => "0010011001000100000100",
			3566 => "1111111011011111100001",
			3567 => "1111111011011111100001",
			3568 => "0000010001100100001000",
			3569 => "0000111111101000000100",
			3570 => "0000001011011111100001",
			3571 => "0000000011011111100001",
			3572 => "0001011101001000000100",
			3573 => "1111111011011111100001",
			3574 => "0000000011011111100001",
			3575 => "1111111011011111100001",
			3576 => "0011111101100100000100",
			3577 => "1111111011100001111111",
			3578 => "0001110011000101001000",
			3579 => "0011010110001100011000",
			3580 => "0001000101111000010100",
			3581 => "0011110101111100001000",
			3582 => "0000110011000000000100",
			3583 => "0000000011100001111111",
			3584 => "0000001011100001111111",
			3585 => "0011101101100100001000",
			3586 => "0001101010111100000100",
			3587 => "0000000011100001111111",
			3588 => "1111111011100001111111",
			3589 => "0000001011100001111111",
			3590 => "1111111011100001111111",
			3591 => "0000010111110000010000",
			3592 => "0001010110101100001000",
			3593 => "0001101110001000000100",
			3594 => "0000000011100001111111",
			3595 => "0000001011100001111111",
			3596 => "0010011001000100000100",
			3597 => "1111111011100001111111",
			3598 => "1111111011100001111111",
			3599 => "0001011101001000010000",
			3600 => "0010001001000100001000",
			3601 => "0001100000010000000100",
			3602 => "0000001011100001111111",
			3603 => "1111111011100001111111",
			3604 => "0001011100010000000100",
			3605 => "1111111011100001111111",
			3606 => "1111110011100001111111",
			3607 => "0000001011100100001000",
			3608 => "0000011000011000000100",
			3609 => "0000000011100001111111",
			3610 => "1111111011100001111111",
			3611 => "0011011100101000000100",
			3612 => "0000001011100001111111",
			3613 => "0000000011100001111111",
			3614 => "1111111011100001111111",
			3615 => "0011111101100100010000",
			3616 => "0010011010100100000100",
			3617 => "0000001011100011011001",
			3618 => "0011000111011100001000",
			3619 => "0010010110000000000100",
			3620 => "1111111011100011011001",
			3621 => "0000001011100011011001",
			3622 => "1111111011100011011001",
			3623 => "0010011111011000011100",
			3624 => "0011101001011100000100",
			3625 => "0000001011100011011001",
			3626 => "0000110011000000001000",
			3627 => "0000001101011100000100",
			3628 => "1111111011100011011001",
			3629 => "0000000011100011011001",
			3630 => "0011110100000100000100",
			3631 => "1111111011100011011001",
			3632 => "0011100100011100001000",
			3633 => "0001010011001000000100",
			3634 => "0000001011100011011001",
			3635 => "0000000011100011011001",
			3636 => "1111111011100011011001",
			3637 => "1111111011100011011001",
			3638 => "0000111101000000001000",
			3639 => "0001101001010100000100",
			3640 => "0000000011100101000101",
			3641 => "0000010011100101000101",
			3642 => "0001010001001000100000",
			3643 => "0010001010100100001000",
			3644 => "0001110011000000000100",
			3645 => "0000000011100101000101",
			3646 => "1111111011100101000101",
			3647 => "0000011000111100000100",
			3648 => "0000001011100101000101",
			3649 => "0010000011001000010000",
			3650 => "0001010110011100001000",
			3651 => "0010001010000100000100",
			3652 => "0000000011100101000101",
			3653 => "0000000011100101000101",
			3654 => "0010110111011100000100",
			3655 => "1111111011100101000101",
			3656 => "0000001011100101000101",
			3657 => "1111111011100101000101",
			3658 => "0010110111011100001000",
			3659 => "0011011110011000000100",
			3660 => "1111111011100101000101",
			3661 => "0000001011100101000101",
			3662 => "0001001000000000000100",
			3663 => "0000000011100101000101",
			3664 => "1111111011100101000101",
			3665 => "0010011010000100111000",
			3666 => "0000001011001000011000",
			3667 => "0001000111110000001000",
			3668 => "0001011111011100000100",
			3669 => "1111111011100111001001",
			3670 => "0000100011100111001001",
			3671 => "0000010111100100000100",
			3672 => "1111111011100111001001",
			3673 => "0011000011010000000100",
			3674 => "1111111011100111001001",
			3675 => "0011000111011100000100",
			3676 => "0000001011100111001001",
			3677 => "1111111011100111001001",
			3678 => "0011100110000100011100",
			3679 => "0000001010111000010100",
			3680 => "0001100000001100010000",
			3681 => "0001011000000000001000",
			3682 => "0010100011000000000100",
			3683 => "0000000011100111001001",
			3684 => "0000001011100111001001",
			3685 => "0000010110010000000100",
			3686 => "0000000011100111001001",
			3687 => "0000000011100111001001",
			3688 => "0000000011100111001001",
			3689 => "0010111010100100000100",
			3690 => "0000000011100111001001",
			3691 => "0000001011100111001001",
			3692 => "1111111011100111001001",
			3693 => "0001100101100000000100",
			3694 => "1111111011100111001001",
			3695 => "0000010110001100000100",
			3696 => "0000000011100111001001",
			3697 => "1111111011100111001001",
			3698 => "0000101000011100010000",
			3699 => "0011000111011100001100",
			3700 => "0011000011010000000100",
			3701 => "1111111011101000110101",
			3702 => "0000010111100100000100",
			3703 => "1111111011101000110101",
			3704 => "0000001011101000110101",
			3705 => "1111111011101000110101",
			3706 => "0010011111011000100100",
			3707 => "0010010111011100000100",
			3708 => "0000001011101000110101",
			3709 => "0000110011000000000100",
			3710 => "1111111011101000110101",
			3711 => "0001110110101100010000",
			3712 => "0001100100000100001000",
			3713 => "0010010101011100000100",
			3714 => "0000001011101000110101",
			3715 => "0000000011101000110101",
			3716 => "0011001110011000000100",
			3717 => "1111111011101000110101",
			3718 => "1111111011101000110101",
			3719 => "0000011000111100000100",
			3720 => "0000001011101000110101",
			3721 => "0000000110111100000100",
			3722 => "0000000011101000110101",
			3723 => "0000000011101000110101",
			3724 => "1111111011101000110101",
			3725 => "0011111101100100010000",
			3726 => "0010011010100100000100",
			3727 => "0000000011101010101001",
			3728 => "0011000111011100001000",
			3729 => "0010110111011100000100",
			3730 => "1111111011101010101001",
			3731 => "0000001011101010101001",
			3732 => "1111111011101010101001",
			3733 => "0010011111011000101000",
			3734 => "0011100100011100100100",
			3735 => "0000101011101000001000",
			3736 => "0011110100101000000100",
			3737 => "0000001011101010101001",
			3738 => "1111111011101010101001",
			3739 => "0011000101010100010000",
			3740 => "0010100100101100001000",
			3741 => "0000010001100100000100",
			3742 => "0000001011101010101001",
			3743 => "0000000011101010101001",
			3744 => "0000010111100100000100",
			3745 => "1111111011101010101001",
			3746 => "0000000011101010101001",
			3747 => "0010001111011000001000",
			3748 => "0000111101001000000100",
			3749 => "0000001011101010101001",
			3750 => "0000001011101010101001",
			3751 => "0000000011101010101001",
			3752 => "1111111011101010101001",
			3753 => "1111111011101010101001",
			3754 => "0001001100000001000100",
			3755 => "0001011001010000101100",
			3756 => "0000010001100100100000",
			3757 => "0001010110101100010100",
			3758 => "0001111011111000010000",
			3759 => "0010111010100100001000",
			3760 => "0001000110000000000100",
			3761 => "0000000011101101111101",
			3762 => "0000000011101101111101",
			3763 => "0010101000111000000100",
			3764 => "0000000011101101111101",
			3765 => "0000001011101101111101",
			3766 => "0000000011101101111101",
			3767 => "0011100111001000001000",
			3768 => "0000000000101000000100",
			3769 => "0000000011101101111101",
			3770 => "1111111011101101111101",
			3771 => "0000000011101101111101",
			3772 => "0000111000000000000100",
			3773 => "1111111011101101111101",
			3774 => "0011110000001000000100",
			3775 => "0000000011101101111101",
			3776 => "0000000011101101111101",
			3777 => "0010001111011000010100",
			3778 => "0010000101101100001000",
			3779 => "0011110101111100000100",
			3780 => "0000000011101101111101",
			3781 => "1111111011101101111101",
			3782 => "0000000010101100000100",
			3783 => "0000000011101101111101",
			3784 => "0001111011111000000100",
			3785 => "0000001011101101111101",
			3786 => "0000000011101101111101",
			3787 => "0000000011101101111101",
			3788 => "0011000101011100010100",
			3789 => "0001001001010000001000",
			3790 => "0010101011000000000100",
			3791 => "0000000011101101111101",
			3792 => "1111111011101101111101",
			3793 => "0001111100110000000100",
			3794 => "0000000011101101111101",
			3795 => "0000010000011000000100",
			3796 => "0000000011101101111101",
			3797 => "0000000011101101111101",
			3798 => "0010010011000000001000",
			3799 => "0001111101001000000100",
			3800 => "0000000011101101111101",
			3801 => "0000000011101101111101",
			3802 => "0011010011010000001000",
			3803 => "0011000101101100000100",
			3804 => "0000000011101101111101",
			3805 => "0000000011101101111101",
			3806 => "0000000011101101111101",
			3807 => "0000100101011000010100",
			3808 => "0010011010100100000100",
			3809 => "0000000011110000001001",
			3810 => "0011000111011100001100",
			3811 => "0010110111011100001000",
			3812 => "0000100100111100000100",
			3813 => "1111111011110000001001",
			3814 => "0000000011110000001001",
			3815 => "0000001011110000001001",
			3816 => "1111111011110000001001",
			3817 => "0010010101111000101100",
			3818 => "0011100010110100101000",
			3819 => "0011001010100100010100",
			3820 => "0001100101001100001100",
			3821 => "0000001011010000000100",
			3822 => "1111111011110000001001",
			3823 => "0010101101001000000100",
			3824 => "0000010011110000001001",
			3825 => "0000001011110000001001",
			3826 => "0011100100010000000100",
			3827 => "1111111011110000001001",
			3828 => "0000000011110000001001",
			3829 => "0001011000000100000100",
			3830 => "0000010011110000001001",
			3831 => "0010000101011100001000",
			3832 => "0011111000001000000100",
			3833 => "0000000011110000001001",
			3834 => "0000001011110000001001",
			3835 => "0000010001100100000100",
			3836 => "0000010011110000001001",
			3837 => "0000001011110000001001",
			3838 => "1111111011110000001001",
			3839 => "0011010101010100000100",
			3840 => "0000000011110000001001",
			3841 => "1111111011110000001001",
			3842 => "0000100101011000010100",
			3843 => "0001000111110000001000",
			3844 => "0001000001110000000100",
			3845 => "0000000011110010011101",
			3846 => "0000000011110010011101",
			3847 => "0001010110011100000100",
			3848 => "0000000011110010011101",
			3849 => "0000001110100000000100",
			3850 => "0000000011110010011101",
			3851 => "0000000011110010011101",
			3852 => "0000010110110100110000",
			3853 => "0000110011000000000100",
			3854 => "0000000011110010011101",
			3855 => "0001101101010000011100",
			3856 => "0010110101010100010000",
			3857 => "0010101000101000001000",
			3858 => "0001100100000100000100",
			3859 => "0000000011110010011101",
			3860 => "0000000011110010011101",
			3861 => "0000100110010100000100",
			3862 => "0000000011110010011101",
			3863 => "0000000011110010011101",
			3864 => "0011101101100000001000",
			3865 => "0010001010000100000100",
			3866 => "0000000011110010011101",
			3867 => "0000000011110010011101",
			3868 => "0000000011110010011101",
			3869 => "0000010110010000000100",
			3870 => "0000000011110010011101",
			3871 => "0000101111001100000100",
			3872 => "0000000011110010011101",
			3873 => "0011111011011000000100",
			3874 => "0000000011110010011101",
			3875 => "0000000011110010011101",
			3876 => "0000010011000000000100",
			3877 => "0000000011110010011101",
			3878 => "0000000011110010011101",
			3879 => "0010011010000101001100",
			3880 => "0011000101010100101000",
			3881 => "0011010101010100100100",
			3882 => "0001100000001100011000",
			3883 => "0010101011111000010000",
			3884 => "0011101110100000001000",
			3885 => "0010001111001000000100",
			3886 => "0000000011110101111001",
			3887 => "0000000011110101111001",
			3888 => "0011100100010000000100",
			3889 => "0000001011110101111001",
			3890 => "0000000011110101111001",
			3891 => "0010110011010000000100",
			3892 => "1111111011110101111001",
			3893 => "0000000011110101111001",
			3894 => "0000101110110000001000",
			3895 => "0000101011001100000100",
			3896 => "1111111011110101111001",
			3897 => "0000000011110101111001",
			3898 => "0000000011110101111001",
			3899 => "1111111011110101111001",
			3900 => "0010001001000100011000",
			3901 => "0001000110000000001000",
			3902 => "0001001100101000000100",
			3903 => "0000000011110101111001",
			3904 => "0000001011110101111001",
			3905 => "0001001001010000001000",
			3906 => "0001011011000000000100",
			3907 => "0000000011110101111001",
			3908 => "1111111011110101111001",
			3909 => "0001001011000000000100",
			3910 => "0000000011110101111001",
			3911 => "0000000011110101111001",
			3912 => "0001011001010100000100",
			3913 => "0000000011110101111001",
			3914 => "0001001000111000000100",
			3915 => "0000001011110101111001",
			3916 => "0000000011110101111001",
			3917 => "0000111111101000010000",
			3918 => "0001110100101100001100",
			3919 => "0001001001001000001000",
			3920 => "0001001100101000000100",
			3921 => "0000000011110101111001",
			3922 => "0000000011110101111001",
			3923 => "0000000011110101111001",
			3924 => "1111111011110101111001",
			3925 => "0001010011000100001000",
			3926 => "0001010110011100000100",
			3927 => "0000000011110101111001",
			3928 => "0000001011110101111001",
			3929 => "0010000011001000000100",
			3930 => "1111111011110101111001",
			3931 => "0000010110110100000100",
			3932 => "0000000011110101111001",
			3933 => "0000000011110101111001",
			3934 => "0010011010000100111100",
			3935 => "0011100110000100111000",
			3936 => "0011000101010100011100",
			3937 => "0011010101010100011000",
			3938 => "0001100000001100010000",
			3939 => "0010101000101000001000",
			3940 => "0001011001010000000100",
			3941 => "0000000011111000100101",
			3942 => "0000001011111000100101",
			3943 => "0000000110111100000100",
			3944 => "1111111011111000100101",
			3945 => "0000000011111000100101",
			3946 => "0000001001101000000100",
			3947 => "1111111011111000100101",
			3948 => "0000000011111000100101",
			3949 => "1111111011111000100101",
			3950 => "0011100011101100010100",
			3951 => "0000011000011000001100",
			3952 => "0010001001000100001000",
			3953 => "0001010000111000000100",
			3954 => "0000000011111000100101",
			3955 => "0000000011111000100101",
			3956 => "0000001011111000100101",
			3957 => "0011001100101000000100",
			3958 => "1111111011111000100101",
			3959 => "0000000011111000100101",
			3960 => "0000011001100000000100",
			3961 => "0000000011111000100101",
			3962 => "0000001011111000100101",
			3963 => "1111111011111000100101",
			3964 => "0000111111101000010000",
			3965 => "0001110100101100001100",
			3966 => "0001001001001000001000",
			3967 => "0001001100101000000100",
			3968 => "0000000011111000100101",
			3969 => "0000000011111000100101",
			3970 => "0000000011111000100101",
			3971 => "1111111011111000100101",
			3972 => "0011011100101000001000",
			3973 => "0000000000000000000100",
			3974 => "0000000011111000100101",
			3975 => "0000000011111000100101",
			3976 => "1111111011111000100101",
			3977 => "0000111101000000001000",
			3978 => "0011100110101100000100",
			3979 => "0000000011111010111001",
			3980 => "0000010011111010111001",
			3981 => "0000100101011000010100",
			3982 => "0000010111100100000100",
			3983 => "1111111011111010111001",
			3984 => "0011000111011100001100",
			3985 => "0000111101001000001000",
			3986 => "0010001111111100000100",
			3987 => "0000000011111010111001",
			3988 => "1111111011111010111001",
			3989 => "0000001011111010111001",
			3990 => "1111111011111010111001",
			3991 => "0011100000110100001000",
			3992 => "0010101011000000000100",
			3993 => "0000001011111010111001",
			3994 => "1111111011111010111001",
			3995 => "0001110110101100001100",
			3996 => "0010010101011100001000",
			3997 => "0001100100000100000100",
			3998 => "0000000011111010111001",
			3999 => "0000000011111010111001",
			4000 => "1111111011111010111001",
			4001 => "0011101111010100010000",
			4002 => "0000000110111100001000",
			4003 => "0000100011111000000100",
			4004 => "0000000011111010111001",
			4005 => "0000000011111010111001",
			4006 => "0011000101010100000100",
			4007 => "0000000011111010111001",
			4008 => "0000001011111010111001",
			4009 => "0000010001110000000100",
			4010 => "0000000011111010111001",
			4011 => "0010000101101100000100",
			4012 => "1111111011111010111001",
			4013 => "0000000011111010111001",
			4014 => "0000000011111000100100",
			4015 => "0010010101101100011000",
			4016 => "0010001001001100000100",
			4017 => "0000000011111110010101",
			4018 => "0010001111111100001100",
			4019 => "0001101110001100000100",
			4020 => "0000000011111110010101",
			4021 => "0011100010010100000100",
			4022 => "0000000011111110010101",
			4023 => "0000000011111110010101",
			4024 => "0001100111100000000100",
			4025 => "0000000011111110010101",
			4026 => "0000000011111110010101",
			4027 => "0011010110001100001000",
			4028 => "0001000110000000000100",
			4029 => "0000000011111110010101",
			4030 => "0000000011111110010101",
			4031 => "1111111011111110010101",
			4032 => "0001101010111100101000",
			4033 => "0000110011001000001000",
			4034 => "0011010110001100000100",
			4035 => "0000000011111110010101",
			4036 => "0000000011111110010101",
			4037 => "0001100101100000010100",
			4038 => "0010101111101000001000",
			4039 => "0001000110000000000100",
			4040 => "0000000011111110010101",
			4041 => "0000000011111110010101",
			4042 => "0000000110111100001000",
			4043 => "0001011010011100000100",
			4044 => "1111111011111110010101",
			4045 => "0000000011111110010101",
			4046 => "0000000011111110010101",
			4047 => "0000100000000000001000",
			4048 => "0001010001001000000100",
			4049 => "0000001011111110010101",
			4050 => "0000000011111110010101",
			4051 => "0000000011111110010101",
			4052 => "0011111101001100000100",
			4053 => "0000000011111110010101",
			4054 => "0000111000000000001100",
			4055 => "0000011000011000001000",
			4056 => "0000110011001000000100",
			4057 => "0000000011111110010101",
			4058 => "0000000011111110010101",
			4059 => "1111111011111110010101",
			4060 => "0011100011101000001000",
			4061 => "0010010101101100000100",
			4062 => "0000000011111110010101",
			4063 => "0000000011111110010101",
			4064 => "0000111100010000000100",
			4065 => "0000000011111110010101",
			4066 => "0010010101111000000100",
			4067 => "1111111011111110010101",
			4068 => "0000000011111110010101",
			4069 => "0000001011001000100000",
			4070 => "0001000111110000001100",
			4071 => "0001000001110000000100",
			4072 => "0000000100000001101001",
			4073 => "0001100011001000000100",
			4074 => "0000000100000001101001",
			4075 => "0000000100000001101001",
			4076 => "0001010110011100001100",
			4077 => "0011010111011100000100",
			4078 => "0000000100000001101001",
			4079 => "0011010101010100000100",
			4080 => "0000000100000001101001",
			4081 => "0000000100000001101001",
			4082 => "0001011000100000000100",
			4083 => "0000000100000001101001",
			4084 => "0000000100000001101001",
			4085 => "0001101010101100101100",
			4086 => "0001110110101100010000",
			4087 => "0001101010001000000100",
			4088 => "0000000100000001101001",
			4089 => "0011001110011000001000",
			4090 => "0010001001001100000100",
			4091 => "0000000100000001101001",
			4092 => "0000000100000001101001",
			4093 => "0000000100000001101001",
			4094 => "0001011100110000000100",
			4095 => "0000000100000001101001",
			4096 => "0000101011010000001100",
			4097 => "0011000101011100000100",
			4098 => "0000000100000001101001",
			4099 => "0000000010101100000100",
			4100 => "0000000100000001101001",
			4101 => "0000000100000001101001",
			4102 => "0000000101101000001000",
			4103 => "0010010101111000000100",
			4104 => "0000000100000001101001",
			4105 => "0000000100000001101001",
			4106 => "0000000100000001101001",
			4107 => "0000101100100100000100",
			4108 => "0000000100000001101001",
			4109 => "0001111101001000000100",
			4110 => "0000000100000001101001",
			4111 => "0001111100101100001100",
			4112 => "0000111001010100001000",
			4113 => "0000010110010000000100",
			4114 => "0000000100000001101001",
			4115 => "0000000100000001101001",
			4116 => "0000000100000001101001",
			4117 => "0001011100101100000100",
			4118 => "0000000100000001101001",
			4119 => "0001010011000100000100",
			4120 => "0000000100000001101001",
			4121 => "0000000100000001101001",
			4122 => "0000111011000000110000",
			4123 => "0010011010100100001000",
			4124 => "0001000110001100000100",
			4125 => "0000011100000011001101",
			4126 => "0000001100000011001101",
			4127 => "0000110011000000000100",
			4128 => "1111111100000011001101",
			4129 => "0000011011101100100000",
			4130 => "0010110111011100010000",
			4131 => "0010010110000000001000",
			4132 => "0001011001010000000100",
			4133 => "0000000100000011001101",
			4134 => "0000000100000011001101",
			4135 => "0000011001100000000100",
			4136 => "0000000100000011001101",
			4137 => "1111111100000011001101",
			4138 => "0000010110010000001000",
			4139 => "0001010110101100000100",
			4140 => "0000001100000011001101",
			4141 => "1111111100000011001101",
			4142 => "0001010110011100000100",
			4143 => "0000000100000011001101",
			4144 => "0000001100000011001101",
			4145 => "1111111100000011001101",
			4146 => "1111111100000011001101",
			4147 => "0000101010000000011100",
			4148 => "0000100101011000010100",
			4149 => "0010011010100100000100",
			4150 => "0000000100000101101001",
			4151 => "0011000111011100001100",
			4152 => "0010000101101100000100",
			4153 => "1111111100000101101001",
			4154 => "0011000011010000000100",
			4155 => "1111111100000101101001",
			4156 => "0000001100000101101001",
			4157 => "1111111100000101101001",
			4158 => "0001110110101100000100",
			4159 => "0000001100000101101001",
			4160 => "1111111100000101101001",
			4161 => "0010011111011000110000",
			4162 => "0011100100011100101100",
			4163 => "0001011000000000001100",
			4164 => "0011010110110100000100",
			4165 => "0000100100000101101001",
			4166 => "0000110011000000000100",
			4167 => "1111111100000101101001",
			4168 => "0000010100000101101001",
			4169 => "0010010101101100010000",
			4170 => "0000000101101000001000",
			4171 => "0001001010000100000100",
			4172 => "0000010100000101101001",
			4173 => "1111111100000101101001",
			4174 => "0011001110011000000100",
			4175 => "0000000100000101101001",
			4176 => "1111111100000101101001",
			4177 => "0011010101010100001000",
			4178 => "0011111101001100000100",
			4179 => "0000010100000101101001",
			4180 => "0000100100000101101001",
			4181 => "0010010011000000000100",
			4182 => "0000010100000101101001",
			4183 => "0000000100000101101001",
			4184 => "1111111100000101101001",
			4185 => "1111111100000101101001",
			4186 => "0000001011001000010000",
			4187 => "0011010111011100000100",
			4188 => "0000000100001000110101",
			4189 => "0011010101010100001000",
			4190 => "0000011001100000000100",
			4191 => "0000000100001000110101",
			4192 => "0000000100001000110101",
			4193 => "0000000100001000110101",
			4194 => "0010000000110000111100",
			4195 => "0010111110011000011000",
			4196 => "0011100011010100000100",
			4197 => "0000000100001000110101",
			4198 => "0001111001010100001100",
			4199 => "0000011001100100000100",
			4200 => "0000000100001000110101",
			4201 => "0000010111100100000100",
			4202 => "0000000100001000110101",
			4203 => "0000000100001000110101",
			4204 => "0000010111100100000100",
			4205 => "0000000100001000110101",
			4206 => "0000000100001000110101",
			4207 => "0011111001111000010100",
			4208 => "0001000110000000001000",
			4209 => "0001100100000100000100",
			4210 => "0000000100001000110101",
			4211 => "0000000100001000110101",
			4212 => "0001110110011100001000",
			4213 => "0010101110111000000100",
			4214 => "0000000100001000110101",
			4215 => "0000000100001000110101",
			4216 => "0000000100001000110101",
			4217 => "0011100100011100001100",
			4218 => "0010011101101000001000",
			4219 => "0010101111101000000100",
			4220 => "0000000100001000110101",
			4221 => "0000000100001000110101",
			4222 => "0000000100001000110101",
			4223 => "0000000100001000110101",
			4224 => "0001000110101100010000",
			4225 => "0011110000000100000100",
			4226 => "0000000100001000110101",
			4227 => "0000001101011000000100",
			4228 => "0000000100001000110101",
			4229 => "0000001000001100000100",
			4230 => "0000000100001000110101",
			4231 => "0000000100001000110101",
			4232 => "0011110111010000000100",
			4233 => "0000000100001000110101",
			4234 => "0011110100011000000100",
			4235 => "0000000100001000110101",
			4236 => "0000000100001000110101",
			4237 => "0000111001010001011100",
			4238 => "0000001011010000101000",
			4239 => "0011001010100100010000",
			4240 => "0001011101000000000100",
			4241 => "0000000100001101000001",
			4242 => "0010101000111000000100",
			4243 => "0000000100001101000001",
			4244 => "0001001100101000000100",
			4245 => "0000000100001101000001",
			4246 => "0000000100001101000001",
			4247 => "0010101000101000010100",
			4248 => "0000000101000100001000",
			4249 => "0000110110101100000100",
			4250 => "0000000100001101000001",
			4251 => "0000000100001101000001",
			4252 => "0010001001000100001000",
			4253 => "0001110001010000000100",
			4254 => "0000000100001101000001",
			4255 => "0000000100001101000001",
			4256 => "0000000100001101000001",
			4257 => "0000000100001101000001",
			4258 => "0011010011010000100100",
			4259 => "0010111010100100011000",
			4260 => "0001100000001100001100",
			4261 => "0000101101110000001000",
			4262 => "0000100000101000000100",
			4263 => "0000000100001101000001",
			4264 => "0000000100001101000001",
			4265 => "0000000100001101000001",
			4266 => "0011100001000000000100",
			4267 => "0000000100001101000001",
			4268 => "0010010101011100000100",
			4269 => "0000000100001101000001",
			4270 => "0000000100001101000001",
			4271 => "0011011011101100000100",
			4272 => "0000000100001101000001",
			4273 => "0001001010000100000100",
			4274 => "0000000100001101000001",
			4275 => "0000000100001101000001",
			4276 => "0001011001010100000100",
			4277 => "0000000100001101000001",
			4278 => "0001001100000000001000",
			4279 => "0001110011000100000100",
			4280 => "0000000100001101000001",
			4281 => "0000000100001101000001",
			4282 => "0000000100001101000001",
			4283 => "0011001001001000011000",
			4284 => "0001001001010000010000",
			4285 => "0011111011010100001000",
			4286 => "0010001001001100000100",
			4287 => "0000000100001101000001",
			4288 => "0000000100001101000001",
			4289 => "0011110100110100000100",
			4290 => "0000000100001101000001",
			4291 => "0000000100001101000001",
			4292 => "0001000100101100000100",
			4293 => "0000000100001101000001",
			4294 => "0000000100001101000001",
			4295 => "0011011100101000001100",
			4296 => "0010111001001000001000",
			4297 => "0000001011111100000100",
			4298 => "0000000100001101000001",
			4299 => "0000000100001101000001",
			4300 => "0000000100001101000001",
			4301 => "0000010001100100000100",
			4302 => "0000000100001101000001",
			4303 => "0000000100001101000001",
			4304 => "0000111101000000001000",
			4305 => "0001101001010100000100",
			4306 => "0000000100001111011101",
			4307 => "0000011100001111011101",
			4308 => "0001010001001000111000",
			4309 => "0010001010100100001000",
			4310 => "0001110011000000000100",
			4311 => "0000000100001111011101",
			4312 => "1111111100001111011101",
			4313 => "0010001001001100010000",
			4314 => "0000001001110100000100",
			4315 => "1111111100001111011101",
			4316 => "0001011101001000001000",
			4317 => "0010101101001000000100",
			4318 => "0000001100001111011101",
			4319 => "0000000100001111011101",
			4320 => "0000000100001111011101",
			4321 => "0011000011010000010000",
			4322 => "0010101100010000001000",
			4323 => "0001000110000000000100",
			4324 => "0000000100001111011101",
			4325 => "0000001100001111011101",
			4326 => "0001001100101000000100",
			4327 => "0000000100001111011101",
			4328 => "1111111100001111011101",
			4329 => "0001010110011100001000",
			4330 => "0010001010000100000100",
			4331 => "0000000100001111011101",
			4332 => "0000000100001111011101",
			4333 => "0010110111011100000100",
			4334 => "1111111100001111011101",
			4335 => "0000001100001111011101",
			4336 => "0010110111011100001000",
			4337 => "0011011110011000000100",
			4338 => "1111111100001111011101",
			4339 => "0000001100001111011101",
			4340 => "0001001000000000000100",
			4341 => "0000000100001111011101",
			4342 => "1111111100001111011101",
			4343 => "0010011010100100000100",
			4344 => "0000001100010001010001",
			4345 => "0000110011000000000100",
			4346 => "1111111100010001010001",
			4347 => "0001010011001000010100",
			4348 => "0010101000111000001000",
			4349 => "0010010101101100000100",
			4350 => "0000001100010001010001",
			4351 => "0000000100010001010001",
			4352 => "0010011001001000000100",
			4353 => "1111111100010001010001",
			4354 => "0010001111001000000100",
			4355 => "0000001100010001010001",
			4356 => "0000000100010001010001",
			4357 => "0010101110111000011100",
			4358 => "0001101010101100001100",
			4359 => "0000111111011000000100",
			4360 => "1111111100010001010001",
			4361 => "0011111000001000000100",
			4362 => "0000000100010001010001",
			4363 => "0000001100010001010001",
			4364 => "0011111101001100001000",
			4365 => "0001010110011100000100",
			4366 => "1111111100010001010001",
			4367 => "0000000100010001010001",
			4368 => "0000010001110000000100",
			4369 => "0000001100010001010001",
			4370 => "0000000100010001010001",
			4371 => "1111111100010001010001",
			4372 => "0000000011111000100100",
			4373 => "0001111100010000011100",
			4374 => "0010111010100100010000",
			4375 => "0001000111110000000100",
			4376 => "0000000100010101001101",
			4377 => "0000011001100100001000",
			4378 => "0001010011001000000100",
			4379 => "0000000100010101001101",
			4380 => "0000000100010101001101",
			4381 => "0000000100010101001101",
			4382 => "0001111100000000000100",
			4383 => "0000000100010101001101",
			4384 => "0011000111011100000100",
			4385 => "0000000100010101001101",
			4386 => "0000000100010101001101",
			4387 => "0010011100101000000100",
			4388 => "0000000100010101001101",
			4389 => "0000000100010101001101",
			4390 => "0011111100111100100100",
			4391 => "0010010101011100001000",
			4392 => "0001111100010000000100",
			4393 => "0000000100010101001101",
			4394 => "0000000100010101001101",
			4395 => "0000010111100100001000",
			4396 => "0011111110101100000100",
			4397 => "0000000100010101001101",
			4398 => "0000000100010101001101",
			4399 => "0011110111000000001100",
			4400 => "0000000010100100000100",
			4401 => "0000000100010101001101",
			4402 => "0010110101010100000100",
			4403 => "0000000100010101001101",
			4404 => "0000000100010101001101",
			4405 => "0010010011000000000100",
			4406 => "0000000100010101001101",
			4407 => "0000000100010101001101",
			4408 => "0011111101001100010100",
			4409 => "0001001111011000001100",
			4410 => "0011010110110100000100",
			4411 => "0000000100010101001101",
			4412 => "0010110111011100000100",
			4413 => "0000000100010101001101",
			4414 => "0000000100010101001101",
			4415 => "0000111111101000000100",
			4416 => "0000000100010101001101",
			4417 => "0000000100010101001101",
			4418 => "0011100011101000010100",
			4419 => "0001011100110000001000",
			4420 => "0000010111100100000100",
			4421 => "0000000100010101001101",
			4422 => "0000000100010101001101",
			4423 => "0001101101010000001000",
			4424 => "0011011011101100000100",
			4425 => "0000000100010101001101",
			4426 => "0000000100010101001101",
			4427 => "0000000100010101001101",
			4428 => "0001110001010000000100",
			4429 => "0000000100010101001101",
			4430 => "0010010101111000000100",
			4431 => "0000000100010101001101",
			4432 => "0001101110101100000100",
			4433 => "0000000100010101001101",
			4434 => "0000000100010101001101",
			4435 => "0000000011111000011100",
			4436 => "0001110110101100011000",
			4437 => "0010001001001100000100",
			4438 => "0000000100011000010001",
			4439 => "0011111101100100010000",
			4440 => "0001000111110000000100",
			4441 => "0000000100011000010001",
			4442 => "0001010110011100000100",
			4443 => "0000000100011000010001",
			4444 => "0001010000111100000100",
			4445 => "0000000100011000010001",
			4446 => "0000000100011000010001",
			4447 => "0000000100011000010001",
			4448 => "0000000100011000010001",
			4449 => "0011010011010000110000",
			4450 => "0001110110101100010000",
			4451 => "0011100010001000000100",
			4452 => "0000000100011000010001",
			4453 => "0001000101010100000100",
			4454 => "0000000100011000010001",
			4455 => "0001100100000100000100",
			4456 => "0000000100011000010001",
			4457 => "0000000100011000010001",
			4458 => "0010100100101100010100",
			4459 => "0011101000101100010000",
			4460 => "0001001001000100001000",
			4461 => "0010111110011000000100",
			4462 => "0000000100011000010001",
			4463 => "0000000100011000010001",
			4464 => "0001000110000000000100",
			4465 => "0000000100011000010001",
			4466 => "0000000100011000010001",
			4467 => "0000000100011000010001",
			4468 => "0001001000000000001000",
			4469 => "0011101100011000000100",
			4470 => "0000000100011000010001",
			4471 => "0000000100011000010001",
			4472 => "0000000100011000010001",
			4473 => "0000000010100100000100",
			4474 => "0000000100011000010001",
			4475 => "0001011101001000000100",
			4476 => "0000000100011000010001",
			4477 => "0001010011000100001100",
			4478 => "0000101000010000000100",
			4479 => "0000000100011000010001",
			4480 => "0001001111011000000100",
			4481 => "0000000100011000010001",
			4482 => "0000000100011000010001",
			4483 => "0000000100011000010001",
			4484 => "0010000000110001011100",
			4485 => "0011000011010000110000",
			4486 => "0001001010000100101000",
			4487 => "0011110101000100011100",
			4488 => "0000001011010000010000",
			4489 => "0011001010100100001000",
			4490 => "0001010110001100000100",
			4491 => "0000000100011011110101",
			4492 => "0000000100011011110101",
			4493 => "0001010011001000000100",
			4494 => "0000000100011011110101",
			4495 => "0000000100011011110101",
			4496 => "0010101101001000000100",
			4497 => "0000000100011011110101",
			4498 => "0011100011101100000100",
			4499 => "0000000100011011110101",
			4500 => "0000000100011011110101",
			4501 => "0001000101011100001000",
			4502 => "0001001010100100000100",
			4503 => "0000000100011011110101",
			4504 => "0000000100011011110101",
			4505 => "0000000100011011110101",
			4506 => "0010111010100100000100",
			4507 => "0000000100011011110101",
			4508 => "0000000100011011110101",
			4509 => "0000101100100100100000",
			4510 => "0001101100000100011000",
			4511 => "0011000111011100001100",
			4512 => "0010101000101000001000",
			4513 => "0001111100000000000100",
			4514 => "0000000100011011110101",
			4515 => "0000000100011011110101",
			4516 => "0000000100011011110101",
			4517 => "0010001001000100000100",
			4518 => "0000000100011011110101",
			4519 => "0011010011010000000100",
			4520 => "0000000100011011110101",
			4521 => "0000000100011011110101",
			4522 => "0001001100101000000100",
			4523 => "0000000100011011110101",
			4524 => "0000000100011011110101",
			4525 => "0011100011101000001000",
			4526 => "0001011011000000000100",
			4527 => "0000000100011011110101",
			4528 => "0000000100011011110101",
			4529 => "0000000100011011110101",
			4530 => "0001101010111100001100",
			4531 => "0000001011100100001000",
			4532 => "0011100110110000000100",
			4533 => "0000000100011011110101",
			4534 => "0000000100011011110101",
			4535 => "0000000100011011110101",
			4536 => "0001001000111000000100",
			4537 => "0000000100011011110101",
			4538 => "0001001100010000000100",
			4539 => "0000000100011011110101",
			4540 => "0000000100011011110101",
			4541 => "0000101011010001000000",
			4542 => "0011111110101100110000",
			4543 => "0000001001110100100100",
			4544 => "0001011000000100010000",
			4545 => "0011001010100100001000",
			4546 => "0000111101000000000100",
			4547 => "0000000100100000001001",
			4548 => "0000000100100000001001",
			4549 => "0000100110011000000100",
			4550 => "0000000100100000001001",
			4551 => "0000000100100000001001",
			4552 => "0001010001010000001000",
			4553 => "0001000101111000000100",
			4554 => "1111111100100000001001",
			4555 => "0000000100100000001001",
			4556 => "0010101011000000001000",
			4557 => "0011011010100100000100",
			4558 => "0000000100100000001001",
			4559 => "0000000100100000001001",
			4560 => "0000000100100000001001",
			4561 => "0011100011010100000100",
			4562 => "0000000100100000001001",
			4563 => "0001101110010000000100",
			4564 => "0000000100100000001001",
			4565 => "0000000100100000001001",
			4566 => "0010110101010100001000",
			4567 => "0010000101011100000100",
			4568 => "0000000100100000001001",
			4569 => "1111111100100000001001",
			4570 => "0001100001111000000100",
			4571 => "0000000100100000001001",
			4572 => "0000000100100000001001",
			4573 => "0000000101101000101000",
			4574 => "0000100000101000100000",
			4575 => "0010111010100100010000",
			4576 => "0010010101011100001000",
			4577 => "0000101101011100000100",
			4578 => "0000000100100000001001",
			4579 => "0000000100100000001001",
			4580 => "0000010110010000000100",
			4581 => "1111111100100000001001",
			4582 => "0000000100100000001001",
			4583 => "0011100001000000001100",
			4584 => "0011110111010000000100",
			4585 => "0000000100100000001001",
			4586 => "0010001111011000000100",
			4587 => "0000000100100000001001",
			4588 => "0000000100100000001001",
			4589 => "0000000100100000001001",
			4590 => "0000111001010000000100",
			4591 => "0000000100100000001001",
			4592 => "0000000100100000001001",
			4593 => "0011111011000100001000",
			4594 => "0011000011010000000100",
			4595 => "0000000100100000001001",
			4596 => "0000000100100000001001",
			4597 => "0001111100101100001100",
			4598 => "0010010101101100001000",
			4599 => "0001011000111000000100",
			4600 => "0000000100100000001001",
			4601 => "1111111100100000001001",
			4602 => "0000000100100000001001",
			4603 => "0000111111101000000100",
			4604 => "0000000100100000001001",
			4605 => "0000111100101100001000",
			4606 => "0000100101101000000100",
			4607 => "0000000100100000001001",
			4608 => "0000000100100000001001",
			4609 => "0000000100100000001001",
			4610 => "0000101011010000111100",
			4611 => "0011111110101100110000",
			4612 => "0000001001110100100100",
			4613 => "0001011000000100010000",
			4614 => "0011001010100100001000",
			4615 => "0000111101000000000100",
			4616 => "0000000100100100001101",
			4617 => "0000000100100100001101",
			4618 => "0000100110011000000100",
			4619 => "0000000100100100001101",
			4620 => "0000000100100100001101",
			4621 => "0001010001010000001000",
			4622 => "0001000101111000000100",
			4623 => "1111111100100100001101",
			4624 => "0000000100100100001101",
			4625 => "0010101011000000001000",
			4626 => "0011011010100100000100",
			4627 => "0000000100100100001101",
			4628 => "0000000100100100001101",
			4629 => "0000000100100100001101",
			4630 => "0011100011010100000100",
			4631 => "0000000100100100001101",
			4632 => "0001101110010000000100",
			4633 => "0000000100100100001101",
			4634 => "0000000100100100001101",
			4635 => "0010110101010100000100",
			4636 => "1111111100100100001101",
			4637 => "0001100001111000000100",
			4638 => "0000000100100100001101",
			4639 => "0000000100100100001101",
			4640 => "0000000101101000100100",
			4641 => "0001110110101100001000",
			4642 => "0001010110101100000100",
			4643 => "0000000100100100001101",
			4644 => "0000000100100100001101",
			4645 => "0011100001000000011000",
			4646 => "0010111010100100001000",
			4647 => "0010011100101000000100",
			4648 => "0000000100100100001101",
			4649 => "0000000100100100001101",
			4650 => "0000111011111000001000",
			4651 => "0010001111011000000100",
			4652 => "0000001100100100001101",
			4653 => "0000000100100100001101",
			4654 => "0011110101111100000100",
			4655 => "0000000100100100001101",
			4656 => "0000000100100100001101",
			4657 => "0000000100100100001101",
			4658 => "0011111011000100001000",
			4659 => "0011000011010000000100",
			4660 => "0000000100100100001101",
			4661 => "0000000100100100001101",
			4662 => "0001111100101100001100",
			4663 => "0010010101101100001000",
			4664 => "0001011000111000000100",
			4665 => "0000000100100100001101",
			4666 => "1111111100100100001101",
			4667 => "0000000100100100001101",
			4668 => "0000111111101000000100",
			4669 => "0000000100100100001101",
			4670 => "0000111100101100001000",
			4671 => "0000100101101000000100",
			4672 => "0000000100100100001101",
			4673 => "0000000100100100001101",
			4674 => "0000000100100100001101",
			4675 => "0001101010111101001100",
			4676 => "0000100110101000111100",
			4677 => "0010101000101000100100",
			4678 => "0011101111110100011100",
			4679 => "0010101000111000001100",
			4680 => "0010011010100100000100",
			4681 => "0000000100100111110001",
			4682 => "0001011100110000000100",
			4683 => "0000000100100111110001",
			4684 => "0000000100100111110001",
			4685 => "0011011010100100001000",
			4686 => "0011000101010100000100",
			4687 => "0000000100100111110001",
			4688 => "0000000100100111110001",
			4689 => "0011010111011100000100",
			4690 => "0000000100100111110001",
			4691 => "0000000100100111110001",
			4692 => "0011101101100000000100",
			4693 => "0000000100100111110001",
			4694 => "0000000100100111110001",
			4695 => "0001011010011100001100",
			4696 => "0011100110110000001000",
			4697 => "0001001101101000000100",
			4698 => "0000000100100111110001",
			4699 => "0000000100100111110001",
			4700 => "0000000100100111110001",
			4701 => "0001010010111000001000",
			4702 => "0001111100010000000100",
			4703 => "0000000100100111110001",
			4704 => "0000000100100111110001",
			4705 => "0000000100100111110001",
			4706 => "0011100100001100000100",
			4707 => "0000000100100111110001",
			4708 => "0000000101101000001000",
			4709 => "0010100011000100000100",
			4710 => "0000000100100111110001",
			4711 => "0000000100100111110001",
			4712 => "0000000100100111110001",
			4713 => "0000010001110000000100",
			4714 => "0000000100100111110001",
			4715 => "0010010101101100001000",
			4716 => "0011110111001100000100",
			4717 => "0000000100100111110001",
			4718 => "0000000100100111110001",
			4719 => "0010011101101000001000",
			4720 => "0010101111101000000100",
			4721 => "0000000100100111110001",
			4722 => "0000000100100111110001",
			4723 => "0001001000000100001000",
			4724 => "0010111001001000000100",
			4725 => "0000000100100111110001",
			4726 => "0000000100100111110001",
			4727 => "0000001001101000000100",
			4728 => "0000000100100111110001",
			4729 => "0001001100010000000100",
			4730 => "0000000100100111110001",
			4731 => "0000000100100111110001",
			4732 => "0000000011111000000100",
			4733 => "0000000100101010100101",
			4734 => "0010101111101000101100",
			4735 => "0010101000111000001000",
			4736 => "0011010110001100000100",
			4737 => "0000000100101010100101",
			4738 => "0000000100101010100101",
			4739 => "0010001010000100011100",
			4740 => "0010111110011000010000",
			4741 => "0000110011100100001000",
			4742 => "0001101110101100000100",
			4743 => "0000000100101010100101",
			4744 => "0000000100101010100101",
			4745 => "0000101101011100000100",
			4746 => "0000000100101010100101",
			4747 => "0000000100101010100101",
			4748 => "0001000101111000001000",
			4749 => "0001100101100000000100",
			4750 => "0000000100101010100101",
			4751 => "0000000100101010100101",
			4752 => "0000000100101010100101",
			4753 => "0000000101010000000100",
			4754 => "0000000100101010100101",
			4755 => "0000000100101010100101",
			4756 => "0010110101010100011000",
			4757 => "0000111001010000001100",
			4758 => "0011000111011100001000",
			4759 => "0011110110011000000100",
			4760 => "0000000100101010100101",
			4761 => "0000000100101010100101",
			4762 => "0000000100101010100101",
			4763 => "0011101111110100000100",
			4764 => "0000000100101010100101",
			4765 => "0011111011000100000100",
			4766 => "0000000100101010100101",
			4767 => "0000000100101010100101",
			4768 => "0011011100101000001000",
			4769 => "0011100100101000000100",
			4770 => "0000000100101010100101",
			4771 => "0000000100101010100101",
			4772 => "0001001111011000001000",
			4773 => "0000000101101000000100",
			4774 => "0000000100101010100101",
			4775 => "0000000100101010100101",
			4776 => "0000000100101010100101",
			4777 => "0001001100000000111100",
			4778 => "0001001000000100111000",
			4779 => "0001001111011000110000",
			4780 => "0000001011001000011100",
			4781 => "0001000111110000001100",
			4782 => "0001000001110000000100",
			4783 => "0000000100101101110001",
			4784 => "0000010111110000000100",
			4785 => "0000000100101101110001",
			4786 => "0000000100101101110001",
			4787 => "0011010111011100001000",
			4788 => "0010010101101100000100",
			4789 => "0000000100101101110001",
			4790 => "0000000100101101110001",
			4791 => "0001001001001000000100",
			4792 => "0000000100101101110001",
			4793 => "0000000100101101110001",
			4794 => "0011100000110100000100",
			4795 => "0000000100101101110001",
			4796 => "0011100001101100001000",
			4797 => "0010010101011100000100",
			4798 => "0000000100101101110001",
			4799 => "1111111100101101110001",
			4800 => "0010111110011000000100",
			4801 => "0000000100101101110001",
			4802 => "0000000100101101110001",
			4803 => "0010011101101000000100",
			4804 => "0000000100101101110001",
			4805 => "0000000100101101110001",
			4806 => "0000000100101101110001",
			4807 => "0001000110101100010100",
			4808 => "0001011000100000001100",
			4809 => "0011110010101000000100",
			4810 => "0000000100101101110001",
			4811 => "0011110100110100000100",
			4812 => "0000000100101101110001",
			4813 => "0000000100101101110001",
			4814 => "0001010001001000000100",
			4815 => "0000000100101101110001",
			4816 => "0000000100101101110001",
			4817 => "0001000100101100010100",
			4818 => "0011000101010100000100",
			4819 => "0000000100101101110001",
			4820 => "0000101000011100000100",
			4821 => "0000000100101101110001",
			4822 => "0001001001010000001000",
			4823 => "0000000000000000000100",
			4824 => "0000000100101101110001",
			4825 => "0000000100101101110001",
			4826 => "0000000100101101110001",
			4827 => "0000000100101101110001",
			4828 => "0000000011111000100100",
			4829 => "0001000111110000001100",
			4830 => "0001000001110000000100",
			4831 => "0000000100110001100101",
			4832 => "0000010111110000000100",
			4833 => "0000000100110001100101",
			4834 => "0000000100110001100101",
			4835 => "0001010001010000001000",
			4836 => "0000111101001000000100",
			4837 => "0000000100110001100101",
			4838 => "0000000100110001100101",
			4839 => "0000010110010000000100",
			4840 => "0000000100110001100101",
			4841 => "0011000101011100001000",
			4842 => "0001111100000000000100",
			4843 => "0000000100110001100101",
			4844 => "0000000100110001100101",
			4845 => "0000000100110001100101",
			4846 => "0011111100111100100100",
			4847 => "0011001110011000000100",
			4848 => "0000000100110001100101",
			4849 => "0000010111100100001000",
			4850 => "0011111110101100000100",
			4851 => "0000000100110001100101",
			4852 => "0000000100110001100101",
			4853 => "0001001100000000001100",
			4854 => "0000010001100100000100",
			4855 => "0000000100110001100101",
			4856 => "0011110111010000000100",
			4857 => "0000000100110001100101",
			4858 => "0000000100110001100101",
			4859 => "0011000101101100000100",
			4860 => "0000000100110001100101",
			4861 => "0000000000000000000100",
			4862 => "0000000100110001100101",
			4863 => "0000000100110001100101",
			4864 => "0000100000101000011000",
			4865 => "0010101100010000000100",
			4866 => "0000000100110001100101",
			4867 => "0011000101010100001000",
			4868 => "0011111101001100000100",
			4869 => "1111111100110001100101",
			4870 => "0000000100110001100101",
			4871 => "0011110110011000000100",
			4872 => "0000000100110001100101",
			4873 => "0011111101001100000100",
			4874 => "0000000100110001100101",
			4875 => "0000000100110001100101",
			4876 => "0000000101101000000100",
			4877 => "0000000100110001100101",
			4878 => "0011101110100100001000",
			4879 => "0010001111111100000100",
			4880 => "0000000100110001100101",
			4881 => "0000000100110001100101",
			4882 => "0001111011111000001000",
			4883 => "0010010101101100000100",
			4884 => "0000000100110001100101",
			4885 => "0000000100110001100101",
			4886 => "0010101011000000000100",
			4887 => "0000000100110001100101",
			4888 => "0000000100110001100101",
			4889 => "0010010101011100011100",
			4890 => "0001101010111100010100",
			4891 => "0000001011010000001100",
			4892 => "0010101000000100001000",
			4893 => "0001000111110000000100",
			4894 => "0000000100110101100001",
			4895 => "0000000100110101100001",
			4896 => "0000000100110101100001",
			4897 => "0001001101101000000100",
			4898 => "0000000100110101100001",
			4899 => "0000000100110101100001",
			4900 => "0011001110011000000100",
			4901 => "0000000100110101100001",
			4902 => "0000000100110101100001",
			4903 => "0011000101010100111100",
			4904 => "0010101000101000101100",
			4905 => "0011000011010000011000",
			4906 => "0001111101001000001100",
			4907 => "0010000101101100000100",
			4908 => "0000000100110101100001",
			4909 => "0010001001000100000100",
			4910 => "0000000100110101100001",
			4911 => "0000000100110101100001",
			4912 => "0001111001010000000100",
			4913 => "0000000100110101100001",
			4914 => "0011100111100000000100",
			4915 => "0000000100110101100001",
			4916 => "0000000100110101100001",
			4917 => "0001111101001000001100",
			4918 => "0011000111011100001000",
			4919 => "0001111100000000000100",
			4920 => "0000000100110101100001",
			4921 => "0000000100110101100001",
			4922 => "0000000100110101100001",
			4923 => "0011101110100100000100",
			4924 => "0000000100110101100001",
			4925 => "0000000100110101100001",
			4926 => "0001001001001000000100",
			4927 => "0000000100110101100001",
			4928 => "0010110111011100001000",
			4929 => "0010011100101000000100",
			4930 => "0000000100110101100001",
			4931 => "0000000100110101100001",
			4932 => "0000000100110101100001",
			4933 => "0010000101101100010000",
			4934 => "0010110111011100001100",
			4935 => "0010001111111100001000",
			4936 => "0011011110011000000100",
			4937 => "0000000100110101100001",
			4938 => "0000000100110101100001",
			4939 => "0000000100110101100001",
			4940 => "0000000100110101100001",
			4941 => "0000011011101100010100",
			4942 => "0001011101001000000100",
			4943 => "0000000100110101100001",
			4944 => "0000001011100100001000",
			4945 => "0000010001100100000100",
			4946 => "0000000100110101100001",
			4947 => "0000000100110101100001",
			4948 => "0011100010110100000100",
			4949 => "0000000100110101100001",
			4950 => "0000000100110101100001",
			4951 => "0000000100110101100001",
			4952 => "0011111101100100001100",
			4953 => "0011000111011100001000",
			4954 => "0010110111011100000100",
			4955 => "1111111100111000000101",
			4956 => "0000001100111000000101",
			4957 => "1111111100111000000101",
			4958 => "0010001111011001000000",
			4959 => "0000111011000000111000",
			4960 => "0011000011010000100000",
			4961 => "0010010101011100010000",
			4962 => "0011111001111000001000",
			4963 => "0000001001110100000100",
			4964 => "0000000100111000000101",
			4965 => "0000001100111000000101",
			4966 => "0010111011101100000100",
			4967 => "1111111100111000000101",
			4968 => "0000000100111000000101",
			4969 => "0010101101001000001000",
			4970 => "0010101000000000000100",
			4971 => "1111111100111000000101",
			4972 => "0000000100111000000101",
			4973 => "0011101110100000000100",
			4974 => "1111111100111000000101",
			4975 => "0000000100111000000101",
			4976 => "0011100001000000010000",
			4977 => "0000100110111100001000",
			4978 => "0000010001100100000100",
			4979 => "0000001100111000000101",
			4980 => "0000000100111000000101",
			4981 => "0000100000000000000100",
			4982 => "0000010100111000000101",
			4983 => "0000001100111000000101",
			4984 => "0000001110101000000100",
			4985 => "1111111100111000000101",
			4986 => "0000001100111000000101",
			4987 => "0001110001010000000100",
			4988 => "0000000100111000000101",
			4989 => "1111111100111000000101",
			4990 => "0010010101111000000100",
			4991 => "0000000100111000000101",
			4992 => "1111111100111000000101",
			4993 => "0011111100111101011000",
			4994 => "0000000011111000110100",
			4995 => "0001000101101100011100",
			4996 => "0001001100101000010000",
			4997 => "0001000111110000001000",
			4998 => "0001000001110000000100",
			4999 => "0000000100111100101001",
			5000 => "0000000100111100101001",
			5001 => "0011111000010100000100",
			5002 => "0000000100111100101001",
			5003 => "0000000100111100101001",
			5004 => "0001111000000000000100",
			5005 => "0000000100111100101001",
			5006 => "0001111001010000000100",
			5007 => "0000000100111100101001",
			5008 => "0000000100111100101001",
			5009 => "0010011101101000001000",
			5010 => "0011100101110100000100",
			5011 => "0000000100111100101001",
			5012 => "0000000100111100101001",
			5013 => "0010110101010100001100",
			5014 => "0010110111011100000100",
			5015 => "0000000100111100101001",
			5016 => "0010011010000100000100",
			5017 => "0000000100111100101001",
			5018 => "0000000100111100101001",
			5019 => "0000000100111100101001",
			5020 => "0001001100000000010100",
			5021 => "0010101000111000000100",
			5022 => "0000000100111100101001",
			5023 => "0000010000011000000100",
			5024 => "0000000100111100101001",
			5025 => "0000010001100100000100",
			5026 => "0000000100111100101001",
			5027 => "0011011100101000000100",
			5028 => "0000000100111100101001",
			5029 => "0000000100111100101001",
			5030 => "0000111100101100001000",
			5031 => "0011100110110000000100",
			5032 => "0000000100111100101001",
			5033 => "0000000100111100101001",
			5034 => "0000110011000100000100",
			5035 => "0000000100111100101001",
			5036 => "0000000100111100101001",
			5037 => "0011111101001100010000",
			5038 => "0011010110001100001000",
			5039 => "0010101001010100000100",
			5040 => "0000000100111100101001",
			5041 => "0000000100111100101001",
			5042 => "0011011001001000000100",
			5043 => "0000000100111100101001",
			5044 => "0000000100111100101001",
			5045 => "0000010001110000000100",
			5046 => "0000000100111100101001",
			5047 => "0010010101101100001100",
			5048 => "0000000010100000001000",
			5049 => "0001000011010000000100",
			5050 => "0000000100111100101001",
			5051 => "0000000100111100101001",
			5052 => "0000000100111100101001",
			5053 => "0001101110101100001100",
			5054 => "0011010101010100000100",
			5055 => "0000000100111100101001",
			5056 => "0000100000101000000100",
			5057 => "0000000100111100101001",
			5058 => "0000000100111100101001",
			5059 => "0011110011111100001000",
			5060 => "0010101011000000000100",
			5061 => "0000000100111100101001",
			5062 => "0000000100111100101001",
			5063 => "0000101001101000000100",
			5064 => "0000000100111100101001",
			5065 => "0000000100111100101001",
			5066 => "0011111100111101000100",
			5067 => "0000101111101100111000",
			5068 => "0010101000101000100000",
			5069 => "0011000101010100011100",
			5070 => "0010110110001100001100",
			5071 => "0000011000011000001000",
			5072 => "0000011001100100000100",
			5073 => "0000000101000000110101",
			5074 => "0000000101000000110101",
			5075 => "0000000101000000110101",
			5076 => "0010101000111000001000",
			5077 => "0000000011111000000100",
			5078 => "0000000101000000110101",
			5079 => "0000000101000000110101",
			5080 => "0000001011001000000100",
			5081 => "0000000101000000110101",
			5082 => "0000000101000000110101",
			5083 => "0000000101000000110101",
			5084 => "0000100110010100010100",
			5085 => "0001001001010000001000",
			5086 => "0001111001011000000100",
			5087 => "0000000101000000110101",
			5088 => "0000000101000000110101",
			5089 => "0001010010111000001000",
			5090 => "0011100110100000000100",
			5091 => "0000000101000000110101",
			5092 => "0000000101000000110101",
			5093 => "0000000101000000110101",
			5094 => "0000000101000000110101",
			5095 => "0011011100101000001000",
			5096 => "0000010111100100000100",
			5097 => "0000000101000000110101",
			5098 => "0000000101000000110101",
			5099 => "0000000101000000110101",
			5100 => "0011111000001000010000",
			5101 => "0010101100010000000100",
			5102 => "0000000101000000110101",
			5103 => "0001001000000100000100",
			5104 => "0000000101000000110101",
			5105 => "0001010000111100000100",
			5106 => "0000000101000000110101",
			5107 => "0000000101000000110101",
			5108 => "0001100000001100001100",
			5109 => "0011001010100100000100",
			5110 => "0000000101000000110101",
			5111 => "0010110011010000000100",
			5112 => "0000000101000000110101",
			5113 => "0000000101000000110101",
			5114 => "0010011001000100010100",
			5115 => "0011110111001100001100",
			5116 => "0000111001010100001000",
			5117 => "0001000111011100000100",
			5118 => "0000000101000000110101",
			5119 => "0000000101000000110101",
			5120 => "0000000101000000110101",
			5121 => "0011110111111100000100",
			5122 => "0000000101000000110101",
			5123 => "0000000101000000110101",
			5124 => "0001001111011000001000",
			5125 => "0011001001001000000100",
			5126 => "0000000101000000110101",
			5127 => "0000000101000000110101",
			5128 => "0010101011000000000100",
			5129 => "0000000101000000110101",
			5130 => "0010101001011000000100",
			5131 => "0000000101000000110101",
			5132 => "0000000101000000110101",
			5133 => "0001101010111101011100",
			5134 => "0000010110010000101000",
			5135 => "0011001110011000010000",
			5136 => "0001001010000100001100",
			5137 => "0010001010100100000100",
			5138 => "0000000101000101010001",
			5139 => "0000001001110100000100",
			5140 => "0000000101000101010001",
			5141 => "0000000101000101010001",
			5142 => "0000000101000101010001",
			5143 => "0001000101101100010000",
			5144 => "0000110011001000001100",
			5145 => "0010010101011100000100",
			5146 => "0000000101000101010001",
			5147 => "0010011001001000000100",
			5148 => "0000000101000101010001",
			5149 => "0000000101000101010001",
			5150 => "0000000101000101010001",
			5151 => "0010001001000100000100",
			5152 => "0000000101000101010001",
			5153 => "0000000101000101010001",
			5154 => "0000000110111100101000",
			5155 => "0000010001100100011100",
			5156 => "0011000011010000001100",
			5157 => "0010001111111100000100",
			5158 => "0000000101000101010001",
			5159 => "0010011100101000000100",
			5160 => "0000000101000101010001",
			5161 => "0000000101000101010001",
			5162 => "0011111101100100001000",
			5163 => "0001010110011100000100",
			5164 => "0000000101000101010001",
			5165 => "0000000101000101010001",
			5166 => "0001110001010000000100",
			5167 => "0000000101000101010001",
			5168 => "0000000101000101010001",
			5169 => "0000010101101100001000",
			5170 => "0011100110110000000100",
			5171 => "0000000101000101010001",
			5172 => "0000000101000101010001",
			5173 => "0000000101000101010001",
			5174 => "0000001111001100001000",
			5175 => "0011010101010100000100",
			5176 => "0000000101000101010001",
			5177 => "0000000101000101010001",
			5178 => "0000000101000101010001",
			5179 => "0011111101001100001000",
			5180 => "0010101000101000000100",
			5181 => "0000000101000101010001",
			5182 => "0000000101000101010001",
			5183 => "0001100000001100001000",
			5184 => "0011011011101100000100",
			5185 => "0000000101000101010001",
			5186 => "0000000101000101010001",
			5187 => "0000101111001100010000",
			5188 => "0011000101010100000100",
			5189 => "0000000101000101010001",
			5190 => "0000111000101000001000",
			5191 => "0000111001010100000100",
			5192 => "0000000101000101010001",
			5193 => "0000000101000101010001",
			5194 => "0000000101000101010001",
			5195 => "0001000011000000001000",
			5196 => "0001101101010100000100",
			5197 => "0000000101000101010001",
			5198 => "0000000101000101010001",
			5199 => "0010101011000000000100",
			5200 => "0000000101000101010001",
			5201 => "0000001000001100000100",
			5202 => "0000000101000101010001",
			5203 => "0000000101000101010001",
			5204 => "0011100010110101001100",
			5205 => "0000001000001101001000",
			5206 => "0001101010111100110100",
			5207 => "0011101100011000100000",
			5208 => "0010010101011100010000",
			5209 => "0010111110011000001000",
			5210 => "0001100001100000000100",
			5211 => "0000000101001000000101",
			5212 => "0000000101001000000101",
			5213 => "0010001001001100000100",
			5214 => "0000001101001000000101",
			5215 => "0000000101001000000101",
			5216 => "0000110011001000001000",
			5217 => "0011010110110100000100",
			5218 => "0000000101001000000101",
			5219 => "1111111101001000000101",
			5220 => "0000010000011000000100",
			5221 => "1111111101001000000101",
			5222 => "0000000101001000000101",
			5223 => "0000100011001100001100",
			5224 => "0001111001011000000100",
			5225 => "1111111101001000000101",
			5226 => "0010101001011000000100",
			5227 => "0000000101001000000101",
			5228 => "0000000101001000000101",
			5229 => "0001010001001000000100",
			5230 => "0000001101001000000101",
			5231 => "0000000101001000000101",
			5232 => "0000101100100100000100",
			5233 => "1111111101001000000101",
			5234 => "0010011100101000000100",
			5235 => "1111111101001000000101",
			5236 => "0000000101101000000100",
			5237 => "0000000101001000000101",
			5238 => "0011100100010000000100",
			5239 => "0000000101001000000101",
			5240 => "0000000101001000000101",
			5241 => "0000000101001000000101",
			5242 => "0010010101111000000100",
			5243 => "1111111101001000000101",
			5244 => "0001101110101100001000",
			5245 => "0001100010010000000100",
			5246 => "0000000101001000000101",
			5247 => "0000000101001000000101",
			5248 => "0000000101001000000101",
			5249 => "0000011000111100010100",
			5250 => "0010101100010000001100",
			5251 => "0010010101011100001000",
			5252 => "0010101010000100000100",
			5253 => "0000000101001100000001",
			5254 => "0000000101001100000001",
			5255 => "0000000101001100000001",
			5256 => "0001000011000000000100",
			5257 => "0000000101001100000001",
			5258 => "0000000101001100000001",
			5259 => "0001101010101101000100",
			5260 => "0000010111100100100100",
			5261 => "0001011100010000010000",
			5262 => "0011100011101100001100",
			5263 => "0010101000111000001000",
			5264 => "0001000111110000000100",
			5265 => "0000000101001100000001",
			5266 => "0000000101001100000001",
			5267 => "0000000101001100000001",
			5268 => "0000000101001100000001",
			5269 => "0001101100000100001100",
			5270 => "0000000010101100001000",
			5271 => "0010001111111100000100",
			5272 => "0000000101001100000001",
			5273 => "0000000101001100000001",
			5274 => "0000000101001100000001",
			5275 => "0011111001111000000100",
			5276 => "1111111101001100000001",
			5277 => "0000000101001100000001",
			5278 => "0000001011100100011000",
			5279 => "0010101000101000010000",
			5280 => "0001000101010100001000",
			5281 => "0011000110001100000100",
			5282 => "0000000101001100000001",
			5283 => "0000000101001100000001",
			5284 => "0010001111001000000100",
			5285 => "0000000101001100000001",
			5286 => "0000000101001100000001",
			5287 => "0011100110110000000100",
			5288 => "0000000101001100000001",
			5289 => "0000000101001100000001",
			5290 => "0010110101011100000100",
			5291 => "0000000101001100000001",
			5292 => "0000000101001100000001",
			5293 => "0000010001110000000100",
			5294 => "0000000101001100000001",
			5295 => "0001011001010000010000",
			5296 => "0000001000110000001100",
			5297 => "0001000011010000001000",
			5298 => "0001001010100100000100",
			5299 => "0000000101001100000001",
			5300 => "0000000101001100000001",
			5301 => "1111111101001100000001",
			5302 => "0000000101001100000001",
			5303 => "0001010011000100010000",
			5304 => "0010000000110000001000",
			5305 => "0011110101000100000100",
			5306 => "0000000101001100000001",
			5307 => "0000000101001100000001",
			5308 => "0000111100010000000100",
			5309 => "0000000101001100000001",
			5310 => "0000000101001100000001",
			5311 => "0000000101001100000001",
			5312 => "0001110110011101101000",
			5313 => "0010110111011100110100",
			5314 => "0010001111001000110000",
			5315 => "0010010101101100011100",
			5316 => "0001100110000100001100",
			5317 => "0000001001110100001000",
			5318 => "0010001001001100000100",
			5319 => "0000000101001111100101",
			5320 => "0000000101001111100101",
			5321 => "0000000101001111100101",
			5322 => "0000100000101000001000",
			5323 => "0011010110110100000100",
			5324 => "0000000101001111100101",
			5325 => "0000000101001111100101",
			5326 => "0000001110110000000100",
			5327 => "0000000101001111100101",
			5328 => "0000000101001111100101",
			5329 => "0011100001101100001100",
			5330 => "0010100011001000000100",
			5331 => "0000000101001111100101",
			5332 => "0001010000111000000100",
			5333 => "0000000101001111100101",
			5334 => "0000000101001111100101",
			5335 => "0000111100110000000100",
			5336 => "0000000101001111100101",
			5337 => "0000000101001111100101",
			5338 => "0000000101001111100101",
			5339 => "0000010110010000010000",
			5340 => "0001010110101100001100",
			5341 => "0011011011101100000100",
			5342 => "0000000101001111100101",
			5343 => "0001111100010000000100",
			5344 => "0000000101001111100101",
			5345 => "0000000101001111100101",
			5346 => "0000000101001111100101",
			5347 => "0000000110111100011000",
			5348 => "0000011000011000001100",
			5349 => "0010001001000100000100",
			5350 => "0000000101001111100101",
			5351 => "0010111100101000000100",
			5352 => "0000000101001111100101",
			5353 => "0000000101001111100101",
			5354 => "0010110101010100000100",
			5355 => "0000000101001111100101",
			5356 => "0011011100101000000100",
			5357 => "0000000101001111100101",
			5358 => "0000000101001111100101",
			5359 => "0010010011000000001000",
			5360 => "0000011101000000000100",
			5361 => "0000001101001111100101",
			5362 => "0000000101001111100101",
			5363 => "0000000101001111100101",
			5364 => "0011101101100100001000",
			5365 => "0011011001001000000100",
			5366 => "0000000101001111100101",
			5367 => "0000000101001111100101",
			5368 => "0000000101001111100101",
			5369 => "0000011011101101101100",
			5370 => "0011000011010000101100",
			5371 => "0001001010000100011100",
			5372 => "0000011001100000011000",
			5373 => "0010110110001100001000",
			5374 => "0011010011110000000100",
			5375 => "0000000101010011000001",
			5376 => "1111111101010011000001",
			5377 => "0011110000001000001000",
			5378 => "0010000101011100000100",
			5379 => "0000000101010011000001",
			5380 => "0000000101010011000001",
			5381 => "0001111101001000000100",
			5382 => "1111111101010011000001",
			5383 => "0000000101010011000001",
			5384 => "1111111101010011000001",
			5385 => "0010111010100100001100",
			5386 => "0001111000111000001000",
			5387 => "0001110101111000000100",
			5388 => "0000000101010011000001",
			5389 => "0000000101010011000001",
			5390 => "1111111101010011000001",
			5391 => "0000000101010011000001",
			5392 => "0011111000001000101100",
			5393 => "0000010110010000010000",
			5394 => "0010001001000100000100",
			5395 => "1111111101010011000001",
			5396 => "0001011111101000001000",
			5397 => "0001111100010000000100",
			5398 => "0000000101010011000001",
			5399 => "0000001101010011000001",
			5400 => "0000000101010011000001",
			5401 => "0010000101101100001100",
			5402 => "0001111001010100001000",
			5403 => "0010101001000000000100",
			5404 => "0000001101010011000001",
			5405 => "0000000101010011000001",
			5406 => "1111111101010011000001",
			5407 => "0001000110000000001000",
			5408 => "0011101111110100000100",
			5409 => "0000000101010011000001",
			5410 => "1111111101010011000001",
			5411 => "0000001011100100000100",
			5412 => "0000000101010011000001",
			5413 => "0000000101010011000001",
			5414 => "0011100001000000001000",
			5415 => "0001001010000100000100",
			5416 => "0000000101010011000001",
			5417 => "0000001101010011000001",
			5418 => "0011110011111100001000",
			5419 => "0010101011000000000100",
			5420 => "1111111101010011000001",
			5421 => "0000000101010011000001",
			5422 => "0000000101010011000001",
			5423 => "1111111101010011000001",
			5424 => "0000011011101101110100",
			5425 => "0011000011010000110100",
			5426 => "0001001010000100100100",
			5427 => "0000011001100000100000",
			5428 => "0001100100110000010000",
			5429 => "0011010110001100001000",
			5430 => "0010110110001100000100",
			5431 => "0000000101010110101111",
			5432 => "0000001101010110101111",
			5433 => "0010010101011100000100",
			5434 => "0000000101010110101111",
			5435 => "0000000101010110101111",
			5436 => "0000010111110000001000",
			5437 => "0011111101001100000100",
			5438 => "1111111101010110101111",
			5439 => "0000000101010110101111",
			5440 => "0001011000000000000100",
			5441 => "0000000101010110101111",
			5442 => "0000001101010110101111",
			5443 => "1111111101010110101111",
			5444 => "0010111010100100001100",
			5445 => "0001111000111000001000",
			5446 => "0001110101111000000100",
			5447 => "0000000101010110101111",
			5448 => "0000000101010110101111",
			5449 => "1111111101010110101111",
			5450 => "0000000101010110101111",
			5451 => "0011111000001000101100",
			5452 => "0000010110010000001100",
			5453 => "0010001001000100000100",
			5454 => "1111111101010110101111",
			5455 => "0001111001010100000100",
			5456 => "0000000101010110101111",
			5457 => "0000001101010110101111",
			5458 => "0010000101101100010000",
			5459 => "0011000101010100001000",
			5460 => "0000000101000100000100",
			5461 => "0000000101010110101111",
			5462 => "0000001101010110101111",
			5463 => "0001010000111000000100",
			5464 => "1111111101010110101111",
			5465 => "0000000101010110101111",
			5466 => "0001000110000000001000",
			5467 => "0011101111110100000100",
			5468 => "0000000101010110101111",
			5469 => "1111111101010110101111",
			5470 => "0000011000011000000100",
			5471 => "0000001101010110101111",
			5472 => "0000000101010110101111",
			5473 => "0011100001000000001000",
			5474 => "0011011010100100000100",
			5475 => "0000000101010110101111",
			5476 => "0000001101010110101111",
			5477 => "0010101011000000001000",
			5478 => "0011111000100100000100",
			5479 => "1111111101010110101111",
			5480 => "0000000101010110101111",
			5481 => "0000000101010110101111",
			5482 => "1111111101010110101111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1943, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3615, initial_addr_3'length));
	end generate gen_rom_3;

	gen_rom_4: if SELECT_ROM = 4 generate
		bank <= (
			0 => "0000110011001000011000",
			1 => "0001100011101000001100",
			2 => "0001011000000000000100",
			3 => "0000000000000010010101",
			4 => "0001011100010000000100",
			5 => "0000000000000010010101",
			6 => "0000000000000010010101",
			7 => "0000001111001100001000",
			8 => "0011101100011000000100",
			9 => "0000000000000010010101",
			10 => "0000000000000010010101",
			11 => "0000000000000010010101",
			12 => "0010110111011100011100",
			13 => "0000010001100100010100",
			14 => "0000101100010100001100",
			15 => "0011110111100000000100",
			16 => "0000000000000010010101",
			17 => "0001011000000000000100",
			18 => "0000000000000010010101",
			19 => "0000000000000010010101",
			20 => "0000111011111000000100",
			21 => "0000000000000010010101",
			22 => "0000000000000010010101",
			23 => "0010010101101100000100",
			24 => "0000000000000010010101",
			25 => "0000000000000010010101",
			26 => "0000101011100100001000",
			27 => "0010010110000000000100",
			28 => "0000000000000010010101",
			29 => "0000000000000010010101",
			30 => "0010001010000100000100",
			31 => "0000000000000010010101",
			32 => "0011000110000000000100",
			33 => "0000000000000010010101",
			34 => "0000111111101000000100",
			35 => "0000000000000010010101",
			36 => "0000000000000010010101",
			37 => "0011011110011000100100",
			38 => "0000001011010000011000",
			39 => "0010001111111100001100",
			40 => "0011110111100000000100",
			41 => "0000000000000100111001",
			42 => "0001111001010100000100",
			43 => "0000000000000100111001",
			44 => "0000000000000100111001",
			45 => "0001110011001000000100",
			46 => "0000000000000100111001",
			47 => "0010100011000000000100",
			48 => "0000000000000100111001",
			49 => "0000000000000100111001",
			50 => "0011101110010000001000",
			51 => "0010101000000100000100",
			52 => "0000000000000100111001",
			53 => "0000000000000100111001",
			54 => "0000000000000100111001",
			55 => "0000101111101100011000",
			56 => "0010011001001000001000",
			57 => "0001001100101000000100",
			58 => "0000000000000100111001",
			59 => "0000000000000100111001",
			60 => "0000111100010000000100",
			61 => "0000000000000100111001",
			62 => "0001000011000000001000",
			63 => "0001001010000100000100",
			64 => "0000000000000100111001",
			65 => "0000000000000100111001",
			66 => "0000000000000100111001",
			67 => "0000011001100000000100",
			68 => "0000000000000100111001",
			69 => "0001001100000000001000",
			70 => "0001011101001000000100",
			71 => "0000000000000100111001",
			72 => "0000000000000100111001",
			73 => "0000001110101000000100",
			74 => "0000000000000100111001",
			75 => "0001111100011100000100",
			76 => "0000000000000100111001",
			77 => "0000000000000100111001",
			78 => "0001011100110000101100",
			79 => "0011001010100100010100",
			80 => "0000001001110100001000",
			81 => "0000000110001000000100",
			82 => "0000000000000111110101",
			83 => "0000000000000111110101",
			84 => "0001100101001100000100",
			85 => "0000000000000111110101",
			86 => "0011100110111000000100",
			87 => "0000000000000111110101",
			88 => "0000000000000111110101",
			89 => "0000110101111000001100",
			90 => "0010110111011100001000",
			91 => "0011111110101100000100",
			92 => "0000000000000111110101",
			93 => "0000000000000111110101",
			94 => "0000000000000111110101",
			95 => "0010110101011100000100",
			96 => "1111111000000111110101",
			97 => "0010010011000000000100",
			98 => "0000000000000111110101",
			99 => "0000000000000111110101",
			100 => "0010110011010000010100",
			101 => "0001011000101000010000",
			102 => "0010101001010100001000",
			103 => "0001111100110000000100",
			104 => "0000000000000111110101",
			105 => "0000000000000111110101",
			106 => "0000101010010100000100",
			107 => "0000000000000111110101",
			108 => "0000000000000111110101",
			109 => "0000000000000111110101",
			110 => "0000010111100100001000",
			111 => "0011110111000000000100",
			112 => "0000000000000111110101",
			113 => "0000001000000111110101",
			114 => "0001111000101000001100",
			115 => "0000011000011000000100",
			116 => "0000000000000111110101",
			117 => "0010011101101000000100",
			118 => "0000000000000111110101",
			119 => "0000000000000111110101",
			120 => "0001111001011000000100",
			121 => "1111111000000111110101",
			122 => "0011011100101000000100",
			123 => "0000000000000111110101",
			124 => "0000000000000111110101",
			125 => "0011101101100000110100",
			126 => "0001101100000100101000",
			127 => "0011000011010000010000",
			128 => "0011110111100000000100",
			129 => "0000000000001010101001",
			130 => "0000001011010000001000",
			131 => "0001010011001000000100",
			132 => "0000000000001010101001",
			133 => "0000000000001010101001",
			134 => "0000000000001010101001",
			135 => "0001110011001000001000",
			136 => "0011010110001100000100",
			137 => "0000000000001010101001",
			138 => "0000000000001010101001",
			139 => "0000011001100000000100",
			140 => "0000000000001010101001",
			141 => "0010101000101000000100",
			142 => "0000000000001010101001",
			143 => "0000011101000000000100",
			144 => "0000000000001010101001",
			145 => "0000000000001010101001",
			146 => "0001011001010100001000",
			147 => "0011111001111000000100",
			148 => "0000000000001010101001",
			149 => "0000000000001010101001",
			150 => "0000000000001010101001",
			151 => "0010011101101000010100",
			152 => "0011011011101100001100",
			153 => "0011110010101000000100",
			154 => "0000000000001010101001",
			155 => "0011110011111100000100",
			156 => "0000000000001010101001",
			157 => "0000000000001010101001",
			158 => "0001011111011000000100",
			159 => "0000000000001010101001",
			160 => "0000000000001010101001",
			161 => "0010001111001000000100",
			162 => "0000000000001010101001",
			163 => "0011001001000100001000",
			164 => "0000101000010000000100",
			165 => "0000000000001010101001",
			166 => "0000000000001010101001",
			167 => "0010011100000000000100",
			168 => "0000000000001010101001",
			169 => "0000000000001010101001",
			170 => "0011110001100000010100",
			171 => "0011010110001100001000",
			172 => "0011110100001100000100",
			173 => "1111111000001100101101",
			174 => "0000001000001100101101",
			175 => "0010010110000000001000",
			176 => "0010100100101100000100",
			177 => "1111111000001100101101",
			178 => "0000000000001100101101",
			179 => "1111111000001100101101",
			180 => "0000011101000000101000",
			181 => "0011010111011100100000",
			182 => "0000111101101000000100",
			183 => "0000010000001100101101",
			184 => "0011010110001100001100",
			185 => "0001011111011000000100",
			186 => "0000000000001100101101",
			187 => "0010010101010100000100",
			188 => "0000000000001100101101",
			189 => "1111111000001100101101",
			190 => "0011100011101100001000",
			191 => "0001000011000000000100",
			192 => "0000100000001100101101",
			193 => "0000000000001100101101",
			194 => "0010011001001000000100",
			195 => "1111111000001100101101",
			196 => "0000001000001100101101",
			197 => "0000001000010000000100",
			198 => "0000001000001100101101",
			199 => "0000100000001100101101",
			200 => "0001000110000000000100",
			201 => "0000000000001100101101",
			202 => "1111111000001100101101",
			203 => "0011011110011000101000",
			204 => "0000000100010100100000",
			205 => "0001011000000000010100",
			206 => "0000110011000000001100",
			207 => "0011100010010100000100",
			208 => "0000000000001111010001",
			209 => "0000000101011000000100",
			210 => "0000000000001111010001",
			211 => "0000000000001111010001",
			212 => "0001111000111000000100",
			213 => "0000000000001111010001",
			214 => "1111111000001111010001",
			215 => "0000111100110000001000",
			216 => "0001101001110000000100",
			217 => "0000000000001111010001",
			218 => "0000000000001111010001",
			219 => "0000000000001111010001",
			220 => "0000111111011000000100",
			221 => "0000000000001111010001",
			222 => "1111111000001111010001",
			223 => "0000100011111000001100",
			224 => "0001111001010100001000",
			225 => "0011100110100000000100",
			226 => "0000000000001111010001",
			227 => "0000000000001111010001",
			228 => "1111111000001111010001",
			229 => "0011100011101100000100",
			230 => "0000001000001111010001",
			231 => "0000001011100100001100",
			232 => "0011011100101000000100",
			233 => "0000000000001111010001",
			234 => "0001100101100000000100",
			235 => "0000000000001111010001",
			236 => "0000000000001111010001",
			237 => "0000110011100100000100",
			238 => "0000001000001111010001",
			239 => "0010010110000000000100",
			240 => "1111111000001111010001",
			241 => "0011000101011100000100",
			242 => "0000000000001111010001",
			243 => "0000000000001111010001",
			244 => "0010101111011000001100",
			245 => "0001111000000100000100",
			246 => "0000000000010001000101",
			247 => "0000000101011000000100",
			248 => "0000000000010001000101",
			249 => "0000001000010001000101",
			250 => "0010000011010000000100",
			251 => "1111111000010001000101",
			252 => "0010000101011100010100",
			253 => "0011001010100100001000",
			254 => "0010010101011100000100",
			255 => "0000000000010001000101",
			256 => "0000001000010001000101",
			257 => "0001111001010000001000",
			258 => "0000110101111000000100",
			259 => "0000000000010001000101",
			260 => "1111111000010001000101",
			261 => "0000001000010001000101",
			262 => "0011001110011000000100",
			263 => "1111111000010001000101",
			264 => "0010100011000100010000",
			265 => "0010110101011100001000",
			266 => "0011111001111000000100",
			267 => "0000000000010001000101",
			268 => "0000000000010001000101",
			269 => "0011011100101000000100",
			270 => "0000001000010001000101",
			271 => "0000000000010001000101",
			272 => "1111111000010001000101",
			273 => "0011110001100000010100",
			274 => "0011111000101100010000",
			275 => "0010010110000000001100",
			276 => "0010001001000100000100",
			277 => "1100011000010011001001",
			278 => "0000000111001000000100",
			279 => "1100011000010011001001",
			280 => "1100110000010011001001",
			281 => "1100011000010011001001",
			282 => "1100100000010011001001",
			283 => "0010101000000100000100",
			284 => "1111001000010011001001",
			285 => "0000110011001000001100",
			286 => "0001000111011100000100",
			287 => "1100100000010011001001",
			288 => "0010101100010000000100",
			289 => "1110001000010011001001",
			290 => "1101000000010011001001",
			291 => "0010001010000100011000",
			292 => "0011000101010100001100",
			293 => "0000111100110000001000",
			294 => "0010111010100100000100",
			295 => "1100100000010011001001",
			296 => "1100111000010011001001",
			297 => "1100011000010011001001",
			298 => "0001100100001000001000",
			299 => "0010110101010100000100",
			300 => "1101001000010011001001",
			301 => "1100011000010011001001",
			302 => "1110000000010011001001",
			303 => "0000011101000000000100",
			304 => "1100100000010011001001",
			305 => "1100011000010011001001",
			306 => "0000010011110001000000",
			307 => "0001010011001000010100",
			308 => "0010101111011000001100",
			309 => "0001101010001000001000",
			310 => "0000010110010000000100",
			311 => "0000000000010101101101",
			312 => "0000000000010101101101",
			313 => "0000000000010101101101",
			314 => "0001111001010000000100",
			315 => "0000000000010101101101",
			316 => "0000000000010101101101",
			317 => "0001000101010100001000",
			318 => "0010000101101100000100",
			319 => "0000000000010101101101",
			320 => "0000000000010101101101",
			321 => "0001000011000000010000",
			322 => "0011111011011000001100",
			323 => "0011010011010000001000",
			324 => "0000010001110000000100",
			325 => "0000000000010101101101",
			326 => "0000000000010101101101",
			327 => "0000000000010101101101",
			328 => "0000000000010101101101",
			329 => "0011010101010100010000",
			330 => "0011000101011100001000",
			331 => "0001001001010100000100",
			332 => "0000000000010101101101",
			333 => "0000000000010101101101",
			334 => "0010110101010100000100",
			335 => "0000000000010101101101",
			336 => "0000000000010101101101",
			337 => "0000000000010101101101",
			338 => "0011001001000100001100",
			339 => "0000110011001000001000",
			340 => "0000110011000000000100",
			341 => "0000000000010101101101",
			342 => "0000000000010101101101",
			343 => "0000000000010101101101",
			344 => "0010010011001000000100",
			345 => "0000000000010101101101",
			346 => "0000000000010101101101",
			347 => "0011111011011100101100",
			348 => "0010101000101000100000",
			349 => "0011001010100100001100",
			350 => "0001111000111000001000",
			351 => "0001110011001000000100",
			352 => "0000000000011000111001",
			353 => "0000000000011000111001",
			354 => "0000000000011000111001",
			355 => "0001011001010100001100",
			356 => "0000110110000000001000",
			357 => "0000111001000100000100",
			358 => "0000000000011000111001",
			359 => "0000000000011000111001",
			360 => "0000000000011000111001",
			361 => "0000111100010000000100",
			362 => "0000000000011000111001",
			363 => "0000000000011000111001",
			364 => "0000011000011000000100",
			365 => "0000000000011000111001",
			366 => "0010011010000100000100",
			367 => "0000000000011000111001",
			368 => "0000000000011000111001",
			369 => "0000010111100100011000",
			370 => "0001000101010100001000",
			371 => "0001011111011000000100",
			372 => "0000000000011000111001",
			373 => "0000000000011000111001",
			374 => "0000011001100100000100",
			375 => "0000000000011000111001",
			376 => "0000101111101100000100",
			377 => "0000000000011000111001",
			378 => "0011010110110100000100",
			379 => "0000000000011000111001",
			380 => "0000000000011000111001",
			381 => "0001001100101000001000",
			382 => "0011001010100100000100",
			383 => "0000000000011000111001",
			384 => "0000000000011000111001",
			385 => "0001001100000000010000",
			386 => "0010000101101100000100",
			387 => "0000000000011000111001",
			388 => "0010110101011100000100",
			389 => "0000000000011000111001",
			390 => "0000100100010100000100",
			391 => "0000000000011000111001",
			392 => "0000000000011000111001",
			393 => "0010010011001000001000",
			394 => "0001100100100000000100",
			395 => "0000000000011000111001",
			396 => "0000000000011000111001",
			397 => "0000000000011000111001",
			398 => "0010110101011100110100",
			399 => "0001110100101100101100",
			400 => "0000101111001100100100",
			401 => "0011101111010100011000",
			402 => "0011101101100000010000",
			403 => "0010110011010000001000",
			404 => "0001000110000000000100",
			405 => "0000000000011011011101",
			406 => "0000000000011011011101",
			407 => "0001010011000100000100",
			408 => "0000000000011011011101",
			409 => "0000000000011011011101",
			410 => "0001101110001000000100",
			411 => "1111111000011011011101",
			412 => "0000000000011011011101",
			413 => "0000010110010000000100",
			414 => "0000000000011011011101",
			415 => "0000101100100100000100",
			416 => "0000000000011011011101",
			417 => "0000001000011011011101",
			418 => "0011001010100100000100",
			419 => "0000000000011011011101",
			420 => "0000000000011011011101",
			421 => "0000001010010000000100",
			422 => "1111111000011011011101",
			423 => "0000000000011011011101",
			424 => "0011011100101000011000",
			425 => "0010101011000000010000",
			426 => "0010010011001000001100",
			427 => "0010010110000000000100",
			428 => "0000000000011011011101",
			429 => "0000000001110100000100",
			430 => "0000000000011011011101",
			431 => "0000001000011011011101",
			432 => "0000000000011011011101",
			433 => "0001110011000100000100",
			434 => "0000000000011011011101",
			435 => "0000000000011011011101",
			436 => "0000011001100000000100",
			437 => "0000000000011011011101",
			438 => "0000000000011011011101",
			439 => "0011110111100000010100",
			440 => "0010010110000000010000",
			441 => "0011001100101000001100",
			442 => "0000000100011000000100",
			443 => "1111111000011101010001",
			444 => "0010101001010100000100",
			445 => "0000001000011101010001",
			446 => "1111111000011101010001",
			447 => "0000001000011101010001",
			448 => "1111111000011101010001",
			449 => "0000010110001100100100",
			450 => "0001101110100100000100",
			451 => "0000010000011101010001",
			452 => "0000000111110100000100",
			453 => "1111111000011101010001",
			454 => "0000111001010100010000",
			455 => "0010010101011100001000",
			456 => "0000000100010100000100",
			457 => "0000001000011101010001",
			458 => "1111111000011101010001",
			459 => "0000010001110000000100",
			460 => "0000000000011101010001",
			461 => "0000001000011101010001",
			462 => "0000000101101000000100",
			463 => "1111111000011101010001",
			464 => "0010110111011100000100",
			465 => "1111111000011101010001",
			466 => "0000001000011101010001",
			467 => "1111111000011101010001",
			468 => "0011111110000000000100",
			469 => "1111111000011110100101",
			470 => "0001011100011100100100",
			471 => "0000010110001100100000",
			472 => "0001101110100000001100",
			473 => "0001111100110000001000",
			474 => "0000010001110000000100",
			475 => "0000010000011110100101",
			476 => "0000001000011110100101",
			477 => "1111111000011110100101",
			478 => "0010110101011100010000",
			479 => "0001110100101100001000",
			480 => "0000101111001100000100",
			481 => "0000000000011110100101",
			482 => "1111111000011110100101",
			483 => "0000101111001100000100",
			484 => "1111111000011110100101",
			485 => "0000000000011110100101",
			486 => "0000001000011110100101",
			487 => "1111111000011110100101",
			488 => "1111111000011110100101",
			489 => "0011111000101100010000",
			490 => "0010010110000000001100",
			491 => "0010001001000100000100",
			492 => "1111111000100000110001",
			493 => "0011110010001100000100",
			494 => "1111111000100000110001",
			495 => "0000010000100000110001",
			496 => "1111111000100000110001",
			497 => "0000010110001100110100",
			498 => "0000110011001000010100",
			499 => "0000000101011000000100",
			500 => "1111111000100000110001",
			501 => "0010010101011100001000",
			502 => "0010101000000000000100",
			503 => "0000010000100000110001",
			504 => "1111111000100000110001",
			505 => "0001000111011100000100",
			506 => "0000010000100000110001",
			507 => "0000100000100000110001",
			508 => "0011011110011000001100",
			509 => "0000011000011000001000",
			510 => "0001011000000100000100",
			511 => "0000000000100000110001",
			512 => "1111111000100000110001",
			513 => "0000010000100000110001",
			514 => "0000000101101000001000",
			515 => "0001111000101000000100",
			516 => "0000100000100000110001",
			517 => "1111111000100000110001",
			518 => "0010111010100100000100",
			519 => "1111111000100000110001",
			520 => "0010001010000100000100",
			521 => "0000101000100000110001",
			522 => "0000001000100000110001",
			523 => "1111111000100000110001",
			524 => "0001001001010001000000",
			525 => "0010110101011100101000",
			526 => "0001011011000000011100",
			527 => "0010011101101000011000",
			528 => "0011010111011100010000",
			529 => "0000000100010100001000",
			530 => "0001000011000000000100",
			531 => "0000000000100010110101",
			532 => "1111111000100010110101",
			533 => "0001101101010000000100",
			534 => "0000000000100010110101",
			535 => "0000000000100010110101",
			536 => "0000000111101100000100",
			537 => "0000000000100010110101",
			538 => "0000000000100010110101",
			539 => "1111111000100010110101",
			540 => "0011000101010100000100",
			541 => "1111111000100010110101",
			542 => "0010001111001000000100",
			543 => "0000001000100010110101",
			544 => "0000000000100010110101",
			545 => "0010101011000000001100",
			546 => "0010010011001000001000",
			547 => "0011111100111100000100",
			548 => "0000000000100010110101",
			549 => "0000001000100010110101",
			550 => "1111111000100010110101",
			551 => "0011001001000100000100",
			552 => "1111111000100010110101",
			553 => "0011000110000000000100",
			554 => "0000001000100010110101",
			555 => "0000000000100010110101",
			556 => "1111111000100010110101",
			557 => "0011110100011001000100",
			558 => "0001111100110000011100",
			559 => "0000001001110100010100",
			560 => "0001000110000000001000",
			561 => "0000000100011000000100",
			562 => "0000000000100110010001",
			563 => "0000000000100110010001",
			564 => "0011001100101000000100",
			565 => "0000000000100110010001",
			566 => "0000101000110100000100",
			567 => "0000000000100110010001",
			568 => "0000000000100110010001",
			569 => "0011100011010100000100",
			570 => "0000000000100110010001",
			571 => "0000000000100110010001",
			572 => "0001001010000100001100",
			573 => "0000110110000000001000",
			574 => "0000110101101100000100",
			575 => "0000000000100110010001",
			576 => "0000000000100110010001",
			577 => "1111111000100110010001",
			578 => "0000101010101000010000",
			579 => "0010110111011100000100",
			580 => "0000000000100110010001",
			581 => "0000010011110000000100",
			582 => "0000000000100110010001",
			583 => "0000011101000000000100",
			584 => "0000000000100110010001",
			585 => "0000000000100110010001",
			586 => "0000100010101100000100",
			587 => "0000000000100110010001",
			588 => "0001001000111000000100",
			589 => "0000000000100110010001",
			590 => "0000000000100110010001",
			591 => "0011111001111000001100",
			592 => "0001000011000000001000",
			593 => "0010011100101000000100",
			594 => "0000000000100110010001",
			595 => "0000000000100110010001",
			596 => "0000000000100110010001",
			597 => "0010011101101000010000",
			598 => "0000111000000000001100",
			599 => "0011110010101000000100",
			600 => "0000000000100110010001",
			601 => "0000010110010000000100",
			602 => "0000000000100110010001",
			603 => "0000000000100110010001",
			604 => "0000000000100110010001",
			605 => "0000011101000000000100",
			606 => "0000000000100110010001",
			607 => "0000001101111000000100",
			608 => "0000000000100110010001",
			609 => "0000101101011000000100",
			610 => "0000000000100110010001",
			611 => "0000000000100110010001",
			612 => "0011111011011100111100",
			613 => "0001011000111000100000",
			614 => "0001111000111000010100",
			615 => "0001010011001000001100",
			616 => "0001001011101100001000",
			617 => "0001010101101100000100",
			618 => "0000000000101001110101",
			619 => "0000000000101001110101",
			620 => "0000000000101001110101",
			621 => "0011001010100100000100",
			622 => "0000000000101001110101",
			623 => "0000000000101001110101",
			624 => "0010100011000000001000",
			625 => "0001001011101100000100",
			626 => "0000000000101001110101",
			627 => "0000000000101001110101",
			628 => "0000000000101001110101",
			629 => "0001000011000000010000",
			630 => "0010111110011000000100",
			631 => "0000000000101001110101",
			632 => "0011110001100000001000",
			633 => "0001011100110000000100",
			634 => "0000000000101001110101",
			635 => "0000000000101001110101",
			636 => "0000000000101001110101",
			637 => "0011100101110000001000",
			638 => "0000101000110100000100",
			639 => "0000000000101001110101",
			640 => "0000000000101001110101",
			641 => "0000000000101001110101",
			642 => "0011010111011100101000",
			643 => "0000100110010100001000",
			644 => "0001111000101000000100",
			645 => "0000000000101001110101",
			646 => "0000000000101001110101",
			647 => "0001101010101100010000",
			648 => "0000010111110000001100",
			649 => "0010001001001100000100",
			650 => "0000000000101001110101",
			651 => "0000010001110000000100",
			652 => "0000000000101001110101",
			653 => "0000000000101001110101",
			654 => "0000000000101001110101",
			655 => "0000101101111000001000",
			656 => "0011101010001000000100",
			657 => "0000000000101001110101",
			658 => "0000000000101001110101",
			659 => "0001110001010000000100",
			660 => "0000000000101001110101",
			661 => "0000000000101001110101",
			662 => "0001011101001000000100",
			663 => "0000000000101001110101",
			664 => "0001001100000000000100",
			665 => "0000000000101001110101",
			666 => "0010010011001000000100",
			667 => "0000000000101001110101",
			668 => "0000000000101001110101",
			669 => "0001001100101000100100",
			670 => "0000110011000000011000",
			671 => "0001111000000100000100",
			672 => "0000000000101101001001",
			673 => "0010000101101100001000",
			674 => "0000000101011000000100",
			675 => "0000000000101101001001",
			676 => "0000001000101101001001",
			677 => "0000110101101100001000",
			678 => "0010101111111100000100",
			679 => "0000000000101101001001",
			680 => "0000000000101101001001",
			681 => "0000000000101101001001",
			682 => "0011001010100100001000",
			683 => "0010010101011100000100",
			684 => "0000000000101101001001",
			685 => "0000000000101101001001",
			686 => "1111111000101101001001",
			687 => "0010101000111000011000",
			688 => "0000011001100000010000",
			689 => "0010011001000100001100",
			690 => "0001010011001000000100",
			691 => "0000000000101101001001",
			692 => "0001101001110000000100",
			693 => "0000000000101101001001",
			694 => "0000001000101101001001",
			695 => "0000000000101101001001",
			696 => "0010110111011100000100",
			697 => "0000000000101101001001",
			698 => "0000000000101101001001",
			699 => "0001011100110000001100",
			700 => "0010111110011000000100",
			701 => "0000000000101101001001",
			702 => "0010110101010100000100",
			703 => "1111111000101101001001",
			704 => "0000000000101101001001",
			705 => "0010101011000000010100",
			706 => "0011011110011000001000",
			707 => "0000010111100100000100",
			708 => "1111111000101101001001",
			709 => "0000000000101101001001",
			710 => "0000010111100100000100",
			711 => "0000001000101101001001",
			712 => "0001111000101000000100",
			713 => "0000000000101101001001",
			714 => "0000000000101101001001",
			715 => "0010000101011100001000",
			716 => "0000010111110000000100",
			717 => "0000000000101101001001",
			718 => "0000000000101101001001",
			719 => "0011110011100000000100",
			720 => "1111111000101101001001",
			721 => "0000000000101101001001",
			722 => "0010101011111001000000",
			723 => "0011000101011100101100",
			724 => "0001000011000000101000",
			725 => "0001011100110000010000",
			726 => "0001000110000000001100",
			727 => "0010101101001000001000",
			728 => "0010110111011100000100",
			729 => "0000000000101111101101",
			730 => "0000000000101111101101",
			731 => "0000000000101111101101",
			732 => "1111111000101111101101",
			733 => "0011111001111000001100",
			734 => "0001111100010000000100",
			735 => "0000000000101111101101",
			736 => "0001001010000100000100",
			737 => "0000000000101111101101",
			738 => "0000001000101111101101",
			739 => "0010001111111100001000",
			740 => "0011100001000100000100",
			741 => "0000000000101111101101",
			742 => "0000000000101111101101",
			743 => "0000000000101111101101",
			744 => "1111111000101111101101",
			745 => "0010101111101000001100",
			746 => "0001110100101100000100",
			747 => "0000000000101111101101",
			748 => "0010000011001000000100",
			749 => "0000000000101111101101",
			750 => "0000000000101111101101",
			751 => "0000011101000000000100",
			752 => "0000001000101111101101",
			753 => "0000000000101111101101",
			754 => "0001001100010000000100",
			755 => "0000000000101111101101",
			756 => "0001001001010000001100",
			757 => "0001111001010000000100",
			758 => "0000000000101111101101",
			759 => "0000011110011000000100",
			760 => "0000000000101111101101",
			761 => "0000000000101111101101",
			762 => "0000000000101111101101",
			763 => "0001011100110001000000",
			764 => "0010101000111000101000",
			765 => "0011111011011100100000",
			766 => "0011001010100100001100",
			767 => "0001110011001000000100",
			768 => "0000000000110011011001",
			769 => "0001111000111000000100",
			770 => "0000000000110011011001",
			771 => "0000000000110011011001",
			772 => "0001110011001000001000",
			773 => "0000000101000000000100",
			774 => "0000000000110011011001",
			775 => "0000000000110011011001",
			776 => "0010100101101100001000",
			777 => "0000111100101000000100",
			778 => "0000000000110011011001",
			779 => "0000000000110011011001",
			780 => "0000000000110011011001",
			781 => "0001000111011100000100",
			782 => "0000000000110011011001",
			783 => "0000000000110011011001",
			784 => "0000010001100100001100",
			785 => "0001010101111000001000",
			786 => "0010111010100100000100",
			787 => "0000000000110011011001",
			788 => "0000000000110011011001",
			789 => "0000000000110011011001",
			790 => "0000110011100100000100",
			791 => "0000000000110011011001",
			792 => "0000111101001000000100",
			793 => "0000000000110011011001",
			794 => "0000000000110011011001",
			795 => "0010101011111000100100",
			796 => "0010110011010000010000",
			797 => "0000011000011000001000",
			798 => "0000001011001000000100",
			799 => "0000000000110011011001",
			800 => "0000000000110011011001",
			801 => "0010101001010100000100",
			802 => "0000000000110011011001",
			803 => "0000000000110011011001",
			804 => "0000010111100100000100",
			805 => "0000000000110011011001",
			806 => "0010110111011100000100",
			807 => "0000000000110011011001",
			808 => "0001111000101000000100",
			809 => "0000000000110011011001",
			810 => "0011100110111000000100",
			811 => "0000000000110011011001",
			812 => "0000000000110011011001",
			813 => "0011001001000100001100",
			814 => "0001001001010100000100",
			815 => "0000000000110011011001",
			816 => "0001001111101000000100",
			817 => "0000000000110011011001",
			818 => "0000000000110011011001",
			819 => "0010011000000100000100",
			820 => "0000000000110011011001",
			821 => "0000000000110011011001",
			822 => "0010110101011101000100",
			823 => "0010011001000100101100",
			824 => "0001110001010000100000",
			825 => "0000001111001100011100",
			826 => "0011111011011100010000",
			827 => "0001011001010100001000",
			828 => "0011001010100100000100",
			829 => "0000000000110110010101",
			830 => "0000000000110110010101",
			831 => "0001111100010000000100",
			832 => "0000000000110110010101",
			833 => "0000000000110110010101",
			834 => "0000001100100100000100",
			835 => "0000001000110110010101",
			836 => "0010101101001000000100",
			837 => "0000000000110110010101",
			838 => "0000000000110110010101",
			839 => "1111111000110110010101",
			840 => "0000111000000000001000",
			841 => "0001101000010100000100",
			842 => "0000000000110110010101",
			843 => "0000001000110110010101",
			844 => "0000000000110110010101",
			845 => "0001011011111000001000",
			846 => "0010000101011100000100",
			847 => "0000000000110110010101",
			848 => "1111111000110110010101",
			849 => "0001011100011100001100",
			850 => "0000011101000000001000",
			851 => "0010011101101000000100",
			852 => "0000000000110110010101",
			853 => "0000000000110110010101",
			854 => "0000000000110110010101",
			855 => "0000000000110110010101",
			856 => "0010010011001000011000",
			857 => "0010101011000000001000",
			858 => "0011111100111100000100",
			859 => "0000000000110110010101",
			860 => "0000000000110110010101",
			861 => "0000011001100000001000",
			862 => "0000010111100100000100",
			863 => "0000000000110110010101",
			864 => "0000000000110110010101",
			865 => "0010001010000100000100",
			866 => "0000000000110110010101",
			867 => "0000000000110110010101",
			868 => "0000000000110110010101",
			869 => "0000000110001000001100",
			870 => "0001111000000000001000",
			871 => "0011100100000000000100",
			872 => "1111111000111000100001",
			873 => "0000001000111000100001",
			874 => "1111111000111000100001",
			875 => "0000101110011100000100",
			876 => "0000010000111000100001",
			877 => "0000010011110000100000",
			878 => "0011010101010100011000",
			879 => "0000000100010100001100",
			880 => "0001111000101000001000",
			881 => "0000011000011000000100",
			882 => "0000000000111000100001",
			883 => "0000001000111000100001",
			884 => "1111111000111000100001",
			885 => "0011100010110000000100",
			886 => "1111111000111000100001",
			887 => "0000011001100000000100",
			888 => "0000000000111000100001",
			889 => "1111111000111000100001",
			890 => "0000100111110100000100",
			891 => "0000000000111000100001",
			892 => "0000001000111000100001",
			893 => "0000111100010000001100",
			894 => "0000001101011100000100",
			895 => "0000000000111000100001",
			896 => "0001011101001000000100",
			897 => "0000001000111000100001",
			898 => "1111111000111000100001",
			899 => "0011001001000100000100",
			900 => "1111111000111000100001",
			901 => "0010110101101100000100",
			902 => "0000001000111000100001",
			903 => "1111111000111000100001",
			904 => "0011111010110000110100",
			905 => "0011100001101100100100",
			906 => "0011100000110100011000",
			907 => "0000001101110100010100",
			908 => "0010011001001000001000",
			909 => "0011110100010000000100",
			910 => "0000000000111100000101",
			911 => "0000000000111100000101",
			912 => "0011101101101100001000",
			913 => "0001101111000000000100",
			914 => "0000000000111100000101",
			915 => "0000000000111100000101",
			916 => "1111111000111100000101",
			917 => "1111111000111100000101",
			918 => "0000011001100000001000",
			919 => "0000010001110000000100",
			920 => "0000000000111100000101",
			921 => "0000001000111100000101",
			922 => "0000000000111100000101",
			923 => "0000010001100100001000",
			924 => "0001000101010100000100",
			925 => "0000000000111100000101",
			926 => "1111111000111100000101",
			927 => "0000100011111000000100",
			928 => "0000000000111100000101",
			929 => "0000000000111100000101",
			930 => "0011011110011000011000",
			931 => "0000000100010100001100",
			932 => "0011110111010000000100",
			933 => "0000000000111100000101",
			934 => "0001111001010000000100",
			935 => "0000001000111100000101",
			936 => "0000000000111100000101",
			937 => "0011110101000100000100",
			938 => "1111111000111100000101",
			939 => "0011111110011100000100",
			940 => "0000000000111100000101",
			941 => "0000000000111100000101",
			942 => "0000011001100000001100",
			943 => "0001001001000100000100",
			944 => "0000000000111100000101",
			945 => "0000010111100100000100",
			946 => "0000001000111100000101",
			947 => "0000000000111100000101",
			948 => "0010101101001000000100",
			949 => "0000000000111100000101",
			950 => "0011100001000000001000",
			951 => "0011110111000000000100",
			952 => "0000000000111100000101",
			953 => "1111111000111100000101",
			954 => "0001001100000000001000",
			955 => "0000111100010000000100",
			956 => "0000000000111100000101",
			957 => "0000000000111100000101",
			958 => "0010111001001000000100",
			959 => "0000000000111100000101",
			960 => "0000000000111100000101",
			961 => "0011111010110000111000",
			962 => "0011100001101100101000",
			963 => "0001011000000000010000",
			964 => "0011100000110100001100",
			965 => "0001001101000000001000",
			966 => "0001011001001000000100",
			967 => "0000000000111111101001",
			968 => "0000000000111111101001",
			969 => "1111111000111111101001",
			970 => "0000000000111111101001",
			971 => "0001001111011000010100",
			972 => "0011010011010000001100",
			973 => "0001011000101000001000",
			974 => "0000000100011000000100",
			975 => "0000000000111111101001",
			976 => "0000001000111111101001",
			977 => "0000000000111111101001",
			978 => "0001011001010100000100",
			979 => "0000000000111111101001",
			980 => "0000000000111111101001",
			981 => "0000000000111111101001",
			982 => "0000010001100100001000",
			983 => "0001000101010100000100",
			984 => "0000000000111111101001",
			985 => "1111111000111111101001",
			986 => "0000100011111000000100",
			987 => "0000000000111111101001",
			988 => "0000000000111111101001",
			989 => "0000010111100100010100",
			990 => "0011011110011000010000",
			991 => "0000111000000000001100",
			992 => "0001101101010000001000",
			993 => "0000001100100100000100",
			994 => "0000000000111111101001",
			995 => "1111111000111111101001",
			996 => "0000000000111111101001",
			997 => "1111111000111111101001",
			998 => "0000000000111111101001",
			999 => "0010110101011100011000",
			1000 => "0000010001100100010000",
			1001 => "0010001111001000001100",
			1002 => "0000101011111100000100",
			1003 => "0000000000111111101001",
			1004 => "0000101111001100000100",
			1005 => "1111111000111111101001",
			1006 => "0000000000111111101001",
			1007 => "0000000000111111101001",
			1008 => "0010001111001000000100",
			1009 => "0000000000111111101001",
			1010 => "1111111000111111101001",
			1011 => "0011011100101000000100",
			1012 => "0000000000111111101001",
			1013 => "0000000100010100001000",
			1014 => "0011111101010100000100",
			1015 => "0000000000111111101001",
			1016 => "0000000000111111101001",
			1017 => "0000000000111111101001",
			1018 => "0001101100000100101100",
			1019 => "0000101010101000100100",
			1020 => "0001111001010100100000",
			1021 => "0011100000110100011100",
			1022 => "0011001010100100001100",
			1023 => "0010101000111000001000",
			1024 => "0000101000110100000100",
			1025 => "0000000001000010100101",
			1026 => "0000000001000010100101",
			1027 => "0000000001000010100101",
			1028 => "0011101101101100001000",
			1029 => "0011110000010100000100",
			1030 => "0000000001000010100101",
			1031 => "0000000001000010100101",
			1032 => "0001011001010100000100",
			1033 => "0000000001000010100101",
			1034 => "0000000001000010100101",
			1035 => "0000000001000010100101",
			1036 => "0000000001000010100101",
			1037 => "0001001000000000000100",
			1038 => "0000000001000010100101",
			1039 => "0000000001000010100101",
			1040 => "0011011110011000010100",
			1041 => "0000001100100100001000",
			1042 => "0000000010101100000100",
			1043 => "0000000001000010100101",
			1044 => "0000000001000010100101",
			1045 => "0001101101010000000100",
			1046 => "0000000001000010100101",
			1047 => "0011110011111100000100",
			1048 => "0000000001000010100101",
			1049 => "0000000001000010100101",
			1050 => "0000011001100000001000",
			1051 => "0011100111100000000100",
			1052 => "0000000001000010100101",
			1053 => "0000000001000010100101",
			1054 => "0000010001100100000100",
			1055 => "0000000001000010100101",
			1056 => "0000101111001100001100",
			1057 => "0001101011011100001000",
			1058 => "0010101011000000000100",
			1059 => "0000000001000010100101",
			1060 => "0000000001000010100101",
			1061 => "0000000001000010100101",
			1062 => "0011110011100000000100",
			1063 => "0000000001000010100101",
			1064 => "0000000001000010100101",
			1065 => "0010101000111000100100",
			1066 => "0001010011001000010000",
			1067 => "0000110011000000001100",
			1068 => "0001111000000100000100",
			1069 => "0000000001000110010001",
			1070 => "0000000101011000000100",
			1071 => "0000000001000110010001",
			1072 => "0000000001000110010001",
			1073 => "0000000001000110010001",
			1074 => "0000110011100100010000",
			1075 => "0000011001100000001100",
			1076 => "0001000110000000001000",
			1077 => "0001001100101000000100",
			1078 => "0000000001000110010001",
			1079 => "0000001001000110010001",
			1080 => "0000000001000110010001",
			1081 => "0000000001000110010001",
			1082 => "0000000001000110010001",
			1083 => "0010110111011100101000",
			1084 => "0000011000011000010100",
			1085 => "0000001011001000001000",
			1086 => "0011110001100000000100",
			1087 => "0000000001000110010001",
			1088 => "0000000001000110010001",
			1089 => "0010110011010000001000",
			1090 => "0000011001100100000100",
			1091 => "0000000001000110010001",
			1092 => "1111111001000110010001",
			1093 => "0000000001000110010001",
			1094 => "0010111110011000000100",
			1095 => "0000000001000110010001",
			1096 => "0011011010100100001000",
			1097 => "0001111000101000000100",
			1098 => "0000000001000110010001",
			1099 => "0000000001000110010001",
			1100 => "0001001001001000000100",
			1101 => "0000000001000110010001",
			1102 => "0000000001000110010001",
			1103 => "0010101011111000011000",
			1104 => "0001011100010000000100",
			1105 => "0000000001000110010001",
			1106 => "0011010101011100001000",
			1107 => "0001100000100000000100",
			1108 => "0000000001000110010001",
			1109 => "0000000001000110010001",
			1110 => "0011110100110100000100",
			1111 => "0000000001000110010001",
			1112 => "0011100111101000000100",
			1113 => "0000000001000110010001",
			1114 => "0000000001000110010001",
			1115 => "0011001001000100001100",
			1116 => "0010000101011100001000",
			1117 => "0000010111110000000100",
			1118 => "0000000001000110010001",
			1119 => "0000000001000110010001",
			1120 => "0000000001000110010001",
			1121 => "0010111001001000000100",
			1122 => "0000000001000110010001",
			1123 => "0000000001000110010001",
			1124 => "0011010111011101001000",
			1125 => "0010101111011000001100",
			1126 => "0001111000000100000100",
			1127 => "0000000001001001010101",
			1128 => "0000000101011000000100",
			1129 => "0000000001001001010101",
			1130 => "0000000001001001010101",
			1131 => "0011000101011100110000",
			1132 => "0010001111111100011000",
			1133 => "0011010110001100001100",
			1134 => "0011110101000100001000",
			1135 => "0000000101011000000100",
			1136 => "0000000001001001010101",
			1137 => "0000000001001001010101",
			1138 => "0000000001001001010101",
			1139 => "0001011001010000001000",
			1140 => "0010001001001100000100",
			1141 => "0000000001001001010101",
			1142 => "0000000001001001010101",
			1143 => "0000000001001001010101",
			1144 => "0000000110111100001100",
			1145 => "0001011000000000000100",
			1146 => "0000000001001001010101",
			1147 => "0001111000101000000100",
			1148 => "0000000001001001010101",
			1149 => "0000000001001001010101",
			1150 => "0011110100110100000100",
			1151 => "0000000001001001010101",
			1152 => "0001101100111100000100",
			1153 => "0000000001001001010101",
			1154 => "0000000001001001010101",
			1155 => "0001011000101000000100",
			1156 => "0000000001001001010101",
			1157 => "0001001000000000000100",
			1158 => "0000000001001001010101",
			1159 => "0000000001001001010101",
			1160 => "0000011111011100010000",
			1161 => "0000001000010000001100",
			1162 => "0001110110101100001000",
			1163 => "0001111100110000000100",
			1164 => "0000000001001001010101",
			1165 => "0000000001001001010101",
			1166 => "0000000001001001010101",
			1167 => "0000000001001001010101",
			1168 => "0000110011001000001000",
			1169 => "0010010101111000000100",
			1170 => "0000000001001001010101",
			1171 => "0000000001001001010101",
			1172 => "0000000001001001010101",
			1173 => "0011100100100100010000",
			1174 => "0010001111001000000100",
			1175 => "1111111001001100010001",
			1176 => "0010001010000100001000",
			1177 => "0000001010111100000100",
			1178 => "0000000001001100010001",
			1179 => "0000001001001100010001",
			1180 => "1111111001001100010001",
			1181 => "0000111000000000101100",
			1182 => "0011001010100100010100",
			1183 => "0010101101001000010000",
			1184 => "0011111001111000001100",
			1185 => "0000001001110100001000",
			1186 => "0000000100110100000100",
			1187 => "0000000001001100010001",
			1188 => "0000001001001100010001",
			1189 => "0000000001001100010001",
			1190 => "0000001001001100010001",
			1191 => "1111111001001100010001",
			1192 => "0000001001110100001000",
			1193 => "0001001010100100000100",
			1194 => "0000000001001100010001",
			1195 => "1111111001001100010001",
			1196 => "0011010111011100001100",
			1197 => "0000101011010000000100",
			1198 => "0000000001001100010001",
			1199 => "0001111001010100000100",
			1200 => "1111111001001100010001",
			1201 => "0000000001001100010001",
			1202 => "0000001001001100010001",
			1203 => "0010110011010000001000",
			1204 => "0000001011001000000100",
			1205 => "0000001001001100010001",
			1206 => "1111111001001100010001",
			1207 => "0001111000101000001000",
			1208 => "0001011000100000000100",
			1209 => "0000001001001100010001",
			1210 => "1111111001001100010001",
			1211 => "0010000101101100000100",
			1212 => "0000001001001100010001",
			1213 => "0010111100101000001000",
			1214 => "0010010101111000000100",
			1215 => "1111111001001100010001",
			1216 => "0000000001001100010001",
			1217 => "0010010011001000000100",
			1218 => "0000001001001100010001",
			1219 => "1111111001001100010001",
			1220 => "0010110101011101001100",
			1221 => "0010101111011000001000",
			1222 => "0011100010010100000100",
			1223 => "0000000001001111001101",
			1224 => "0000000001001111001101",
			1225 => "0011101101100000100100",
			1226 => "0001011000000000001100",
			1227 => "0011011110011000001000",
			1228 => "0000110011000000000100",
			1229 => "0000000001001111001101",
			1230 => "0000000001001111001101",
			1231 => "0000000001001111001101",
			1232 => "0001000011000000001100",
			1233 => "0011111001111000001000",
			1234 => "0001011000101000000100",
			1235 => "0000000001001111001101",
			1236 => "0000000001001111001101",
			1237 => "0000000001001111001101",
			1238 => "0001011100101100000100",
			1239 => "0000000001001111001101",
			1240 => "0000011000011000000100",
			1241 => "0000000001001111001101",
			1242 => "0000000001001111001101",
			1243 => "0011011011101100001100",
			1244 => "0011110101000100000100",
			1245 => "0000000001001111001101",
			1246 => "0000111000000000000100",
			1247 => "0000000001001111001101",
			1248 => "0000000001001111001101",
			1249 => "0001011011111000001100",
			1250 => "0000010001100100000100",
			1251 => "0000000001001111001101",
			1252 => "0011110100111100000100",
			1253 => "0000000001001111001101",
			1254 => "0000000001001111001101",
			1255 => "0011000101011100000100",
			1256 => "0000000001001111001101",
			1257 => "0000000001001111001101",
			1258 => "0010010011001000010000",
			1259 => "0010101011000000001000",
			1260 => "0011111100111100000100",
			1261 => "0000000001001111001101",
			1262 => "0000000001001111001101",
			1263 => "0000011001100000000100",
			1264 => "0000000001001111001101",
			1265 => "0000000001001111001101",
			1266 => "0000000001001111001101",
			1267 => "0000000110001000001100",
			1268 => "0011111110000000000100",
			1269 => "1111111001010001110001",
			1270 => "0011101111100100000100",
			1271 => "0000001001010001110001",
			1272 => "1111111001010001110001",
			1273 => "0000111000000000100000",
			1274 => "0011010111011100011100",
			1275 => "0000001011010000001000",
			1276 => "0010101000111000000100",
			1277 => "0000001001010001110001",
			1278 => "0000000001010001110001",
			1279 => "0011100101110100000100",
			1280 => "1111111001010001110001",
			1281 => "0001101101010000001000",
			1282 => "0000001011001100000100",
			1283 => "0000001001010001110001",
			1284 => "1111111001010001110001",
			1285 => "0011110011111100000100",
			1286 => "0000001001010001110001",
			1287 => "1111111001010001110001",
			1288 => "0000001001010001110001",
			1289 => "0010010011001000100100",
			1290 => "0010110111011100010000",
			1291 => "0000000100010100001100",
			1292 => "0010101111101000001000",
			1293 => "0010111110011000000100",
			1294 => "1111111001010001110001",
			1295 => "0000001001010001110001",
			1296 => "1111111001010001110001",
			1297 => "1111111001010001110001",
			1298 => "0000011101000000001100",
			1299 => "0010101011111000000100",
			1300 => "0000001001010001110001",
			1301 => "0011010111011100000100",
			1302 => "1111111001010001110001",
			1303 => "0000001001010001110001",
			1304 => "0001001000111000000100",
			1305 => "1111111001010001110001",
			1306 => "0000000001010001110001",
			1307 => "1111111001010001110001",
			1308 => "0010101000111000101000",
			1309 => "0011111011011100100000",
			1310 => "0001111000111000010100",
			1311 => "0001111111011000000100",
			1312 => "0000000001010101001101",
			1313 => "0011001010100100000100",
			1314 => "0000000001010101001101",
			1315 => "0000011000011000000100",
			1316 => "0000000001010101001101",
			1317 => "0010001111001000000100",
			1318 => "0000000001010101001101",
			1319 => "0000000001010101001101",
			1320 => "0000110110000000001000",
			1321 => "0001010101101100000100",
			1322 => "0000000001010101001101",
			1323 => "0000000001010101001101",
			1324 => "0000000001010101001101",
			1325 => "0011010110001100000100",
			1326 => "0000000001010101001101",
			1327 => "0000000001010101001101",
			1328 => "0011010111011100100100",
			1329 => "0001011011000000011100",
			1330 => "0000001000110000011000",
			1331 => "0000010001100100010000",
			1332 => "0001011000000100001000",
			1333 => "0011111001111000000100",
			1334 => "0000000001010101001101",
			1335 => "0000000001010101001101",
			1336 => "0011110010010000000100",
			1337 => "0000000001010101001101",
			1338 => "1111111001010101001101",
			1339 => "0001100101100000000100",
			1340 => "0000000001010101001101",
			1341 => "0000000001010101001101",
			1342 => "0000000001010101001101",
			1343 => "0001010011000100000100",
			1344 => "0000000001010101001101",
			1345 => "0000000001010101001101",
			1346 => "0000011001100000001000",
			1347 => "0011100101110100000100",
			1348 => "0000000001010101001101",
			1349 => "0000000001010101001101",
			1350 => "0001011000000000000100",
			1351 => "0000000001010101001101",
			1352 => "0001111001010000001000",
			1353 => "0000001000001000000100",
			1354 => "0000000001010101001101",
			1355 => "0000000001010101001101",
			1356 => "0011000110000000001000",
			1357 => "0001110001001000000100",
			1358 => "0000000001010101001101",
			1359 => "0000000001010101001101",
			1360 => "0011011100101000000100",
			1361 => "0000000001010101001101",
			1362 => "0000000001010101001101",
			1363 => "0001000011000001011100",
			1364 => "0001001001000100111000",
			1365 => "0011010111011100101000",
			1366 => "0011001010100100010100",
			1367 => "0000011001100000010000",
			1368 => "0010010101011100001000",
			1369 => "0010101111011000000100",
			1370 => "0000000001011000101001",
			1371 => "1111111001011000101001",
			1372 => "0010000101101100000100",
			1373 => "0000001001011000101001",
			1374 => "0000000001011000101001",
			1375 => "1111111001011000101001",
			1376 => "0001111100101100010000",
			1377 => "0000110011000000001000",
			1378 => "0011100000110100000100",
			1379 => "0000000001011000101001",
			1380 => "0000001001011000101001",
			1381 => "0000011001100000000100",
			1382 => "1111111001011000101001",
			1383 => "0000000001011000101001",
			1384 => "0000000001011000101001",
			1385 => "0011010101010100001000",
			1386 => "0010001001000100000100",
			1387 => "0000000001011000101001",
			1388 => "0000001001011000101001",
			1389 => "0011001001001000000100",
			1390 => "0000000001011000101001",
			1391 => "0000000001011000101001",
			1392 => "0000101010010100011100",
			1393 => "0010110111011100010000",
			1394 => "0010011001000100001100",
			1395 => "0010101000111000000100",
			1396 => "0000001001011000101001",
			1397 => "0010001001001100000100",
			1398 => "1111111001011000101001",
			1399 => "0000000001011000101001",
			1400 => "1111111001011000101001",
			1401 => "0001110100101100001000",
			1402 => "0010011010000100000100",
			1403 => "0000001001011000101001",
			1404 => "0000000001011000101001",
			1405 => "0000000001011000101001",
			1406 => "0010111001001000000100",
			1407 => "1111111001011000101001",
			1408 => "0000000001011000101001",
			1409 => "0010010110000000000100",
			1410 => "1111111001011000101001",
			1411 => "0010001001000100001000",
			1412 => "0011100010011000000100",
			1413 => "1111111001011000101001",
			1414 => "0000001001011000101001",
			1415 => "0000000010100000000100",
			1416 => "1111111001011000101001",
			1417 => "0000001001011000101001",
			1418 => "0000010011110001100000",
			1419 => "0011011110011000111000",
			1420 => "0000010110010000100000",
			1421 => "0010110111011100011000",
			1422 => "0010101111011000001100",
			1423 => "0011100000110100001000",
			1424 => "0001000101010100000100",
			1425 => "0000000001011100010101",
			1426 => "0000000001011100010101",
			1427 => "0000000001011100010101",
			1428 => "0000101110011100001000",
			1429 => "0000000100110100000100",
			1430 => "0000000001011100010101",
			1431 => "0000000001011100010101",
			1432 => "0000000001011100010101",
			1433 => "0001000101011100000100",
			1434 => "0000000001011100010101",
			1435 => "0000000001011100010101",
			1436 => "0011100100111000010100",
			1437 => "0001011100010000001100",
			1438 => "0010110011010000001000",
			1439 => "0010010101011100000100",
			1440 => "0000000001011100010101",
			1441 => "0000000001011100010101",
			1442 => "0000000001011100010101",
			1443 => "0000000100010100000100",
			1444 => "0000000001011100010101",
			1445 => "0000000001011100010101",
			1446 => "0000000001011100010101",
			1447 => "0000010111100100010000",
			1448 => "0001100001100000001100",
			1449 => "0000001011001000001000",
			1450 => "0000000000011100000100",
			1451 => "0000000001011100010101",
			1452 => "0000000001011100010101",
			1453 => "0000000001011100010101",
			1454 => "0000000001011100010101",
			1455 => "0001001010000100001000",
			1456 => "0010000101101100000100",
			1457 => "0000000001011100010101",
			1458 => "0000000001011100010101",
			1459 => "0000011000011000000100",
			1460 => "0000000001011100010101",
			1461 => "0011100011101100001000",
			1462 => "0001111000101000000100",
			1463 => "0000000001011100010101",
			1464 => "0000000001011100010101",
			1465 => "0000000001011100010101",
			1466 => "0000101101011000010100",
			1467 => "0001000101010100001000",
			1468 => "0001000011010000000100",
			1469 => "0000000001011100010101",
			1470 => "0000000001011100010101",
			1471 => "0000110011001000001000",
			1472 => "0000111111011000000100",
			1473 => "0000000001011100010101",
			1474 => "0000000001011100010101",
			1475 => "0000000001011100010101",
			1476 => "0000000001011100010101",
			1477 => "0010110101011101010000",
			1478 => "0010101111011000001000",
			1479 => "0011100010010100000100",
			1480 => "0000000001011111011001",
			1481 => "0000000001011111011001",
			1482 => "0011101101100000100100",
			1483 => "0001011000000000001100",
			1484 => "0011011110011000001000",
			1485 => "0000110011000000000100",
			1486 => "0000000001011111011001",
			1487 => "0000000001011111011001",
			1488 => "0000000001011111011001",
			1489 => "0001000011000000001100",
			1490 => "0001011000101000001000",
			1491 => "0011111001111000000100",
			1492 => "0000000001011111011001",
			1493 => "0000000001011111011001",
			1494 => "0000000001011111011001",
			1495 => "0001011100101100000100",
			1496 => "0000000001011111011001",
			1497 => "0000011000011000000100",
			1498 => "0000000001011111011001",
			1499 => "0000000001011111011001",
			1500 => "0011001110011000001000",
			1501 => "0001100100001000000100",
			1502 => "0000000001011111011001",
			1503 => "0000000001011111011001",
			1504 => "0001110001010000001100",
			1505 => "0000111100010000000100",
			1506 => "0000000001011111011001",
			1507 => "0001010001010000000100",
			1508 => "0000000001011111011001",
			1509 => "0000000001011111011001",
			1510 => "0001011000000000001000",
			1511 => "0011100111100000000100",
			1512 => "0000000001011111011001",
			1513 => "0000000001011111011001",
			1514 => "0011111101001100000100",
			1515 => "0000000001011111011001",
			1516 => "0000000001011111011001",
			1517 => "0010010011001000010000",
			1518 => "0010101011000000001000",
			1519 => "0011111100111100000100",
			1520 => "0000000001011111011001",
			1521 => "0000000001011111011001",
			1522 => "0000011001100000000100",
			1523 => "0000000001011111011001",
			1524 => "0000000001011111011001",
			1525 => "0000000001011111011001",
			1526 => "0010100011000101010000",
			1527 => "0000011111011100111100",
			1528 => "0001011011000000110000",
			1529 => "0000111000000000011100",
			1530 => "0010110111011100010000",
			1531 => "0001101000110100001000",
			1532 => "0000001011010000000100",
			1533 => "0000000001100001111101",
			1534 => "1111111001100001111101",
			1535 => "0011011110011000000100",
			1536 => "0000000001100001111101",
			1537 => "0000001001100001111101",
			1538 => "0011011011101100000100",
			1539 => "0000001001100001111101",
			1540 => "0011010101011100000100",
			1541 => "1111111001100001111101",
			1542 => "0000000001100001111101",
			1543 => "0010010101101100000100",
			1544 => "1111111001100001111101",
			1545 => "0000000110111100001000",
			1546 => "0001111001010000000100",
			1547 => "0000001001100001111101",
			1548 => "0000000001100001111101",
			1549 => "0001110100101100000100",
			1550 => "1111111001100001111101",
			1551 => "0000000001100001111101",
			1552 => "0001011000100000001000",
			1553 => "0010001001000100000100",
			1554 => "0000001001100001111101",
			1555 => "0000000001100001111101",
			1556 => "1111111001100001111101",
			1557 => "0001010001011000001100",
			1558 => "0001011100000000001000",
			1559 => "0010101000000000000100",
			1560 => "1111111001100001111101",
			1561 => "0000000001100001111101",
			1562 => "1111111001100001111101",
			1563 => "0000111011111000000100",
			1564 => "0000000001100001111101",
			1565 => "0000000001100001111101",
			1566 => "1111111001100001111101",
			1567 => "0001100100110000111000",
			1568 => "0001111000111000011100",
			1569 => "0001111111011000000100",
			1570 => "0000000001100110000001",
			1571 => "0010101000111000010000",
			1572 => "0011001010100100000100",
			1573 => "0000000001100110000001",
			1574 => "0000011000011000000100",
			1575 => "0000000001100110000001",
			1576 => "0010001111001000000100",
			1577 => "0000000001100110000001",
			1578 => "0000000001100110000001",
			1579 => "0011001100101000000100",
			1580 => "0000000001100110000001",
			1581 => "0000000001100110000001",
			1582 => "0000111111011000001000",
			1583 => "0011100010011000000100",
			1584 => "0000000001100110000001",
			1585 => "0000000001100110000001",
			1586 => "0011100010110000001100",
			1587 => "0011001100101000000100",
			1588 => "0000000001100110000001",
			1589 => "0011001001001000000100",
			1590 => "0000000001100110000001",
			1591 => "0000000001100110000001",
			1592 => "0011100011101100000100",
			1593 => "0000000001100110000001",
			1594 => "0000000001100110000001",
			1595 => "0011110011111101000100",
			1596 => "0001011001010100011100",
			1597 => "0010010101011100001000",
			1598 => "0000000110111100000100",
			1599 => "0000000001100110000001",
			1600 => "0000000001100110000001",
			1601 => "0011111001111000001000",
			1602 => "0000100011011100000100",
			1603 => "0000000001100110000001",
			1604 => "0000000001100110000001",
			1605 => "0011110010101000001000",
			1606 => "0000001011001100000100",
			1607 => "0000000001100110000001",
			1608 => "0000000001100110000001",
			1609 => "0000000001100110000001",
			1610 => "0011000101011100010000",
			1611 => "0011010101010100001100",
			1612 => "0011000011010000001000",
			1613 => "0011110110011000000100",
			1614 => "0000000001100110000001",
			1615 => "0000000001100110000001",
			1616 => "0000000001100110000001",
			1617 => "0000000001100110000001",
			1618 => "0010101011000000001100",
			1619 => "0000000101101000000100",
			1620 => "0000000001100110000001",
			1621 => "0010110101101100000100",
			1622 => "0000000001100110000001",
			1623 => "0000000001100110000001",
			1624 => "0010111001000100000100",
			1625 => "0000000001100110000001",
			1626 => "0001001100010000000100",
			1627 => "0000000001100110000001",
			1628 => "0000000001100110000001",
			1629 => "0001001100000000000100",
			1630 => "0000000001100110000001",
			1631 => "0000000001100110000001",
			1632 => "0000110011001001000100",
			1633 => "0000010001110000010100",
			1634 => "0000011000111100000100",
			1635 => "0000000001101010010101",
			1636 => "0001000101101100001100",
			1637 => "0001010101111000001000",
			1638 => "0001011101101000000100",
			1639 => "0000000001101010010101",
			1640 => "0000000001101010010101",
			1641 => "0000000001101010010101",
			1642 => "0000000001101010010101",
			1643 => "0000010111100100010100",
			1644 => "0001000111011100001100",
			1645 => "0001001011101100001000",
			1646 => "0001111000000100000100",
			1647 => "0000000001101010010101",
			1648 => "0000000001101010010101",
			1649 => "0000000001101010010101",
			1650 => "0000000001110100000100",
			1651 => "0000000001101010010101",
			1652 => "0000001001101010010101",
			1653 => "0001100111101000011000",
			1654 => "0001111000111000001100",
			1655 => "0011000110001100000100",
			1656 => "0000000001101010010101",
			1657 => "0010010101101100000100",
			1658 => "0000000001101010010101",
			1659 => "0000000001101010010101",
			1660 => "0000110110000000001000",
			1661 => "0010101111111100000100",
			1662 => "0000000001101010010101",
			1663 => "0000000001101010010101",
			1664 => "0000000001101010010101",
			1665 => "0000000001101010010101",
			1666 => "0001011011000000101100",
			1667 => "0001101101010000011100",
			1668 => "0000101101011100011000",
			1669 => "0010101000101000001100",
			1670 => "0001101000110100001000",
			1671 => "0000001011001000000100",
			1672 => "0000000001101010010101",
			1673 => "1111111001101010010101",
			1674 => "0000000001101010010101",
			1675 => "0000011000011000000100",
			1676 => "0000000001101010010101",
			1677 => "0011100011101100000100",
			1678 => "0000000001101010010101",
			1679 => "0000000001101010010101",
			1680 => "1111111001101010010101",
			1681 => "0000111000000000000100",
			1682 => "0000000001101010010101",
			1683 => "0001001111011000001000",
			1684 => "0011001001000100000100",
			1685 => "0000000001101010010101",
			1686 => "0000000001101010010101",
			1687 => "0000000001101010010101",
			1688 => "0000000110010100000100",
			1689 => "0000000001101010010101",
			1690 => "0011000101010100000100",
			1691 => "0000000001101010010101",
			1692 => "0000101111001100001100",
			1693 => "0000111001010000000100",
			1694 => "0000000001101010010101",
			1695 => "0011011100101000000100",
			1696 => "0000001001101010010101",
			1697 => "0000000001101010010101",
			1698 => "0010101011000000000100",
			1699 => "0000000001101010010101",
			1700 => "0000000001101010010101",
			1701 => "0001111111011000000100",
			1702 => "1111111001101101000001",
			1703 => "0000110011000000001000",
			1704 => "0000000101011000000100",
			1705 => "0000000001101101000001",
			1706 => "0000001001101101000001",
			1707 => "0010110111011100011100",
			1708 => "0001011000101000010000",
			1709 => "0001111000111000000100",
			1710 => "0000000001101101000001",
			1711 => "0010101000000000000100",
			1712 => "1111111001101101000001",
			1713 => "0000010110010000000100",
			1714 => "0000000001101101000001",
			1715 => "0000000001101101000001",
			1716 => "0000111011111000000100",
			1717 => "1111111001101101000001",
			1718 => "0000010111100100000100",
			1719 => "0000000001101101000001",
			1720 => "0000000001101101000001",
			1721 => "0010101011111000011000",
			1722 => "0001111000101000001000",
			1723 => "0001101010110100000100",
			1724 => "0000000001101101000001",
			1725 => "0000001001101101000001",
			1726 => "0000000101101000001000",
			1727 => "0001011000111000000100",
			1728 => "0000000001101101000001",
			1729 => "1111111001101101000001",
			1730 => "0001011000101000000100",
			1731 => "0000000001101101000001",
			1732 => "0000001001101101000001",
			1733 => "0011001001000100001100",
			1734 => "0010000101011100001000",
			1735 => "0000010111110000000100",
			1736 => "0000000001101101000001",
			1737 => "0000000001101101000001",
			1738 => "1111111001101101000001",
			1739 => "0000001110101000000100",
			1740 => "0000000001101101000001",
			1741 => "0000010101010100000100",
			1742 => "0000000001101101000001",
			1743 => "0000000001101101000001",
			1744 => "0001001001010001101000",
			1745 => "0001010011001000100000",
			1746 => "0001011111011000011100",
			1747 => "0001101010001000010000",
			1748 => "0010111011101100001100",
			1749 => "0010110110110100000100",
			1750 => "1111111001110000010111",
			1751 => "0000010110010000000100",
			1752 => "0000000001110000010111",
			1753 => "0000001001110000010111",
			1754 => "1111111001110000010111",
			1755 => "0011100110110000001000",
			1756 => "0000010001110000000100",
			1757 => "0000000001110000010111",
			1758 => "0000001001110000010111",
			1759 => "1111111001110000010111",
			1760 => "1111111001110000010111",
			1761 => "0000110011001000011000",
			1762 => "0001000111011100000100",
			1763 => "1111111001110000010111",
			1764 => "0001000110000000001100",
			1765 => "0001000101101100001000",
			1766 => "0000110101111000000100",
			1767 => "0000000001110000010111",
			1768 => "0000001001110000010111",
			1769 => "0000001001110000010111",
			1770 => "0010001001000100000100",
			1771 => "0000000001110000010111",
			1772 => "1111111001110000010111",
			1773 => "0010001111001000011100",
			1774 => "0010110111011100010000",
			1775 => "0000010110010000001000",
			1776 => "0001111000000100000100",
			1777 => "0000001001110000010111",
			1778 => "1111111001110000010111",
			1779 => "0001111001010000000100",
			1780 => "0000000001110000010111",
			1781 => "0000000001110000010111",
			1782 => "0001011001010000000100",
			1783 => "0000000001110000010111",
			1784 => "0010101011111000000100",
			1785 => "0000001001110000010111",
			1786 => "0000000001110000010111",
			1787 => "0001001100000000001000",
			1788 => "0011100101110000000100",
			1789 => "0000000001110000010111",
			1790 => "1111111001110000010111",
			1791 => "0010010011001000001000",
			1792 => "0011001100101000000100",
			1793 => "0000000001110000010111",
			1794 => "0000001001110000010111",
			1795 => "0000000001110000010111",
			1796 => "1111111001110000010111",
			1797 => "0000101011001000011000",
			1798 => "0011001010100100001000",
			1799 => "0011111000101100000100",
			1800 => "1111111001110010000001",
			1801 => "0000001001110010000001",
			1802 => "0001111000000000001000",
			1803 => "0011110101001000000100",
			1804 => "1111111001110010000001",
			1805 => "0000001001110010000001",
			1806 => "0011110100000100000100",
			1807 => "1111111001110010000001",
			1808 => "1111111001110010000001",
			1809 => "0000010110001100011100",
			1810 => "0001001100110000011000",
			1811 => "0011001100101000010100",
			1812 => "0001100000000100010000",
			1813 => "0001000101111000001000",
			1814 => "0001001010000100000100",
			1815 => "0000001001110010000001",
			1816 => "0000010001110010000001",
			1817 => "0010000101101100000100",
			1818 => "0000001001110010000001",
			1819 => "1111111001110010000001",
			1820 => "1111111001110010000001",
			1821 => "0000001001110010000001",
			1822 => "1111111001110010000001",
			1823 => "1111111001110010000001",
			1824 => "0011110100001100001100",
			1825 => "0011111110000000000100",
			1826 => "1111111001110011110101",
			1827 => "0000100111101000000100",
			1828 => "0000001001110011110101",
			1829 => "1111111001110011110101",
			1830 => "0000011101000000100100",
			1831 => "0000111101101000001000",
			1832 => "0000000101011000000100",
			1833 => "0000000001110011110101",
			1834 => "0000001001110011110101",
			1835 => "0011100101001000000100",
			1836 => "0000010001110011110101",
			1837 => "0000000010100100001100",
			1838 => "0011100011010100001000",
			1839 => "0010011001000100000100",
			1840 => "0000001001110011110101",
			1841 => "1111111001110011110101",
			1842 => "1111111001110011110101",
			1843 => "0011100101110100000100",
			1844 => "1111111001110011110101",
			1845 => "0000101011010000000100",
			1846 => "0000001001110011110101",
			1847 => "0000000001110011110101",
			1848 => "0011110011100000001000",
			1849 => "0001000110000000000100",
			1850 => "0000000001110011110101",
			1851 => "1111111001110011110101",
			1852 => "0000001001110011110101",
			1853 => "0011110001100000010000",
			1854 => "0010010110000000001100",
			1855 => "0001100000100000000100",
			1856 => "1111111001110101111001",
			1857 => "0001111000000000000100",
			1858 => "0000011001110101111001",
			1859 => "1111111001110101111001",
			1860 => "1111111001110101111001",
			1861 => "0000011101000000101100",
			1862 => "0010110111011100100000",
			1863 => "0010101000111000001100",
			1864 => "0011100010011000000100",
			1865 => "0000001001110101111001",
			1866 => "0011010110001100000100",
			1867 => "0000001001110101111001",
			1868 => "0000010001110101111001",
			1869 => "0011100011011000001000",
			1870 => "0000101011010000000100",
			1871 => "0000010001110101111001",
			1872 => "1111111001110101111001",
			1873 => "0000010001100100001000",
			1874 => "0010110011010000000100",
			1875 => "1111111001110101111001",
			1876 => "0000000001110101111001",
			1877 => "0000001001110101111001",
			1878 => "0000101011100100001000",
			1879 => "0011101101100000000100",
			1880 => "0000010001110101111001",
			1881 => "1111111001110101111001",
			1882 => "0000011001110101111001",
			1883 => "0001000110000000000100",
			1884 => "0000000001110101111001",
			1885 => "1111111001110101111001",
			1886 => "0010101000111000101000",
			1887 => "0001001100101000011000",
			1888 => "0011001010100100001100",
			1889 => "0001111000000100000100",
			1890 => "0000000001111000111101",
			1891 => "0000000101011000000100",
			1892 => "0000000001111000111101",
			1893 => "0000000001111000111101",
			1894 => "0000110011000000001000",
			1895 => "0001010110000000000100",
			1896 => "0000000001111000111101",
			1897 => "0000000001111000111101",
			1898 => "0000000001111000111101",
			1899 => "0001000110000000001000",
			1900 => "0001111111011000000100",
			1901 => "0000000001111000111101",
			1902 => "0000000001111000111101",
			1903 => "0000110011000000000100",
			1904 => "0000000001111000111101",
			1905 => "0000000001111000111101",
			1906 => "0010110111011100010100",
			1907 => "0000101011010000010000",
			1908 => "0000001100001000001100",
			1909 => "0001011001010100000100",
			1910 => "0000000001111000111101",
			1911 => "0001011000101000000100",
			1912 => "0000000001111000111101",
			1913 => "0000000001111000111101",
			1914 => "0000000001111000111101",
			1915 => "0000000001111000111101",
			1916 => "0010101011111000010100",
			1917 => "0001011001010000001100",
			1918 => "0011100111001000001000",
			1919 => "0010101101001000000100",
			1920 => "0000000001111000111101",
			1921 => "0000000001111000111101",
			1922 => "0000000001111000111101",
			1923 => "0000011111011100000100",
			1924 => "0000000001111000111101",
			1925 => "0000000001111000111101",
			1926 => "0011001001000100001100",
			1927 => "0010000101011100001000",
			1928 => "0000010111110000000100",
			1929 => "0000000001111000111101",
			1930 => "0000000001111000111101",
			1931 => "0000000001111000111101",
			1932 => "0010011000000100000100",
			1933 => "0000000001111000111101",
			1934 => "0000000001111000111101",
			1935 => "0011110111100000010100",
			1936 => "0010010110000000010000",
			1937 => "0010001001000100000100",
			1938 => "1111111001111011000001",
			1939 => "0000010011110000001000",
			1940 => "0001011001001000000100",
			1941 => "1111111001111011000001",
			1942 => "0000001001111011000001",
			1943 => "1111111001111011000001",
			1944 => "1111111001111011000001",
			1945 => "0000011101000000100100",
			1946 => "0001101110100000000100",
			1947 => "0000001001111011000001",
			1948 => "0011010111011100010100",
			1949 => "0000111101101000000100",
			1950 => "0000001001111011000001",
			1951 => "0001011100110000001000",
			1952 => "0011001010100100000100",
			1953 => "0000000001111011000001",
			1954 => "1111111001111011000001",
			1955 => "0001111101001000000100",
			1956 => "1111111001111011000001",
			1957 => "0000001001111011000001",
			1958 => "0000001111001100001000",
			1959 => "0011100011101100000100",
			1960 => "0000001001111011000001",
			1961 => "1111111001111011000001",
			1962 => "0000001001111011000001",
			1963 => "0011010101011100001000",
			1964 => "0010110101011100000100",
			1965 => "1111111001111011000001",
			1966 => "0000001001111011000001",
			1967 => "1111111001111011000001",
			1968 => "0011011110011000100000",
			1969 => "0000001011010000011000",
			1970 => "0010001111111100001100",
			1971 => "0011110111100000000100",
			1972 => "0000000001111101101101",
			1973 => "0001111001010100000100",
			1974 => "0000000001111101101101",
			1975 => "0000000001111101101101",
			1976 => "0001110011001000000100",
			1977 => "0000000001111101101101",
			1978 => "0010100011000000000100",
			1979 => "0000000001111101101101",
			1980 => "0000000001111101101101",
			1981 => "0001110001010000000100",
			1982 => "0000000001111101101101",
			1983 => "0000000001111101101101",
			1984 => "0000101111101100100000",
			1985 => "0010011001001000001000",
			1986 => "0001001100101000000100",
			1987 => "0000000001111101101101",
			1988 => "0000000001111101101101",
			1989 => "0000111100010000000100",
			1990 => "0000000001111101101101",
			1991 => "0001000011000000001000",
			1992 => "0000001101110100000100",
			1993 => "0000000001111101101101",
			1994 => "0000000001111101101101",
			1995 => "0000001000010000000100",
			1996 => "0000000001111101101101",
			1997 => "0000000100010100000100",
			1998 => "0000000001111101101101",
			1999 => "0000000001111101101101",
			2000 => "0000011001100000000100",
			2001 => "0000000001111101101101",
			2002 => "0001001100000000001000",
			2003 => "0001011101001000000100",
			2004 => "0000000001111101101101",
			2005 => "0000000001111101101101",
			2006 => "0000001110101000000100",
			2007 => "0000000001111101101101",
			2008 => "0001111100011100000100",
			2009 => "0000000001111101101101",
			2010 => "0000000001111101101101",
			2011 => "0000011111011100101100",
			2012 => "0001111111011000000100",
			2013 => "1111111001111111101001",
			2014 => "0010101111011000001000",
			2015 => "0000000101011000000100",
			2016 => "1111111001111111101001",
			2017 => "0000001001111111101001",
			2018 => "0010100011001000000100",
			2019 => "1111111001111111101001",
			2020 => "0000100011111000010000",
			2021 => "0001111000000100001000",
			2022 => "0000000101000000000100",
			2023 => "0000000001111111101001",
			2024 => "0000001001111111101001",
			2025 => "0011100100001100000100",
			2026 => "0000000001111111101001",
			2027 => "1111111001111111101001",
			2028 => "0010010101011100000100",
			2029 => "1111111001111111101001",
			2030 => "0000101010010100000100",
			2031 => "0000000001111111101001",
			2032 => "0000000001111111101001",
			2033 => "0001011100000000001100",
			2034 => "0001110100101100000100",
			2035 => "0000000001111111101001",
			2036 => "0011001000000100000100",
			2037 => "0000000001111111101001",
			2038 => "0000000001111111101001",
			2039 => "0011110011100000000100",
			2040 => "1111111001111111101001",
			2041 => "0000000001111111101001",
			2042 => "0000000110001000001100",
			2043 => "0000111000101000000100",
			2044 => "1111111010000001110101",
			2045 => "0001001100000000000100",
			2046 => "0000001010000001110101",
			2047 => "1111111010000001110101",
			2048 => "0001000111011100001100",
			2049 => "0011101100011000000100",
			2050 => "0000000010000001110101",
			2051 => "0001010101111000000100",
			2052 => "0000000010000001110101",
			2053 => "1111111010000001110101",
			2054 => "0000110011001000001100",
			2055 => "0011010110001100000100",
			2056 => "0000000010000001110101",
			2057 => "0000000000000000000100",
			2058 => "0000000010000001110101",
			2059 => "0000001010000001110101",
			2060 => "0010001111001000011000",
			2061 => "0001001001000100001000",
			2062 => "0011110100111100000100",
			2063 => "1111111010000001110101",
			2064 => "0000000010000001110101",
			2065 => "0011011011101100001000",
			2066 => "0010111011101100000100",
			2067 => "0000001010000001110101",
			2068 => "1111111010000001110101",
			2069 => "0011011010100100000100",
			2070 => "0000001010000001110101",
			2071 => "0000000010000001110101",
			2072 => "0001001100000000000100",
			2073 => "1111111010000001110101",
			2074 => "0010010011001000000100",
			2075 => "0000000010000001110101",
			2076 => "1111111010000001110101",
			2077 => "0011000101010100111100",
			2078 => "0010101000111000010100",
			2079 => "0000110011001000010000",
			2080 => "0001111111011000000100",
			2081 => "0000000010000100101001",
			2082 => "0000000001110100001000",
			2083 => "0011101101000100000100",
			2084 => "0000000010000100101001",
			2085 => "0000000010000100101001",
			2086 => "0000000010000100101001",
			2087 => "0000000010000100101001",
			2088 => "0000010001100100011100",
			2089 => "0000101100010100001100",
			2090 => "0011101001011100000100",
			2091 => "0000000010000100101001",
			2092 => "0011101101100000000100",
			2093 => "0000000010000100101001",
			2094 => "0000000010000100101001",
			2095 => "0000011001100100000100",
			2096 => "0000000010000100101001",
			2097 => "0001011000000100001000",
			2098 => "0001011111011000000100",
			2099 => "0000000010000100101001",
			2100 => "0000000010000100101001",
			2101 => "0000000010000100101001",
			2102 => "0000011101000000001000",
			2103 => "0011100100111000000100",
			2104 => "0000000010000100101001",
			2105 => "0000000010000100101001",
			2106 => "0000000010000100101001",
			2107 => "0001011100010000001100",
			2108 => "0001011100000000001000",
			2109 => "0001010011000000000100",
			2110 => "0000000010000100101001",
			2111 => "0000000010000100101001",
			2112 => "0000000010000100101001",
			2113 => "0001011100011100010000",
			2114 => "0000010110110100001100",
			2115 => "0010101111101000001000",
			2116 => "0010110101011100000100",
			2117 => "0000000010000100101001",
			2118 => "0000000010000100101001",
			2119 => "0000000010000100101001",
			2120 => "0000000010000100101001",
			2121 => "0000000010000100101001",
			2122 => "0011110000100101001000",
			2123 => "0000110011001000100000",
			2124 => "0001010011001000010000",
			2125 => "0010100011000000001000",
			2126 => "0011111000101100000100",
			2127 => "0000000010000111110101",
			2128 => "0000000010000111110101",
			2129 => "0000110110000000000100",
			2130 => "0000000010000111110101",
			2131 => "0000000010000111110101",
			2132 => "0000010111100100001000",
			2133 => "0000000001110100000100",
			2134 => "0000000010000111110101",
			2135 => "0000000010000111110101",
			2136 => "0001001001000100000100",
			2137 => "0000000010000111110101",
			2138 => "0000000010000111110101",
			2139 => "0000000101101000100000",
			2140 => "0000011000011000001100",
			2141 => "0000001011001000001000",
			2142 => "0011110111100000000100",
			2143 => "0000000010000111110101",
			2144 => "0000000010000111110101",
			2145 => "0000000010000111110101",
			2146 => "0001111000101000010000",
			2147 => "0000010011110000001000",
			2148 => "0010001010000100000100",
			2149 => "0000000010000111110101",
			2150 => "0000000010000111110101",
			2151 => "0001011001010000000100",
			2152 => "0000000010000111110101",
			2153 => "0000000010000111110101",
			2154 => "0000000010000111110101",
			2155 => "0000101101110000000100",
			2156 => "0000000010000111110101",
			2157 => "0000000010000111110101",
			2158 => "0011111011011000010100",
			2159 => "0011100110000100001100",
			2160 => "0010000011001000001000",
			2161 => "0001101101010000000100",
			2162 => "0000000010000111110101",
			2163 => "0000000010000111110101",
			2164 => "0000000010000111110101",
			2165 => "0000111101001000000100",
			2166 => "0000000010000111110101",
			2167 => "0000000010000111110101",
			2168 => "0001111100101100000100",
			2169 => "0000000010000111110101",
			2170 => "0000000010100000000100",
			2171 => "0000000010000111110101",
			2172 => "0000000010000111110101",
			2173 => "0011111000101100010000",
			2174 => "0010010110000000001100",
			2175 => "0010001001000100000100",
			2176 => "1111111010001001111001",
			2177 => "0011000011010000000100",
			2178 => "1111111010001001111001",
			2179 => "0000001010001001111001",
			2180 => "1111111010001001111001",
			2181 => "0000010110001100110000",
			2182 => "0010101101001000010100",
			2183 => "0000000101011000000100",
			2184 => "1111111010001001111001",
			2185 => "0011100110111000001100",
			2186 => "0011010110110100000100",
			2187 => "0000000010001001111001",
			2188 => "0000001011100100000100",
			2189 => "0000001010001001111001",
			2190 => "0000010010001001111001",
			2191 => "1111111010001001111001",
			2192 => "0010110011010000001100",
			2193 => "0000011000011000000100",
			2194 => "1111111010001001111001",
			2195 => "0010000101101100000100",
			2196 => "0000011010001001111001",
			2197 => "1111111010001001111001",
			2198 => "0001111000101000000100",
			2199 => "0000010010001001111001",
			2200 => "0000101011100100000100",
			2201 => "1111111010001001111001",
			2202 => "0011001100101000000100",
			2203 => "0000000010001001111001",
			2204 => "0000010010001001111001",
			2205 => "1111111010001001111001",
			2206 => "0011111000101100010000",
			2207 => "0010010110000000001100",
			2208 => "0010001001000100000100",
			2209 => "1111111010001011101101",
			2210 => "0001011000111000000100",
			2211 => "1111111010001011101101",
			2212 => "0000001010001011101101",
			2213 => "1111111010001011101101",
			2214 => "0000010110001100101000",
			2215 => "0010101111011000000100",
			2216 => "0000001010001011101101",
			2217 => "0010010101011100001000",
			2218 => "0001010011000000000100",
			2219 => "0000000010001011101101",
			2220 => "1111111010001011101101",
			2221 => "0000000010100100001100",
			2222 => "0001111001010100000100",
			2223 => "0000001010001011101101",
			2224 => "0000110011100100000100",
			2225 => "1111111010001011101101",
			2226 => "1111111010001011101101",
			2227 => "0000111000000000001000",
			2228 => "0001000101010100000100",
			2229 => "0000000010001011101101",
			2230 => "0000001010001011101101",
			2231 => "0000100110010100000100",
			2232 => "0000001010001011101101",
			2233 => "0000000010001011101101",
			2234 => "1111111010001011101101",
			2235 => "0000000110001000001100",
			2236 => "0000111000101000000100",
			2237 => "1111111010001110010001",
			2238 => "0001001100000000000100",
			2239 => "0000001010001110010001",
			2240 => "1111111010001110010001",
			2241 => "0001011000000000011000",
			2242 => "0001011111011000001100",
			2243 => "0011100110110000001000",
			2244 => "0001100100110000000100",
			2245 => "0000000010001110010001",
			2246 => "0000001010001110010001",
			2247 => "1111111010001110010001",
			2248 => "0001110001010000001000",
			2249 => "0011001010100100000100",
			2250 => "0000000010001110010001",
			2251 => "1111111010001110010001",
			2252 => "0000001010001110010001",
			2253 => "0010001001000100011100",
			2254 => "0010011101101000010100",
			2255 => "0011110110011000001100",
			2256 => "0001010011000100001000",
			2257 => "0000101101011100000100",
			2258 => "0000001010001110010001",
			2259 => "0000000010001110010001",
			2260 => "1111111010001110010001",
			2261 => "0001101110101100000100",
			2262 => "1111111010001110010001",
			2263 => "0000000010001110010001",
			2264 => "0011110001100000000100",
			2265 => "0000000010001110010001",
			2266 => "0000001010001110010001",
			2267 => "0001111000101000000100",
			2268 => "0000000010001110010001",
			2269 => "0011110011100000001100",
			2270 => "0011001001000100000100",
			2271 => "1111111010001110010001",
			2272 => "0011011100101000000100",
			2273 => "0000001010001110010001",
			2274 => "1111111010001110010001",
			2275 => "0000001010001110010001",
			2276 => "0011110100011001000000",
			2277 => "0001111100110000011100",
			2278 => "0000001001110100010100",
			2279 => "0011110111100000010000",
			2280 => "0010001001000100000100",
			2281 => "0000000010010001100101",
			2282 => "0010001010000100001000",
			2283 => "0000011000011000000100",
			2284 => "0000000010010001100101",
			2285 => "0000000010010001100101",
			2286 => "0000000010010001100101",
			2287 => "0000000010010001100101",
			2288 => "0011100011010100000100",
			2289 => "0000000010010001100101",
			2290 => "0000000010010001100101",
			2291 => "0001001010000100001100",
			2292 => "0000110110000000001000",
			2293 => "0000110101101100000100",
			2294 => "0000000010010001100101",
			2295 => "0000000010010001100101",
			2296 => "1111111010010001100101",
			2297 => "0000101010101000001100",
			2298 => "0001110110101100001000",
			2299 => "0000010111110000000100",
			2300 => "0000000010010001100101",
			2301 => "0000000010010001100101",
			2302 => "0000000010010001100101",
			2303 => "0000100010101100000100",
			2304 => "0000000010010001100101",
			2305 => "0001001000111000000100",
			2306 => "0000000010010001100101",
			2307 => "0000000010010001100101",
			2308 => "0011111001111000001100",
			2309 => "0001000011000000001000",
			2310 => "0010011100101000000100",
			2311 => "0000000010010001100101",
			2312 => "0000000010010001100101",
			2313 => "0000000010010001100101",
			2314 => "0010011101101000010000",
			2315 => "0000111000000000001100",
			2316 => "0001101000010100000100",
			2317 => "0000000010010001100101",
			2318 => "0011110011111100000100",
			2319 => "0000000010010001100101",
			2320 => "0000000010010001100101",
			2321 => "0000000010010001100101",
			2322 => "0000011101000000000100",
			2323 => "0000000010010001100101",
			2324 => "0000001101111000000100",
			2325 => "0000000010010001100101",
			2326 => "0000101101011000000100",
			2327 => "0000000010010001100101",
			2328 => "0000000010010001100101",
			2329 => "0011111000101100001100",
			2330 => "0001111000000000001000",
			2331 => "0001100000100000000100",
			2332 => "1111111010010011100001",
			2333 => "0000001010010011100001",
			2334 => "1111111010010011100001",
			2335 => "0010000011001000110000",
			2336 => "0011010110001100001100",
			2337 => "0010101111011000000100",
			2338 => "0000001010010011100001",
			2339 => "0001001010100100000100",
			2340 => "0000000010010011100001",
			2341 => "1111111010010011100001",
			2342 => "0011100111001000010000",
			2343 => "0011111100111100001100",
			2344 => "0001111000101000001000",
			2345 => "0001011100110000000100",
			2346 => "0000000010010011100001",
			2347 => "0000001010010011100001",
			2348 => "1111111010010011100001",
			2349 => "0000001010010011100001",
			2350 => "0011000101101100010000",
			2351 => "0010001111001000001000",
			2352 => "0001000111011100000100",
			2353 => "1111111010010011100001",
			2354 => "0000000010010011100001",
			2355 => "0001011100010000000100",
			2356 => "0000000010010011100001",
			2357 => "1111111010010011100001",
			2358 => "0000001010010011100001",
			2359 => "1111111010010011100001",
			2360 => "0001001100101000100100",
			2361 => "0000110011000000011000",
			2362 => "0001111000000100000100",
			2363 => "0000000010010110101101",
			2364 => "0010000101101100001000",
			2365 => "0000000101011000000100",
			2366 => "0000000010010110101101",
			2367 => "0000001010010110101101",
			2368 => "0000110101101100001000",
			2369 => "0000111100101000000100",
			2370 => "0000000010010110101101",
			2371 => "0000000010010110101101",
			2372 => "0000000010010110101101",
			2373 => "0011001010100100001000",
			2374 => "0010010101011100000100",
			2375 => "0000000010010110101101",
			2376 => "0000000010010110101101",
			2377 => "1111111010010110101101",
			2378 => "0010101000111000010100",
			2379 => "0011100010011000010000",
			2380 => "0001111000000000001000",
			2381 => "0011010110001100000100",
			2382 => "0000000010010110101101",
			2383 => "0000000010010110101101",
			2384 => "0001011001000100000100",
			2385 => "0000000010010110101101",
			2386 => "0000000010010110101101",
			2387 => "0000001010010110101101",
			2388 => "0001011100110000001100",
			2389 => "0001101101010000001000",
			2390 => "0010101100010000000100",
			2391 => "0000000010010110101101",
			2392 => "1111111010010110101101",
			2393 => "0000000010010110101101",
			2394 => "0010101011000000010100",
			2395 => "0011011110011000001000",
			2396 => "0000010111100100000100",
			2397 => "1111111010010110101101",
			2398 => "0000000010010110101101",
			2399 => "0000010111100100000100",
			2400 => "0000001010010110101101",
			2401 => "0001111000101000000100",
			2402 => "0000000010010110101101",
			2403 => "0000000010010110101101",
			2404 => "0010000101011100001000",
			2405 => "0000010111110000000100",
			2406 => "0000000010010110101101",
			2407 => "0000000010010110101101",
			2408 => "0011110011100000000100",
			2409 => "1111111010010110101101",
			2410 => "0000000010010110101101",
			2411 => "0001011100110000111100",
			2412 => "0010101000111000101000",
			2413 => "0011111011011100100000",
			2414 => "0011001010100100001100",
			2415 => "0001110011001000000100",
			2416 => "0000000010011010010001",
			2417 => "0001111000111000000100",
			2418 => "0000000010011010010001",
			2419 => "0000000010011010010001",
			2420 => "0001110011001000001000",
			2421 => "0000000101000000000100",
			2422 => "0000000010011010010001",
			2423 => "0000000010011010010001",
			2424 => "0010100101101100001000",
			2425 => "0000111100101000000100",
			2426 => "0000000010011010010001",
			2427 => "0000000010011010010001",
			2428 => "0000000010011010010001",
			2429 => "0001000111011100000100",
			2430 => "0000000010011010010001",
			2431 => "0000000010011010010001",
			2432 => "0000010001100100001100",
			2433 => "0001010101111000001000",
			2434 => "0010111010100100000100",
			2435 => "0000000010011010010001",
			2436 => "0000000010011010010001",
			2437 => "0000000010011010010001",
			2438 => "0000011101000000000100",
			2439 => "0000000010011010010001",
			2440 => "0000000010011010010001",
			2441 => "0010101011111000100100",
			2442 => "0010110011010000010000",
			2443 => "0000011000011000001000",
			2444 => "0000001011001000000100",
			2445 => "0000000010011010010001",
			2446 => "0000000010011010010001",
			2447 => "0010101001010100000100",
			2448 => "0000000010011010010001",
			2449 => "0000000010011010010001",
			2450 => "0000010111100100000100",
			2451 => "0000000010011010010001",
			2452 => "0010110111011100000100",
			2453 => "0000000010011010010001",
			2454 => "0001111000101000000100",
			2455 => "0000000010011010010001",
			2456 => "0011100110111000000100",
			2457 => "0000000010011010010001",
			2458 => "0000000010011010010001",
			2459 => "0011001001000100001100",
			2460 => "0001001001010100000100",
			2461 => "0000000010011010010001",
			2462 => "0001001111101000000100",
			2463 => "0000000010011010010001",
			2464 => "0000000010011010010001",
			2465 => "0010011000000100000100",
			2466 => "0000000010011010010001",
			2467 => "0000000010011010010001",
			2468 => "0011111010110000110000",
			2469 => "0011100001101100100000",
			2470 => "0000001001110100011100",
			2471 => "0011100000110100010100",
			2472 => "0011001010100100001000",
			2473 => "0000000100111100000100",
			2474 => "0000000010011101100101",
			2475 => "0000000010011101100101",
			2476 => "0000001011001000001000",
			2477 => "0000001011100000000100",
			2478 => "0000000010011101100101",
			2479 => "0000000010011101100101",
			2480 => "0000000010011101100101",
			2481 => "0000100011011100000100",
			2482 => "0000000010011101100101",
			2483 => "0000001010011101100101",
			2484 => "0000000010011101100101",
			2485 => "0000010001100100001000",
			2486 => "0001000101010100000100",
			2487 => "0000000010011101100101",
			2488 => "1111111010011101100101",
			2489 => "0000100011111000000100",
			2490 => "0000000010011101100101",
			2491 => "0000000010011101100101",
			2492 => "0011011110011000011000",
			2493 => "0000000100010100001100",
			2494 => "0011110111010000000100",
			2495 => "0000000010011101100101",
			2496 => "0001111001010000000100",
			2497 => "0000001010011101100101",
			2498 => "0000000010011101100101",
			2499 => "0011110101000100000100",
			2500 => "1111111010011101100101",
			2501 => "0011111110011100000100",
			2502 => "0000000010011101100101",
			2503 => "0000000010011101100101",
			2504 => "0000011001100000001100",
			2505 => "0001001001000100000100",
			2506 => "0000000010011101100101",
			2507 => "0000010111100100000100",
			2508 => "0000001010011101100101",
			2509 => "0000000010011101100101",
			2510 => "0000110011100100000100",
			2511 => "0000000010011101100101",
			2512 => "0001111001011000000100",
			2513 => "1111111010011101100101",
			2514 => "0001001100000000001000",
			2515 => "0001110001001000000100",
			2516 => "0000000010011101100101",
			2517 => "0000000010011101100101",
			2518 => "0010111001001000000100",
			2519 => "0000000010011101100101",
			2520 => "0000000010011101100101",
			2521 => "0011100000110100011000",
			2522 => "0000010110010000000100",
			2523 => "0000000010100000001001",
			2524 => "0011100010010100001100",
			2525 => "0011101101101100001000",
			2526 => "0000001010111100000100",
			2527 => "0000000010100000001001",
			2528 => "0000000010100000001001",
			2529 => "0000000010100000001001",
			2530 => "0011101111000100000100",
			2531 => "0000000010100000001001",
			2532 => "0000000010100000001001",
			2533 => "0001101110000100110000",
			2534 => "0001011111011000001000",
			2535 => "0000001101110100000100",
			2536 => "0000000010100000001001",
			2537 => "0000000010100000001001",
			2538 => "0001000101010100001000",
			2539 => "0001100101001100000100",
			2540 => "0000000010100000001001",
			2541 => "0000000010100000001001",
			2542 => "0000011001100000010000",
			2543 => "0000010001110000001000",
			2544 => "0001011100101100000100",
			2545 => "0000000010100000001001",
			2546 => "0000000010100000001001",
			2547 => "0001100100110000000100",
			2548 => "0000000010100000001001",
			2549 => "0000000010100000001001",
			2550 => "0000100100010100001000",
			2551 => "0010110011010000000100",
			2552 => "0000000010100000001001",
			2553 => "0000000010100000001001",
			2554 => "0011000110000000000100",
			2555 => "0000000010100000001001",
			2556 => "0000000010100000001001",
			2557 => "0001111100101100000100",
			2558 => "0000000010100000001001",
			2559 => "0000000010100000000100",
			2560 => "0000000010100000001001",
			2561 => "0000000010100000001001",
			2562 => "0010001111111100101000",
			2563 => "0001100010110100001100",
			2564 => "0011001010100100001000",
			2565 => "0001010011001000000100",
			2566 => "0000000010100011101101",
			2567 => "0000000010100011101101",
			2568 => "0000000010100011101101",
			2569 => "0011100110110000010100",
			2570 => "0000100000000000010000",
			2571 => "0010000011010000000100",
			2572 => "0000000010100011101101",
			2573 => "0010101101001000000100",
			2574 => "0000000010100011101101",
			2575 => "0010011100101000000100",
			2576 => "0000000010100011101101",
			2577 => "0000000010100011101101",
			2578 => "0000000010100011101101",
			2579 => "0011100011101000000100",
			2580 => "0000000010100011101101",
			2581 => "0000000010100011101101",
			2582 => "0001011001010000101100",
			2583 => "0011010101010100011100",
			2584 => "0000110101111000010000",
			2585 => "0001011000000100001100",
			2586 => "0010101111011000001000",
			2587 => "0001010101101100000100",
			2588 => "0000000010100011101101",
			2589 => "0000000010100011101101",
			2590 => "0000000010100011101101",
			2591 => "0000000010100011101101",
			2592 => "0011101111000100001000",
			2593 => "0001110011001000000100",
			2594 => "0000000010100011101101",
			2595 => "0000000010100011101101",
			2596 => "0000000010100011101101",
			2597 => "0001111001010000001000",
			2598 => "0001111101001000000100",
			2599 => "0000000010100011101101",
			2600 => "0000000010100011101101",
			2601 => "0001011000000000000100",
			2602 => "0000000010100011101101",
			2603 => "0000000010100011101101",
			2604 => "0011011010100100001100",
			2605 => "0001111101001000000100",
			2606 => "0000000010100011101101",
			2607 => "0010101001011000000100",
			2608 => "0000000010100011101101",
			2609 => "0000000010100011101101",
			2610 => "0010111100101000001100",
			2611 => "0001111001010000001000",
			2612 => "0011111110000000000100",
			2613 => "0000000010100011101101",
			2614 => "0000000010100011101101",
			2615 => "0000000010100011101101",
			2616 => "0010010011001000000100",
			2617 => "0000000010100011101101",
			2618 => "0000000010100011101101",
			2619 => "0010101000111000101000",
			2620 => "0011111011011100100000",
			2621 => "0001111000111000010100",
			2622 => "0001111111011000000100",
			2623 => "0000000010100111001001",
			2624 => "0011001010100100000100",
			2625 => "0000000010100111001001",
			2626 => "0000011000011000000100",
			2627 => "0000000010100111001001",
			2628 => "0010001111001000000100",
			2629 => "0000000010100111001001",
			2630 => "0000000010100111001001",
			2631 => "0000110110000000001000",
			2632 => "0001010101101100000100",
			2633 => "0000000010100111001001",
			2634 => "0000000010100111001001",
			2635 => "0000000010100111001001",
			2636 => "0001000101010100000100",
			2637 => "0000000010100111001001",
			2638 => "0000000010100111001001",
			2639 => "0010110111011100100000",
			2640 => "0000010001100100011000",
			2641 => "0001011000000100001000",
			2642 => "0011010110001100000100",
			2643 => "0000000010100111001001",
			2644 => "0000000010100111001001",
			2645 => "0000111011111000001000",
			2646 => "0000011000111100000100",
			2647 => "0000000010100111001001",
			2648 => "1111111010100111001001",
			2649 => "0010101001011000000100",
			2650 => "0000000010100111001001",
			2651 => "0000000010100111001001",
			2652 => "0010010101101100000100",
			2653 => "0000000010100111001001",
			2654 => "0000000010100111001001",
			2655 => "0000000101101000011000",
			2656 => "0001111000101000001100",
			2657 => "0001011011000000001000",
			2658 => "0010011010000100000100",
			2659 => "0000000010100111001001",
			2660 => "0000000010100111001001",
			2661 => "0000000010100111001001",
			2662 => "0001011110111000000100",
			2663 => "0000000010100111001001",
			2664 => "0001001101001000000100",
			2665 => "0000000010100111001001",
			2666 => "0000000010100111001001",
			2667 => "0010001010000100000100",
			2668 => "0000000010100111001001",
			2669 => "0000101111001100001000",
			2670 => "0000101101111000000100",
			2671 => "0000000010100111001001",
			2672 => "0000000010100111001001",
			2673 => "0000000010100111001001",
			2674 => "0010010101011100011000",
			2675 => "0000001011010000010100",
			2676 => "0011001110011000001100",
			2677 => "0011010110001100001000",
			2678 => "0000000100111100000100",
			2679 => "0000000010101001110101",
			2680 => "0000001010101001110101",
			2681 => "0000000010101001110101",
			2682 => "0000111001000100000100",
			2683 => "0000000010101001110101",
			2684 => "0000000010101001110101",
			2685 => "1111111010101001110101",
			2686 => "0000001101110100010100",
			2687 => "0010011001001000001000",
			2688 => "0000000011100000000100",
			2689 => "0000000010101001110101",
			2690 => "0000001010101001110101",
			2691 => "0011101101101100001000",
			2692 => "0001101111000000000100",
			2693 => "0000000010101001110101",
			2694 => "0000000010101001110101",
			2695 => "1111111010101001110101",
			2696 => "0000001010101000000100",
			2697 => "0000001010101001110101",
			2698 => "0000010111100100010100",
			2699 => "0001000101010100000100",
			2700 => "0000000010101001110101",
			2701 => "0000010001110000001000",
			2702 => "0001011011111000000100",
			2703 => "0000000010101001110101",
			2704 => "0000000010101001110101",
			2705 => "0001100100110000000100",
			2706 => "0000000010101001110101",
			2707 => "0000001010101001110101",
			2708 => "0000000010100100000100",
			2709 => "1111111010101001110101",
			2710 => "0000100110010100001000",
			2711 => "0010110101010100000100",
			2712 => "0000000010101001110101",
			2713 => "0000000010101001110101",
			2714 => "0001011101001000000100",
			2715 => "0000000010101001110101",
			2716 => "0000000010101001110101",
			2717 => "0001001001010000101100",
			2718 => "0000001010111100000100",
			2719 => "1111111010101011010001",
			2720 => "0000010110110100100100",
			2721 => "0010110101011100011000",
			2722 => "0001101110100000001100",
			2723 => "0001111100110000001000",
			2724 => "0011010110110100000100",
			2725 => "0000001010101011010001",
			2726 => "0000001010101011010001",
			2727 => "1111111010101011010001",
			2728 => "0011100000110100000100",
			2729 => "1111111010101011010001",
			2730 => "0001011011000000000100",
			2731 => "0000000010101011010001",
			2732 => "0000001010101011010001",
			2733 => "0010101011000000001000",
			2734 => "0011110000001000000100",
			2735 => "0000000010101011010001",
			2736 => "0000001010101011010001",
			2737 => "0000000010101011010001",
			2738 => "1111111010101011010001",
			2739 => "1111111010101011010001",
			2740 => "0011110100011000111100",
			2741 => "0000100010100100110000",
			2742 => "0001011101001000011000",
			2743 => "0010001111111100010000",
			2744 => "0010101000111000001100",
			2745 => "0011100100100100000100",
			2746 => "0000000010101110101101",
			2747 => "0011100010011000000100",
			2748 => "0000000010101110101101",
			2749 => "0000001010101110101101",
			2750 => "1111111010101110101101",
			2751 => "0011010110001100000100",
			2752 => "0000000010101110101101",
			2753 => "1111111010101110101101",
			2754 => "0000011000011000001000",
			2755 => "0001011000101000000100",
			2756 => "0000000010101110101101",
			2757 => "1111111010101110101101",
			2758 => "0001111000101000001100",
			2759 => "0010101000101000000100",
			2760 => "0000000010101110101101",
			2761 => "0010011010000100000100",
			2762 => "0000001010101110101101",
			2763 => "0000000010101110101101",
			2764 => "1111111010101110101101",
			2765 => "0000010001100100000100",
			2766 => "1111111010101110101101",
			2767 => "0000100110010100000100",
			2768 => "0000000010101110101101",
			2769 => "0000000010101110101101",
			2770 => "0011111001111000001100",
			2771 => "0001011000101000001000",
			2772 => "0011001010100100000100",
			2773 => "0000000010101110101101",
			2774 => "0000001010101110101101",
			2775 => "1111111010101110101101",
			2776 => "0011001100101000011100",
			2777 => "0010000101011100001100",
			2778 => "0000101010010100001000",
			2779 => "0001101010101100000100",
			2780 => "0000000010101110101101",
			2781 => "0000001010101110101101",
			2782 => "1111111010101110101101",
			2783 => "0011110101100100000100",
			2784 => "1111111010101110101101",
			2785 => "0011110011111100001000",
			2786 => "0000011001100000000100",
			2787 => "0000001010101110101101",
			2788 => "0000000010101110101101",
			2789 => "1111111010101110101101",
			2790 => "0010000011001000001000",
			2791 => "0000100101101000000100",
			2792 => "0000001010101110101101",
			2793 => "0000000010101110101101",
			2794 => "0000000010101110101101",
			2795 => "0001101101010001001000",
			2796 => "0000100100010100111000",
			2797 => "0011111011011100100000",
			2798 => "0011100001101100011100",
			2799 => "0011100000110100010000",
			2800 => "0000001011001000001000",
			2801 => "0011110001000000000100",
			2802 => "0000000010110010000001",
			2803 => "0000000010110010000001",
			2804 => "0000011000011000000100",
			2805 => "0000000010110010000001",
			2806 => "0000000010110010000001",
			2807 => "0000011001100000001000",
			2808 => "0000111000101000000100",
			2809 => "0000000010110010000001",
			2810 => "0000000010110010000001",
			2811 => "0000000010110010000001",
			2812 => "1111111010110010000001",
			2813 => "0011100011101100001000",
			2814 => "0001100100000100000100",
			2815 => "0000000010110010000001",
			2816 => "0000001010110010000001",
			2817 => "0001111001010100000100",
			2818 => "0000000010110010000001",
			2819 => "0011110000001000000100",
			2820 => "0000000010110010000001",
			2821 => "0001101000010100000100",
			2822 => "0000000010110010000001",
			2823 => "0000000010110010000001",
			2824 => "0010000101011100001100",
			2825 => "0000111000000000000100",
			2826 => "0000000010110010000001",
			2827 => "0010011100101000000100",
			2828 => "0000000010110010000001",
			2829 => "0000000010110010000001",
			2830 => "1111111010110010000001",
			2831 => "0011111011011000010100",
			2832 => "0011100110000100001100",
			2833 => "0000011101000000001000",
			2834 => "0000010111100100000100",
			2835 => "0000000010110010000001",
			2836 => "0000000010110010000001",
			2837 => "0000000010110010000001",
			2838 => "0011110100110100000100",
			2839 => "0000000010110010000001",
			2840 => "0000000010110010000001",
			2841 => "0001111100101100000100",
			2842 => "0000000010110010000001",
			2843 => "0000000010100000000100",
			2844 => "0000000010110010000001",
			2845 => "0010001000111000000100",
			2846 => "0000000010110010000001",
			2847 => "0000000010110010000001",
			2848 => "0011110100011000110100",
			2849 => "0000100010100100101000",
			2850 => "0000100011111000100000",
			2851 => "0001111001010100011100",
			2852 => "0001000011000000010000",
			2853 => "0001001001000100001000",
			2854 => "0010001111111100000100",
			2855 => "0000000010110101001101",
			2856 => "1111111010110101001101",
			2857 => "0000000100011000000100",
			2858 => "0000000010110101001101",
			2859 => "0000001010110101001101",
			2860 => "0011001100101000000100",
			2861 => "1111111010110101001101",
			2862 => "0000011001100000000100",
			2863 => "0000000010110101001101",
			2864 => "0000000010110101001101",
			2865 => "1111111010110101001101",
			2866 => "0010110011010000000100",
			2867 => "0000000010110101001101",
			2868 => "0000001010110101001101",
			2869 => "0000010001100100000100",
			2870 => "1111111010110101001101",
			2871 => "0000100110010100000100",
			2872 => "0000000010110101001101",
			2873 => "0000000010110101001101",
			2874 => "0011111001111000001100",
			2875 => "0001011000101000001000",
			2876 => "0011001010100100000100",
			2877 => "0000000010110101001101",
			2878 => "0000001010110101001101",
			2879 => "1111111010110101001101",
			2880 => "0011001100101000011100",
			2881 => "0010000101011100001100",
			2882 => "0000101010010100001000",
			2883 => "0001101010101100000100",
			2884 => "0000000010110101001101",
			2885 => "0000001010110101001101",
			2886 => "1111111010110101001101",
			2887 => "0011110101100100000100",
			2888 => "1111111010110101001101",
			2889 => "0011110011111100001000",
			2890 => "0000011001100000000100",
			2891 => "0000001010110101001101",
			2892 => "0000000010110101001101",
			2893 => "1111111010110101001101",
			2894 => "0010000011001000001000",
			2895 => "0001010110011100000100",
			2896 => "0000001010110101001101",
			2897 => "0000000010110101001101",
			2898 => "0000000010110101001101",
			2899 => "0011111000101100010100",
			2900 => "0010010110000000010000",
			2901 => "0011001100101000001100",
			2902 => "0000000100011000000100",
			2903 => "1111111010110111011001",
			2904 => "0001110011001000000100",
			2905 => "0000001010110111011001",
			2906 => "1111111010110111011001",
			2907 => "0000001010110111011001",
			2908 => "1111111010110111011001",
			2909 => "0000010110001100110000",
			2910 => "0000111101101000000100",
			2911 => "0000001010110111011001",
			2912 => "0011011011101100011000",
			2913 => "0011001010100100001100",
			2914 => "0010010101011100001000",
			2915 => "0000000100010100000100",
			2916 => "0000000010110111011001",
			2917 => "1111111010110111011001",
			2918 => "0000001010110111011001",
			2919 => "0011110000100100001000",
			2920 => "0000110011100100000100",
			2921 => "1111111010110111011001",
			2922 => "1111111010110111011001",
			2923 => "0000000010110111011001",
			2924 => "0000001101110100001000",
			2925 => "0010011001001000000100",
			2926 => "0000000010110111011001",
			2927 => "1111111010110111011001",
			2928 => "0010101100010000000100",
			2929 => "0000001010110111011001",
			2930 => "0001000110000000000100",
			2931 => "0000000010110111011001",
			2932 => "0000001010110111011001",
			2933 => "1111111010110111011001",
			2934 => "0000010111100100101100",
			2935 => "0010010101101100100100",
			2936 => "0011001010100100010000",
			2937 => "0001110011001000000100",
			2938 => "0000000010111010100101",
			2939 => "0010101101001000001000",
			2940 => "0000000110001000000100",
			2941 => "0000000010111010100101",
			2942 => "0000000010111010100101",
			2943 => "0000000010111010100101",
			2944 => "0001001001000100001100",
			2945 => "0000110011000000001000",
			2946 => "0010100011000000000100",
			2947 => "0000000010111010100101",
			2948 => "0000000010111010100101",
			2949 => "0000000010111010100101",
			2950 => "0001001101101000000100",
			2951 => "0000000010111010100101",
			2952 => "0000000010111010100101",
			2953 => "0011111000010100000100",
			2954 => "0000000010111010100101",
			2955 => "0000000010111010100101",
			2956 => "0001011111011000001100",
			2957 => "0011100110110000001000",
			2958 => "0011100010010100000100",
			2959 => "0000000010111010100101",
			2960 => "0000000010111010100101",
			2961 => "0000000010111010100101",
			2962 => "0011001001000100101000",
			2963 => "0000100100010100100000",
			2964 => "0001001010000100010000",
			2965 => "0011111100111100001000",
			2966 => "0001110011001000000100",
			2967 => "0000000010111010100101",
			2968 => "0000000010111010100101",
			2969 => "0000001000010000000100",
			2970 => "0000000010111010100101",
			2971 => "0000000010111010100101",
			2972 => "0011011010100100001000",
			2973 => "0001111101001000000100",
			2974 => "0000000010111010100101",
			2975 => "0000000010111010100101",
			2976 => "0001110110101100000100",
			2977 => "0000000010111010100101",
			2978 => "0000000010111010100101",
			2979 => "0001110001001000000100",
			2980 => "0000000010111010100101",
			2981 => "0000000010111010100101",
			2982 => "0010010011001000000100",
			2983 => "0000000010111010100101",
			2984 => "0000000010111010100101",
			2985 => "0000000011111000101000",
			2986 => "0001110110101100100100",
			2987 => "0011001110011000001000",
			2988 => "0000000000000100000100",
			2989 => "0000000010111101110001",
			2990 => "0000001010111101110001",
			2991 => "0011011010100100010000",
			2992 => "0010001001000100001000",
			2993 => "0011001010100100000100",
			2994 => "0000000010111101110001",
			2995 => "1111111010111101110001",
			2996 => "0000011000011000000100",
			2997 => "0000000010111101110001",
			2998 => "0000000010111101110001",
			2999 => "0001011001010100000100",
			3000 => "0000000010111101110001",
			3001 => "0001001111011000000100",
			3002 => "0000001010111101110001",
			3003 => "0000000010111101110001",
			3004 => "1111111010111101110001",
			3005 => "0000111000000000011100",
			3006 => "0011010111011100011000",
			3007 => "0000101011010000001000",
			3008 => "0011010110001100000100",
			3009 => "0000000010111101110001",
			3010 => "0000000010111101110001",
			3011 => "0011001010100100001000",
			3012 => "0010010101010100000100",
			3013 => "0000000010111101110001",
			3014 => "0000001010111101110001",
			3015 => "0001111001010100000100",
			3016 => "1111111010111101110001",
			3017 => "0000000010111101110001",
			3018 => "0000001010111101110001",
			3019 => "0000111100010000000100",
			3020 => "1111111010111101110001",
			3021 => "0000010011110000010000",
			3022 => "0001111001010100000100",
			3023 => "1111111010111101110001",
			3024 => "0001011101001000000100",
			3025 => "1111111010111101110001",
			3026 => "0010001001000100000100",
			3027 => "0000001010111101110001",
			3028 => "0000000010111101110001",
			3029 => "0001001100000000000100",
			3030 => "1111111010111101110001",
			3031 => "0011110010101000000100",
			3032 => "0000000010111101110001",
			3033 => "0001111100011100000100",
			3034 => "0000001010111101110001",
			3035 => "0000000010111101110001",
			3036 => "0010110011010000110000",
			3037 => "0001000110000000100100",
			3038 => "0010101101001000100000",
			3039 => "0001001001000100011100",
			3040 => "0000010110010000010000",
			3041 => "0011001010100100001000",
			3042 => "0000001001110100000100",
			3043 => "0000000011000000110101",
			3044 => "0000000011000000110101",
			3045 => "0000110110000000000100",
			3046 => "0000000011000000110101",
			3047 => "0000000011000000110101",
			3048 => "0011111110101100001000",
			3049 => "0010001111111100000100",
			3050 => "0000000011000000110101",
			3051 => "0000000011000000110101",
			3052 => "0000000011000000110101",
			3053 => "0000000011000000110101",
			3054 => "0000000011000000110101",
			3055 => "0010101001010100000100",
			3056 => "1111111011000000110101",
			3057 => "0000011000011000000100",
			3058 => "0000000011000000110101",
			3059 => "0000000011000000110101",
			3060 => "0011101101100000011000",
			3061 => "0001010011000100010100",
			3062 => "0011000111011100000100",
			3063 => "0000000011000000110101",
			3064 => "0001111000101000001000",
			3065 => "0011111110000000000100",
			3066 => "0000000011000000110101",
			3067 => "0000001011000000110101",
			3068 => "0000110011001000000100",
			3069 => "0000000011000000110101",
			3070 => "0000000011000000110101",
			3071 => "0000000011000000110101",
			3072 => "0001101010101100000100",
			3073 => "0000000011000000110101",
			3074 => "0000011001100000000100",
			3075 => "0000000011000000110101",
			3076 => "0001001100000000001000",
			3077 => "0000001101111000000100",
			3078 => "0000000011000000110101",
			3079 => "0000000011000000110101",
			3080 => "0000001110101000000100",
			3081 => "0000000011000000110101",
			3082 => "0000111011111000000100",
			3083 => "0000000011000000110101",
			3084 => "0000000011000000110101",
			3085 => "0011100000110100100100",
			3086 => "0001111000000000011000",
			3087 => "0001000101010100010000",
			3088 => "0000010110010000000100",
			3089 => "1111111011000011111001",
			3090 => "0000110101101100001000",
			3091 => "0000110111011100000100",
			3092 => "0000000011000011111001",
			3093 => "0000000011000011111001",
			3094 => "0000000011000011111001",
			3095 => "0001100000100000000100",
			3096 => "0000000011000011111001",
			3097 => "0000001011000011111001",
			3098 => "0010101010000100001000",
			3099 => "0010100101101100000100",
			3100 => "0000000011000011111001",
			3101 => "0000000011000011111001",
			3102 => "1111111011000011111001",
			3103 => "0010001001001100001000",
			3104 => "0000000110010100000100",
			3105 => "0000000011000011111001",
			3106 => "1111111011000011111001",
			3107 => "0000001101110100000100",
			3108 => "1111111011000011111001",
			3109 => "0011100111001000010100",
			3110 => "0001111000101000001100",
			3111 => "0001000101111000001000",
			3112 => "0011011110011000000100",
			3113 => "0000000011000011111001",
			3114 => "0000001011000011111001",
			3115 => "0000000011000011111001",
			3116 => "0011011100101000000100",
			3117 => "1111111011000011111001",
			3118 => "0000000011000011111001",
			3119 => "0010011101101000010000",
			3120 => "0000010001100100001000",
			3121 => "0011011011101100000100",
			3122 => "0000000011000011111001",
			3123 => "1111111011000011111001",
			3124 => "0010010101101100000100",
			3125 => "0000001011000011111001",
			3126 => "1111111011000011111001",
			3127 => "0010101011111000001000",
			3128 => "0010010011000000000100",
			3129 => "0000001011000011111001",
			3130 => "0000000011000011111001",
			3131 => "0001001100000000000100",
			3132 => "1111111011000011111001",
			3133 => "0000000011000011111001",
			3134 => "0011111011011100111000",
			3135 => "0001111001010100110100",
			3136 => "0001111101001000101000",
			3137 => "0000111100010000011100",
			3138 => "0001011000000000010000",
			3139 => "0001111000111000001000",
			3140 => "0011001010100100000100",
			3141 => "0000000011000111001101",
			3142 => "1111111011000111001101",
			3143 => "0000111001000100000100",
			3144 => "0000000011000111001101",
			3145 => "1111111011000111001101",
			3146 => "0010011001000100001000",
			3147 => "0000000100011000000100",
			3148 => "0000000011000111001101",
			3149 => "0000001011000111001101",
			3150 => "1111111011000111001101",
			3151 => "0000011001100000000100",
			3152 => "1111111011000111001101",
			3153 => "0000001010111100000100",
			3154 => "0000000011000111001101",
			3155 => "0000001011000111001101",
			3156 => "0000011000011000000100",
			3157 => "0000000011000111001101",
			3158 => "0010000000110000000100",
			3159 => "0000001011000111001101",
			3160 => "0000000011000111001101",
			3161 => "1111111011000111001101",
			3162 => "0001000111011100001100",
			3163 => "0001010101111000001000",
			3164 => "0011100110111000000100",
			3165 => "0000001011000111001101",
			3166 => "1111111011000111001101",
			3167 => "1111111011000111001101",
			3168 => "0000110011100100001100",
			3169 => "0011111000001000000100",
			3170 => "0000001011000111001101",
			3171 => "0001100010000100000100",
			3172 => "0000000011000111001101",
			3173 => "0000001011000111001101",
			3174 => "0000010011110000010100",
			3175 => "0010010110000000010000",
			3176 => "0010000101101100001000",
			3177 => "0011101111010100000100",
			3178 => "0000000011000111001101",
			3179 => "0000001011000111001101",
			3180 => "0000000110111100000100",
			3181 => "0000000011000111001101",
			3182 => "1111111011000111001101",
			3183 => "0000001011000111001101",
			3184 => "0000101101011000000100",
			3185 => "1111111011000111001101",
			3186 => "0000000011000111001101",
			3187 => "0001100100110000110100",
			3188 => "0001111000111000011100",
			3189 => "0001111111011000000100",
			3190 => "0000000011001011000001",
			3191 => "0010101000111000010000",
			3192 => "0011001010100100000100",
			3193 => "0000000011001011000001",
			3194 => "0000011000011000000100",
			3195 => "0000000011001011000001",
			3196 => "0010001111001000000100",
			3197 => "0000000011001011000001",
			3198 => "0000000011001011000001",
			3199 => "0011001100101000000100",
			3200 => "0000000011001011000001",
			3201 => "0000000011001011000001",
			3202 => "0000111111011000001100",
			3203 => "0000011001100100000100",
			3204 => "0000000011001011000001",
			3205 => "0000110110000000000100",
			3206 => "0000000011001011000001",
			3207 => "0000000011001011000001",
			3208 => "0010110111011100000100",
			3209 => "0000000011001011000001",
			3210 => "0010110101010100000100",
			3211 => "0000000011001011000001",
			3212 => "0000000011001011000001",
			3213 => "0011110011111101000000",
			3214 => "0001011001010100011000",
			3215 => "0010010101011100001000",
			3216 => "0000000110111100000100",
			3217 => "0000000011001011000001",
			3218 => "0000000011001011000001",
			3219 => "0000010001110000000100",
			3220 => "0000000011001011000001",
			3221 => "0001000111011100000100",
			3222 => "0000000011001011000001",
			3223 => "0000001100001000000100",
			3224 => "0000000011001011000001",
			3225 => "0000000011001011000001",
			3226 => "0011000101011100010000",
			3227 => "0011010101010100001100",
			3228 => "0011000011010000001000",
			3229 => "0011110110011000000100",
			3230 => "0000000011001011000001",
			3231 => "0000000011001011000001",
			3232 => "0000000011001011000001",
			3233 => "0000000011001011000001",
			3234 => "0010101011000000001100",
			3235 => "0000000101101000000100",
			3236 => "0000000011001011000001",
			3237 => "0010110101101100000100",
			3238 => "0000000011001011000001",
			3239 => "0000000011001011000001",
			3240 => "0010111001000100000100",
			3241 => "0000000011001011000001",
			3242 => "0001001100010000000100",
			3243 => "0000000011001011000001",
			3244 => "0000000011001011000001",
			3245 => "0001001100000000000100",
			3246 => "0000000011001011000001",
			3247 => "0000000011001011000001",
			3248 => "0001001001010000110100",
			3249 => "0001111111011000000100",
			3250 => "1111111011001100101101",
			3251 => "0000010110110100101100",
			3252 => "0010110111011100010100",
			3253 => "0010101111011000001000",
			3254 => "0000000101011000000100",
			3255 => "0000000011001100101101",
			3256 => "0000001011001100101101",
			3257 => "0001111000000100000100",
			3258 => "0000001011001100101101",
			3259 => "0000010110010000000100",
			3260 => "0000000011001100101101",
			3261 => "0000000011001100101101",
			3262 => "0001111000101000001100",
			3263 => "0010011101101000001000",
			3264 => "0001101010110100000100",
			3265 => "0000000011001100101101",
			3266 => "0000001011001100101101",
			3267 => "1111111011001100101101",
			3268 => "0011111011110100001000",
			3269 => "0001011000000000000100",
			3270 => "0000000011001100101101",
			3271 => "1111111011001100101101",
			3272 => "0000000011001100101101",
			3273 => "1111111011001100101101",
			3274 => "1111111011001100101101",
			3275 => "0010101011111001100000",
			3276 => "0001010011001000010000",
			3277 => "0001011111011000001100",
			3278 => "0001101010001000000100",
			3279 => "1111111011010000010001",
			3280 => "0011100100111000000100",
			3281 => "0000001011010000010001",
			3282 => "0000000011010000010001",
			3283 => "1111111011010000010001",
			3284 => "0000010111100100100100",
			3285 => "0010101000111000001100",
			3286 => "0001001100101000000100",
			3287 => "0000000011010000010001",
			3288 => "0000000110011000000100",
			3289 => "0000000011010000010001",
			3290 => "0000001011010000010001",
			3291 => "0010110011010000010000",
			3292 => "0011001110011000001000",
			3293 => "0001100101001100000100",
			3294 => "0000000011010000010001",
			3295 => "0000000011010000010001",
			3296 => "0000001011001000000100",
			3297 => "0000000011010000010001",
			3298 => "1111111011010000010001",
			3299 => "0001010110101100000100",
			3300 => "0000000011010000010001",
			3301 => "0000001011010000010001",
			3302 => "0001001010000100010100",
			3303 => "0011111100111100001000",
			3304 => "0001111000000100000100",
			3305 => "0000000011010000010001",
			3306 => "1111111011010000010001",
			3307 => "0000111000000000000100",
			3308 => "0000000011010000010001",
			3309 => "0010011101101000000100",
			3310 => "1111111011010000010001",
			3311 => "0000000011010000010001",
			3312 => "0000100110010100001100",
			3313 => "0010101000101000000100",
			3314 => "0000000011010000010001",
			3315 => "0001111000101000000100",
			3316 => "0000001011010000010001",
			3317 => "0000000011010000010001",
			3318 => "0001101010110000000100",
			3319 => "1111111011010000010001",
			3320 => "0000010011010000000100",
			3321 => "0000000011010000010001",
			3322 => "0000000011010000010001",
			3323 => "0011001001000100001100",
			3324 => "0000111011000000000100",
			3325 => "1111111011010000010001",
			3326 => "0011010101010100000100",
			3327 => "0000000011010000010001",
			3328 => "0000000011010000010001",
			3329 => "0010011000000100000100",
			3330 => "0000000011010000010001",
			3331 => "0000000011010000010001",
			3332 => "0010010101011100011000",
			3333 => "0000001011010000010100",
			3334 => "0011001110011000001100",
			3335 => "0010101000000000001000",
			3336 => "0000001100111000000100",
			3337 => "0000000011010011110101",
			3338 => "0000000011010011110101",
			3339 => "0000000011010011110101",
			3340 => "0000111001000100000100",
			3341 => "0000000011010011110101",
			3342 => "0000000011010011110101",
			3343 => "0000000011010011110101",
			3344 => "0001000011000000101100",
			3345 => "0011110011111100101000",
			3346 => "0011010110110100001000",
			3347 => "0010101111011000000100",
			3348 => "0000000011010011110101",
			3349 => "0000000011010011110101",
			3350 => "0000011001100000010000",
			3351 => "0001000111011100001000",
			3352 => "0001010101111000000100",
			3353 => "0000000011010011110101",
			3354 => "0000000011010011110101",
			3355 => "0000101110110100000100",
			3356 => "0000000011010011110101",
			3357 => "0000000011010011110101",
			3358 => "0001000101010100001000",
			3359 => "0000110011001000000100",
			3360 => "0000000011010011110101",
			3361 => "0000000011010011110101",
			3362 => "0010110111011100000100",
			3363 => "0000000011010011110101",
			3364 => "0000000011010011110101",
			3365 => "0000000011010011110101",
			3366 => "0001011100101100001100",
			3367 => "0010110101011100000100",
			3368 => "1111111011010011110101",
			3369 => "0010110101101100000100",
			3370 => "0000000011010011110101",
			3371 => "0000000011010011110101",
			3372 => "0000011000011000001100",
			3373 => "0010000101011100001000",
			3374 => "0000010111110000000100",
			3375 => "0000000011010011110101",
			3376 => "0000000011010011110101",
			3377 => "0000000011010011110101",
			3378 => "0010001010000100001100",
			3379 => "0011010101010100001000",
			3380 => "0001001111101000000100",
			3381 => "0000000011010011110101",
			3382 => "0000000011010011110101",
			3383 => "0000000011010011110101",
			3384 => "0010101011000000001000",
			3385 => "0000111111101000000100",
			3386 => "0000000011010011110101",
			3387 => "0000000011010011110101",
			3388 => "0000000011010011110101",
			3389 => "0010101111011000001000",
			3390 => "0011100010010100000100",
			3391 => "0000000011010111000001",
			3392 => "0000000011010111000001",
			3393 => "0001011100110000100100",
			3394 => "0011101001110000001000",
			3395 => "0011011110011000000100",
			3396 => "0000000011010111000001",
			3397 => "0000000011010111000001",
			3398 => "0011010111011100011000",
			3399 => "0011001010100100001100",
			3400 => "0010010101011100000100",
			3401 => "0000000011010111000001",
			3402 => "0010101101001000000100",
			3403 => "0000000011010111000001",
			3404 => "0000000011010111000001",
			3405 => "0000110011000000000100",
			3406 => "0000000011010111000001",
			3407 => "0010010101101100000100",
			3408 => "0000000011010111000001",
			3409 => "0000000011010111000001",
			3410 => "0000000011010111000001",
			3411 => "0000010111100100011000",
			3412 => "0011011110011000001000",
			3413 => "0000001110101000000100",
			3414 => "0000000011010111000001",
			3415 => "0000000011010111000001",
			3416 => "0001101000101100001100",
			3417 => "0000001011001000001000",
			3418 => "0000000000011100000100",
			3419 => "0000000011010111000001",
			3420 => "0000000011010111000001",
			3421 => "0000000011010111000001",
			3422 => "0000000011010111000001",
			3423 => "0001111000101000010000",
			3424 => "0000011000011000000100",
			3425 => "0000000011010111000001",
			3426 => "0000001101110100001000",
			3427 => "0001011100101100000100",
			3428 => "0000000011010111000001",
			3429 => "0000000011010111000001",
			3430 => "0000000011010111000001",
			3431 => "0011001001000100001100",
			3432 => "0011000111011100000100",
			3433 => "0000000011010111000001",
			3434 => "0001110001001000000100",
			3435 => "0000000011010111000001",
			3436 => "0000000011010111000001",
			3437 => "0010011000000100000100",
			3438 => "0000000011010111000001",
			3439 => "0000000011010111000001",
			3440 => "0001001001010000111100",
			3441 => "0001111111011000000100",
			3442 => "1111111011011000111111",
			3443 => "0010010011001000110100",
			3444 => "0010110111011100011000",
			3445 => "0010101111011000001000",
			3446 => "0000000101011000000100",
			3447 => "0000000011011000111111",
			3448 => "0000001011011000111111",
			3449 => "0000010110010000001000",
			3450 => "0000000000000000000100",
			3451 => "0000000011011000111111",
			3452 => "1111111011011000111111",
			3453 => "0000000110010100000100",
			3454 => "0000000011011000111111",
			3455 => "0000000011011000111111",
			3456 => "0001111000101000001100",
			3457 => "0010011101101000001000",
			3458 => "0001101010110100000100",
			3459 => "0000000011011000111111",
			3460 => "0000001011011000111111",
			3461 => "0000000011011000111111",
			3462 => "0001101010101100001000",
			3463 => "0010001010000100000100",
			3464 => "1111111011011000111111",
			3465 => "0000000011011000111111",
			3466 => "0001001111011000000100",
			3467 => "0000000011011000111111",
			3468 => "0000001011011000111111",
			3469 => "1111111011011000111111",
			3470 => "1111111011011000111111",
			3471 => "0011111000101100010000",
			3472 => "0010010110000000001100",
			3473 => "0010001001000100000100",
			3474 => "1111111011011010100001",
			3475 => "0011000011010000000100",
			3476 => "1111111011011010100001",
			3477 => "0000001011011010100001",
			3478 => "1111111011011010100001",
			3479 => "0000010110001100100000",
			3480 => "0010101111011000000100",
			3481 => "0000001011011010100001",
			3482 => "0010010101011100001000",
			3483 => "0001010011000000000100",
			3484 => "0000000011011010100001",
			3485 => "1111111011011010100001",
			3486 => "0000000010100100001000",
			3487 => "0001111001010100000100",
			3488 => "0000001011011010100001",
			3489 => "1111111011011010100001",
			3490 => "0010110101011100001000",
			3491 => "0010001001000100000100",
			3492 => "0000001011011010100001",
			3493 => "0000000011011010100001",
			3494 => "0000001011011010100001",
			3495 => "1111111011011010100001",
			3496 => "0011011110011000101000",
			3497 => "0000000100010100100000",
			3498 => "0001011000000000010100",
			3499 => "0000110011000000001100",
			3500 => "0011100010010100000100",
			3501 => "0000000011011100111101",
			3502 => "0000000101011000000100",
			3503 => "0000000011011100111101",
			3504 => "0000001011011100111101",
			3505 => "0001111000111000000100",
			3506 => "0000000011011100111101",
			3507 => "1111111011011100111101",
			3508 => "0000111100110000001000",
			3509 => "0001101001110000000100",
			3510 => "0000000011011100111101",
			3511 => "0000001011011100111101",
			3512 => "0000000011011100111101",
			3513 => "0000111111011000000100",
			3514 => "0000000011011100111101",
			3515 => "1111111011011100111101",
			3516 => "0000100011111000001100",
			3517 => "0001111001010100001000",
			3518 => "0011100110100000000100",
			3519 => "0000000011011100111101",
			3520 => "0000000011011100111101",
			3521 => "1111111011011100111101",
			3522 => "0001011101001000001000",
			3523 => "0000110011100100000100",
			3524 => "0000001011011100111101",
			3525 => "0000000011011100111101",
			3526 => "0000111100010000000100",
			3527 => "1111111011011100111101",
			3528 => "0000011001100000000100",
			3529 => "0000001011011100111101",
			3530 => "0011111010110000000100",
			3531 => "0000001011011100111101",
			3532 => "0001111001011000000100",
			3533 => "1111111011011100111101",
			3534 => "0000000011011100111101",
			3535 => "0001101100000100100000",
			3536 => "0000101010101000011000",
			3537 => "0001111001010100010100",
			3538 => "0011110111100000001100",
			3539 => "0011001100101000000100",
			3540 => "0000000011011111100001",
			3541 => "0010110101010100000100",
			3542 => "0000000011011111100001",
			3543 => "0000000011011111100001",
			3544 => "0000111101001000000100",
			3545 => "0000000011011111100001",
			3546 => "0000000011011111100001",
			3547 => "0000000011011111100001",
			3548 => "0001001000000000000100",
			3549 => "0000000011011111100001",
			3550 => "0000000011011111100001",
			3551 => "0011011110011000010100",
			3552 => "0000101100001000001000",
			3553 => "0000000010101100000100",
			3554 => "0000000011011111100001",
			3555 => "0000000011011111100001",
			3556 => "0001101101010000000100",
			3557 => "0000000011011111100001",
			3558 => "0000111000000000000100",
			3559 => "0000000011011111100001",
			3560 => "0000000011011111100001",
			3561 => "0000011001100000001000",
			3562 => "0011100111100000000100",
			3563 => "0000000011011111100001",
			3564 => "0000000011011111100001",
			3565 => "0000010001100100000100",
			3566 => "0000000011011111100001",
			3567 => "0000101111001100001100",
			3568 => "0001101011011100001000",
			3569 => "0010101011000000000100",
			3570 => "0000000011011111100001",
			3571 => "0000000011011111100001",
			3572 => "0000000011011111100001",
			3573 => "0011110011100000000100",
			3574 => "0000000011011111100001",
			3575 => "0000000011011111100001",
			3576 => "0010101000111000101000",
			3577 => "0001001100101000011000",
			3578 => "0011001010100100001100",
			3579 => "0001111000000100000100",
			3580 => "0000000011100010100101",
			3581 => "0000000101011000000100",
			3582 => "0000000011100010100101",
			3583 => "0000000011100010100101",
			3584 => "0000110011000000001000",
			3585 => "0001010110000000000100",
			3586 => "0000000011100010100101",
			3587 => "0000000011100010100101",
			3588 => "0000000011100010100101",
			3589 => "0001000110000000001000",
			3590 => "0001111111011000000100",
			3591 => "0000000011100010100101",
			3592 => "0000000011100010100101",
			3593 => "0000110011000000000100",
			3594 => "0000000011100010100101",
			3595 => "0000000011100010100101",
			3596 => "0010110111011100010100",
			3597 => "0000101011010000010000",
			3598 => "0000001100001000001100",
			3599 => "0001011001010100000100",
			3600 => "0000000011100010100101",
			3601 => "0001011000101000000100",
			3602 => "0000000011100010100101",
			3603 => "0000000011100010100101",
			3604 => "0000000011100010100101",
			3605 => "0000000011100010100101",
			3606 => "0010101011111000010100",
			3607 => "0001011001010000001100",
			3608 => "0011100111001000001000",
			3609 => "0010101101001000000100",
			3610 => "0000000011100010100101",
			3611 => "0000000011100010100101",
			3612 => "0000000011100010100101",
			3613 => "0000011111011100000100",
			3614 => "0000000011100010100101",
			3615 => "0000000011100010100101",
			3616 => "0011001001000100001100",
			3617 => "0010000101011100001000",
			3618 => "0000010111110000000100",
			3619 => "0000000011100010100101",
			3620 => "0000000011100010100101",
			3621 => "0000000011100010100101",
			3622 => "0010011000000100000100",
			3623 => "0000000011100010100101",
			3624 => "0000000011100010100101",
			3625 => "0010110101011100110100",
			3626 => "0001110100101100101100",
			3627 => "0000101111001100100100",
			3628 => "0011101111010100011000",
			3629 => "0011101101100000010000",
			3630 => "0010110011010000001000",
			3631 => "0001000110000000000100",
			3632 => "0000000011100100110001",
			3633 => "0000000011100100110001",
			3634 => "0001010011000100000100",
			3635 => "0000000011100100110001",
			3636 => "0000000011100100110001",
			3637 => "0010011100101000000100",
			3638 => "0000000011100100110001",
			3639 => "0000000011100100110001",
			3640 => "0000101100100100001000",
			3641 => "0001100100100000000100",
			3642 => "0000000011100100110001",
			3643 => "0000000011100100110001",
			3644 => "0000000011100100110001",
			3645 => "0011001010100100000100",
			3646 => "0000000011100100110001",
			3647 => "0000000011100100110001",
			3648 => "0000001010010000000100",
			3649 => "1111111011100100110001",
			3650 => "0000000011100100110001",
			3651 => "0011011100101000001100",
			3652 => "0010101000100000001000",
			3653 => "0011111100111100000100",
			3654 => "0000000011100100110001",
			3655 => "0000001011100100110001",
			3656 => "0000000011100100110001",
			3657 => "0000011001100000000100",
			3658 => "0000000011100100110001",
			3659 => "0000000011100100110001",
			3660 => "0001011100110000110000",
			3661 => "0011001010100100010100",
			3662 => "0000001001110100001000",
			3663 => "0000000110001000000100",
			3664 => "0000000011100111110101",
			3665 => "0000000011100111110101",
			3666 => "0001100101001100000100",
			3667 => "0000000011100111110101",
			3668 => "0011100110111000000100",
			3669 => "0000000011100111110101",
			3670 => "0000000011100111110101",
			3671 => "0000110011000000001000",
			3672 => "0000101011110100000100",
			3673 => "0000000011100111110101",
			3674 => "0000000011100111110101",
			3675 => "0011111011011000010000",
			3676 => "0010110101011100001000",
			3677 => "0000110101111000000100",
			3678 => "0000000011100111110101",
			3679 => "1111111011100111110101",
			3680 => "0010010011000000000100",
			3681 => "0000000011100111110101",
			3682 => "0000000011100111110101",
			3683 => "0000000011100111110101",
			3684 => "0010110011010000010100",
			3685 => "0001011000101000010000",
			3686 => "0010101001010100001000",
			3687 => "0001111100110000000100",
			3688 => "0000000011100111110101",
			3689 => "0000000011100111110101",
			3690 => "0000010111100100000100",
			3691 => "0000000011100111110101",
			3692 => "0000000011100111110101",
			3693 => "0000000011100111110101",
			3694 => "0000010111100100001000",
			3695 => "0011110111000000000100",
			3696 => "0000000011100111110101",
			3697 => "0000001011100111110101",
			3698 => "0001111000101000001100",
			3699 => "0000011000011000000100",
			3700 => "0000000011100111110101",
			3701 => "0010011101101000000100",
			3702 => "0000000011100111110101",
			3703 => "0000000011100111110101",
			3704 => "0001111001011000000100",
			3705 => "0000000011100111110101",
			3706 => "0011011100101000000100",
			3707 => "0000000011100111110101",
			3708 => "0000000011100111110101",
			3709 => "0011110111100000010100",
			3710 => "0010010110000000010000",
			3711 => "0011001100101000001100",
			3712 => "0000000100011000000100",
			3713 => "1111111011101001111001",
			3714 => "0010101001010100000100",
			3715 => "0000001011101001111001",
			3716 => "1111111011101001111001",
			3717 => "0000001011101001111001",
			3718 => "1111111011101001111001",
			3719 => "0000010110001100101100",
			3720 => "0000111001010100100000",
			3721 => "0010010101011100001100",
			3722 => "0000000100010100001000",
			3723 => "0000010111110000000100",
			3724 => "0000001011101001111001",
			3725 => "0000000011101001111001",
			3726 => "1111111011101001111001",
			3727 => "0000000101011000000100",
			3728 => "1111111011101001111001",
			3729 => "0000010001110000001000",
			3730 => "0000111000000000000100",
			3731 => "0000000011101001111001",
			3732 => "1111111011101001111001",
			3733 => "0001111000101000000100",
			3734 => "0000010011101001111001",
			3735 => "0000001011101001111001",
			3736 => "0000000101101000000100",
			3737 => "1111111011101001111001",
			3738 => "0010110111011100000100",
			3739 => "1111111011101001111001",
			3740 => "0000001011101001111001",
			3741 => "1111111011101001111001",
			3742 => "0011110111100000010000",
			3743 => "0010010110000000001100",
			3744 => "0010001001000100000100",
			3745 => "1111111011101100010101",
			3746 => "0011000011010000000100",
			3747 => "1111111011101100010101",
			3748 => "0000001011101100010101",
			3749 => "1111111011101100010101",
			3750 => "0000111000000000011100",
			3751 => "0011010111011100010100",
			3752 => "0011110001100000000100",
			3753 => "0000011011101100010101",
			3754 => "0010001001000100001100",
			3755 => "0000110011100100001000",
			3756 => "0000000100010100000100",
			3757 => "0000001011101100010101",
			3758 => "0000000011101100010101",
			3759 => "0000010011101100010101",
			3760 => "1111111011101100010101",
			3761 => "0011011001001000000100",
			3762 => "0000010011101100010101",
			3763 => "1111111011101100010101",
			3764 => "0010001010000100011100",
			3765 => "0010110111011100010000",
			3766 => "0000000100010100001100",
			3767 => "0010101111101000001000",
			3768 => "0001011100010000000100",
			3769 => "1111111011101100010101",
			3770 => "0000001011101100010101",
			3771 => "1111111011101100010101",
			3772 => "1111111011101100010101",
			3773 => "0010101001000000001000",
			3774 => "0000011001100000000100",
			3775 => "0000001011101100010101",
			3776 => "0000000011101100010101",
			3777 => "1111111011101100010101",
			3778 => "0000011101000000000100",
			3779 => "0000000011101100010101",
			3780 => "1111111011101100010101",
			3781 => "0011101101100000110100",
			3782 => "0011100000110100010100",
			3783 => "0011001110011000001000",
			3784 => "0001110101111000000100",
			3785 => "0000000011101111011001",
			3786 => "0000000011101111011001",
			3787 => "0001110011001000001000",
			3788 => "0001111111011000000100",
			3789 => "0000000011101111011001",
			3790 => "0000000011101111011001",
			3791 => "0000000011101111011001",
			3792 => "0001000101111000010100",
			3793 => "0011001110011000001000",
			3794 => "0000000011001100000100",
			3795 => "0000000011101111011001",
			3796 => "0000000011101111011001",
			3797 => "0011010110001100000100",
			3798 => "0000000011101111011001",
			3799 => "0001111000101000000100",
			3800 => "0000000011101111011001",
			3801 => "0000000011101111011001",
			3802 => "0001001001010100000100",
			3803 => "0000000011101111011001",
			3804 => "0011010101010100000100",
			3805 => "0000000011101111011001",
			3806 => "0000000011101111011001",
			3807 => "0010011101101000010100",
			3808 => "0000001000110000010000",
			3809 => "0011001010100100001000",
			3810 => "0000111000000000000100",
			3811 => "0000000011101111011001",
			3812 => "0000000011101111011001",
			3813 => "0001011111011000000100",
			3814 => "0000000011101111011001",
			3815 => "0000000011101111011001",
			3816 => "0000000011101111011001",
			3817 => "0000011001100000000100",
			3818 => "0000000011101111011001",
			3819 => "0011110011100000010100",
			3820 => "0011000110000000001100",
			3821 => "0000101000010000001000",
			3822 => "0000100110010100000100",
			3823 => "0000000011101111011001",
			3824 => "0000000011101111011001",
			3825 => "0000000011101111011001",
			3826 => "0010011000000000000100",
			3827 => "0000000011101111011001",
			3828 => "0000000011101111011001",
			3829 => "0000000011101111011001",
			3830 => "0011111011011100101000",
			3831 => "0001011001010100011000",
			3832 => "0011001010100100001100",
			3833 => "0001111000111000001000",
			3834 => "0001110011001000000100",
			3835 => "0000000011110010011101",
			3836 => "0000000011110010011101",
			3837 => "0000000011110010011101",
			3838 => "0000110110000000001000",
			3839 => "0000111001000100000100",
			3840 => "0000000011110010011101",
			3841 => "0000000011110010011101",
			3842 => "0000000011110010011101",
			3843 => "0000011000011000001000",
			3844 => "0010011001001000000100",
			3845 => "0000000011110010011101",
			3846 => "0000000011110010011101",
			3847 => "0010010110000000000100",
			3848 => "0000000011110010011101",
			3849 => "0000000011110010011101",
			3850 => "0011100111001000010100",
			3851 => "0001011001010100001100",
			3852 => "0011010110001100001000",
			3853 => "0011011101000000000100",
			3854 => "0000000011110010011101",
			3855 => "0000000011110010011101",
			3856 => "0000000011110010011101",
			3857 => "0001010100101100000100",
			3858 => "0000000011110010011101",
			3859 => "0000000011110010011101",
			3860 => "0011101111010100000100",
			3861 => "0000000011110010011101",
			3862 => "0000001011001100001100",
			3863 => "0001101110001000001000",
			3864 => "0001100101001100000100",
			3865 => "0000000011110010011101",
			3866 => "0000000011110010011101",
			3867 => "0000000011110010011101",
			3868 => "0000001010111000001100",
			3869 => "0001110100101100000100",
			3870 => "0000000011110010011101",
			3871 => "0011001001001000000100",
			3872 => "0000000011110010011101",
			3873 => "0000000011110010011101",
			3874 => "0001110100101100000100",
			3875 => "0000000011110010011101",
			3876 => "0010001010000100000100",
			3877 => "0000000011110010011101",
			3878 => "0000000011110010011101",
			3879 => "0011111000101100010000",
			3880 => "0010010110000000001100",
			3881 => "0010001001000100000100",
			3882 => "1111111011110100010001",
			3883 => "0001011000111000000100",
			3884 => "1111111011110100010001",
			3885 => "0000010011110100010001",
			3886 => "1111111011110100010001",
			3887 => "0000010110001100101000",
			3888 => "0000111101101000000100",
			3889 => "0000010011110100010001",
			3890 => "0000000010100100001000",
			3891 => "0001110110101100000100",
			3892 => "0000001011110100010001",
			3893 => "1111111011110100010001",
			3894 => "0011011110011000010000",
			3895 => "0000000100010100001000",
			3896 => "0001100100110000000100",
			3897 => "0000001011110100010001",
			3898 => "0000010011110100010001",
			3899 => "0001101101010000000100",
			3900 => "1111111011110100010001",
			3901 => "0000000011110100010001",
			3902 => "0011101101100000000100",
			3903 => "0000011011110100010001",
			3904 => "0011111011110100000100",
			3905 => "1111111011110100010001",
			3906 => "0000001011110100010001",
			3907 => "1111111011110100010001",
			3908 => "0011110000100101001000",
			3909 => "0000110011001000100000",
			3910 => "0001010011001000010000",
			3911 => "0010100011000000001000",
			3912 => "0011111000101100000100",
			3913 => "0000000011110111011101",
			3914 => "0000000011110111011101",
			3915 => "0000110110000000000100",
			3916 => "0000000011110111011101",
			3917 => "0000000011110111011101",
			3918 => "0000010111100100001000",
			3919 => "0000000001110100000100",
			3920 => "0000000011110111011101",
			3921 => "0000000011110111011101",
			3922 => "0001001001000100000100",
			3923 => "0000000011110111011101",
			3924 => "0000000011110111011101",
			3925 => "0000000101101000100000",
			3926 => "0000011000011000001100",
			3927 => "0000001011001000001000",
			3928 => "0011110111100000000100",
			3929 => "0000000011110111011101",
			3930 => "0000000011110111011101",
			3931 => "0000000011110111011101",
			3932 => "0001111000101000010000",
			3933 => "0000010011110000001000",
			3934 => "0010001010000100000100",
			3935 => "0000000011110111011101",
			3936 => "0000000011110111011101",
			3937 => "0001011001010000000100",
			3938 => "0000000011110111011101",
			3939 => "0000000011110111011101",
			3940 => "0000000011110111011101",
			3941 => "0000101101110000000100",
			3942 => "0000000011110111011101",
			3943 => "0000000011110111011101",
			3944 => "0011011011101100001000",
			3945 => "0000111000000000000100",
			3946 => "0000000011110111011101",
			3947 => "0000000011110111011101",
			3948 => "0010110101011100010000",
			3949 => "0010010101101100001000",
			3950 => "0000011000011000000100",
			3951 => "0000000011110111011101",
			3952 => "0000000011110111011101",
			3953 => "0010100100101100000100",
			3954 => "0000000011110111011101",
			3955 => "0000000011110111011101",
			3956 => "0010010011001000000100",
			3957 => "0000000011110111011101",
			3958 => "0000000011110111011101",
			3959 => "0011111011011100111100",
			3960 => "0001011000111000100000",
			3961 => "0001111000111000010100",
			3962 => "0001010011001000001100",
			3963 => "0001001011101100001000",
			3964 => "0001010101101100000100",
			3965 => "0000000011111011000001",
			3966 => "0000000011111011000001",
			3967 => "0000000011111011000001",
			3968 => "0011001010100100000100",
			3969 => "0000000011111011000001",
			3970 => "0000000011111011000001",
			3971 => "0010100011000000001000",
			3972 => "0001001011101100000100",
			3973 => "0000000011111011000001",
			3974 => "0000000011111011000001",
			3975 => "0000000011111011000001",
			3976 => "0001000011000000010000",
			3977 => "0010111110011000000100",
			3978 => "0000000011111011000001",
			3979 => "0011110001100000001000",
			3980 => "0001011100110000000100",
			3981 => "0000000011111011000001",
			3982 => "0000000011111011000001",
			3983 => "0000000011111011000001",
			3984 => "0011100101110000001000",
			3985 => "0000101000110100000100",
			3986 => "0000000011111011000001",
			3987 => "0000000011111011000001",
			3988 => "0000000011111011000001",
			3989 => "0011010111011100100100",
			3990 => "0000100110010100001000",
			3991 => "0001111000101000000100",
			3992 => "0000000011111011000001",
			3993 => "0000000011111011000001",
			3994 => "0001101010101100001100",
			3995 => "0001111001010100001000",
			3996 => "0000011001100100000100",
			3997 => "0000000011111011000001",
			3998 => "0000000011111011000001",
			3999 => "0000000011111011000001",
			4000 => "0000101101111000001000",
			4001 => "0011100100101000000100",
			4002 => "0000000011111011000001",
			4003 => "0000000011111011000001",
			4004 => "0001110001010000000100",
			4005 => "0000000011111011000001",
			4006 => "0000000011111011000001",
			4007 => "0001000110000000000100",
			4008 => "0000000011111011000001",
			4009 => "0001001100000000001000",
			4010 => "0000001000001100000100",
			4011 => "0000000011111011000001",
			4012 => "0000000011111011000001",
			4013 => "0010010011001000000100",
			4014 => "0000000011111011000001",
			4015 => "0000000011111011000001",
			4016 => "0011111000101100010000",
			4017 => "0010010110000000001100",
			4018 => "0010001001000100000100",
			4019 => "1111111011111101000101",
			4020 => "0011000011010000000100",
			4021 => "1111111011111101000101",
			4022 => "0000001011111101000101",
			4023 => "1111111011111101000101",
			4024 => "0010000011001000110000",
			4025 => "0011010110001100001100",
			4026 => "0010101111011000000100",
			4027 => "0000001011111101000101",
			4028 => "0011110100111100000100",
			4029 => "1111111011111101000101",
			4030 => "0000000011111101000101",
			4031 => "0011100111001000010000",
			4032 => "0011111100111100001100",
			4033 => "0001111000101000001000",
			4034 => "0001010011000100000100",
			4035 => "0000001011111101000101",
			4036 => "1111111011111101000101",
			4037 => "1111111011111101000101",
			4038 => "0000001011111101000101",
			4039 => "0011000101101100010000",
			4040 => "0010001111001000001000",
			4041 => "0001000110000000000100",
			4042 => "0000000011111101000101",
			4043 => "0000001011111101000101",
			4044 => "0001011100010000000100",
			4045 => "0000000011111101000101",
			4046 => "1111111011111101000101",
			4047 => "0000001011111101000101",
			4048 => "1111111011111101000101",
			4049 => "0011100000110100011000",
			4050 => "0000010110010000000100",
			4051 => "0000000011111111101001",
			4052 => "0011100010010100001100",
			4053 => "0011101101101100001000",
			4054 => "0000001010111100000100",
			4055 => "0000000011111111101001",
			4056 => "0000000011111111101001",
			4057 => "0000000011111111101001",
			4058 => "0011101111000100000100",
			4059 => "0000000011111111101001",
			4060 => "0000000011111111101001",
			4061 => "0001101110000100110000",
			4062 => "0001011111011000001000",
			4063 => "0000001101110100000100",
			4064 => "0000000011111111101001",
			4065 => "0000000011111111101001",
			4066 => "0000010001110000001100",
			4067 => "0001011100101100001000",
			4068 => "0011100011011000000100",
			4069 => "0000000011111111101001",
			4070 => "0000000011111111101001",
			4071 => "0000000011111111101001",
			4072 => "0000010111100100001100",
			4073 => "0001001100101000000100",
			4074 => "0000000011111111101001",
			4075 => "0001100100110000000100",
			4076 => "0000000011111111101001",
			4077 => "0000000011111111101001",
			4078 => "0000100100010100001000",
			4079 => "0010011001001000000100",
			4080 => "0000000011111111101001",
			4081 => "0000000011111111101001",
			4082 => "0011100001000000000100",
			4083 => "0000000011111111101001",
			4084 => "0000000011111111101001",
			4085 => "0001111100101100000100",
			4086 => "0000000011111111101001",
			4087 => "0000000010100000000100",
			4088 => "0000000011111111101001",
			4089 => "0000000011111111101001",
			4090 => "0000011111011101001100",
			4091 => "0001000111011100100000",
			4092 => "0010110011010000010100",
			4093 => "0011101100011000010000",
			4094 => "0001100110000100001100",
			4095 => "0000110101101100001000",
			4096 => "0001010101011100000100",
			4097 => "0000000100000010100101",
			4098 => "0000000100000010100101",
			4099 => "1111111100000010100101",
			4100 => "0000001100000010100101",
			4101 => "1111111100000010100101",
			4102 => "0000110011000000001000",
			4103 => "0001010110000000000100",
			4104 => "0000000100000010100101",
			4105 => "0000000100000010100101",
			4106 => "1111111100000010100101",
			4107 => "0011101111010100011000",
			4108 => "0011111011110100010100",
			4109 => "0001100101001100010000",
			4110 => "0011100011101100001000",
			4111 => "0000010011110000000100",
			4112 => "0000000100000010100101",
			4113 => "1111111100000010100101",
			4114 => "0001111000101000000100",
			4115 => "1111111100000010100101",
			4116 => "0000000100000010100101",
			4117 => "0000001100000010100101",
			4118 => "1111111100000010100101",
			4119 => "0011101101100100001000",
			4120 => "0000010111100100000100",
			4121 => "0000001100000010100101",
			4122 => "0000000100000010100101",
			4123 => "0000001110110000000100",
			4124 => "1111111100000010100101",
			4125 => "0011111011011000000100",
			4126 => "0000000100000010100101",
			4127 => "0000000100000010100101",
			4128 => "0001011100000000001100",
			4129 => "0001110100101100000100",
			4130 => "0000000100000010100101",
			4131 => "0011001000000100000100",
			4132 => "0000000100000010100101",
			4133 => "0000000100000010100101",
			4134 => "0011110011100000000100",
			4135 => "1111111100000010100101",
			4136 => "0000000100000010100101",
			4137 => "0010001010000101000100",
			4138 => "0001101101010000110000",
			4139 => "0000000111111000101000",
			4140 => "0011111011011100011000",
			4141 => "0000100111000100010000",
			4142 => "0001000011000000001000",
			4143 => "0001011000000100000100",
			4144 => "0000000100000101010001",
			4145 => "0000000100000101010001",
			4146 => "0010001111001000000100",
			4147 => "0000000100000101010001",
			4148 => "0000000100000101010001",
			4149 => "0001001010000100000100",
			4150 => "0000000100000101010001",
			4151 => "0000000100000101010001",
			4152 => "0001111000101000001100",
			4153 => "0011100111001000001000",
			4154 => "0010001001001100000100",
			4155 => "0000000100000101010001",
			4156 => "0000001100000101010001",
			4157 => "0000000100000101010001",
			4158 => "0000000100000101010001",
			4159 => "0010110011010000000100",
			4160 => "1111111100000101010001",
			4161 => "0000000100000101010001",
			4162 => "0001000111011100001000",
			4163 => "0000000101101000000100",
			4164 => "0000000100000101010001",
			4165 => "0000000100000101010001",
			4166 => "0000001011001100000100",
			4167 => "0000000100000101010001",
			4168 => "0010101000101000000100",
			4169 => "0000001100000101010001",
			4170 => "0000000100000101010001",
			4171 => "0010101101001000010000",
			4172 => "0000010110110100001100",
			4173 => "0010110101011100000100",
			4174 => "0000000100000101010001",
			4175 => "0000000100111000000100",
			4176 => "0000000100000101010001",
			4177 => "0000000100000101010001",
			4178 => "0000000100000101010001",
			4179 => "1111111100000101010001",
			4180 => "0011111110000000000100",
			4181 => "1111111100000111001101",
			4182 => "0000010011110000100000",
			4183 => "0001001001010000011100",
			4184 => "0011010111011100011000",
			4185 => "0000000100010100001100",
			4186 => "0001111000101000001000",
			4187 => "0000011000011000000100",
			4188 => "0000000100000111001101",
			4189 => "0000001100000111001101",
			4190 => "1111111100000111001101",
			4191 => "0011100010110000000100",
			4192 => "1111111100000111001101",
			4193 => "0010101011111000000100",
			4194 => "0000000100000111001101",
			4195 => "1111111100000111001101",
			4196 => "0000001100000111001101",
			4197 => "1111111100000111001101",
			4198 => "0000111100010000010000",
			4199 => "0011000011010000000100",
			4200 => "1111111100000111001101",
			4201 => "0000001011111100000100",
			4202 => "1111111100000111001101",
			4203 => "0001000011000000000100",
			4204 => "0000001100000111001101",
			4205 => "1111111100000111001101",
			4206 => "0011001001000100000100",
			4207 => "1111111100000111001101",
			4208 => "0011011001001000000100",
			4209 => "0000001100000111001101",
			4210 => "1111111100000111001101",
			4211 => "0011000101010100111100",
			4212 => "0010101000111000010100",
			4213 => "0000110011001000010000",
			4214 => "0001111111011000000100",
			4215 => "0000000100001010010001",
			4216 => "0000000001110100001000",
			4217 => "0011101101000100000100",
			4218 => "0000000100001010010001",
			4219 => "0000000100001010010001",
			4220 => "0000000100001010010001",
			4221 => "0000000100001010010001",
			4222 => "0000010001100100011100",
			4223 => "0000101100010100001100",
			4224 => "0011101001011100000100",
			4225 => "0000000100001010010001",
			4226 => "0011101101100000000100",
			4227 => "0000000100001010010001",
			4228 => "0000000100001010010001",
			4229 => "0000011001100100000100",
			4230 => "0000000100001010010001",
			4231 => "0001011000000100001000",
			4232 => "0001011111011000000100",
			4233 => "0000000100001010010001",
			4234 => "0000000100001010010001",
			4235 => "0000000100001010010001",
			4236 => "0000011101000000001000",
			4237 => "0011100100111000000100",
			4238 => "0000000100001010010001",
			4239 => "0000000100001010010001",
			4240 => "0000000100001010010001",
			4241 => "0001011100010000001100",
			4242 => "0001011100000000001000",
			4243 => "0001010011000000000100",
			4244 => "0000000100001010010001",
			4245 => "0000000100001010010001",
			4246 => "0000000100001010010001",
			4247 => "0001011100011100011000",
			4248 => "0000010110110100010100",
			4249 => "0000001100001000001100",
			4250 => "0000001010101100000100",
			4251 => "0000000100001010010001",
			4252 => "0011010111011100000100",
			4253 => "0000000100001010010001",
			4254 => "0000000100001010010001",
			4255 => "0010101111101000000100",
			4256 => "0000000100001010010001",
			4257 => "0000000100001010010001",
			4258 => "0000000100001010010001",
			4259 => "0000000100001010010001",
			4260 => "0000000011111000101000",
			4261 => "0001110110101100100100",
			4262 => "0011001110011000001000",
			4263 => "0000000000000100000100",
			4264 => "0000000100001101001101",
			4265 => "0000001100001101001101",
			4266 => "0011011010100100010000",
			4267 => "0010001001000100001000",
			4268 => "0011001010100100000100",
			4269 => "0000000100001101001101",
			4270 => "1111111100001101001101",
			4271 => "0000011000011000000100",
			4272 => "0000000100001101001101",
			4273 => "0000000100001101001101",
			4274 => "0001011001010100000100",
			4275 => "0000000100001101001101",
			4276 => "0001001111011000000100",
			4277 => "0000001100001101001101",
			4278 => "0000000100001101001101",
			4279 => "1111111100001101001101",
			4280 => "0000100000101000100100",
			4281 => "0001111000101000011100",
			4282 => "0011100101110100001000",
			4283 => "0000000011001100000100",
			4284 => "0000000100001101001101",
			4285 => "1111111100001101001101",
			4286 => "0011100011101100001000",
			4287 => "0001100100110000000100",
			4288 => "0000000100001101001101",
			4289 => "0000001100001101001101",
			4290 => "0001100101001100000100",
			4291 => "1111111100001101001101",
			4292 => "0000010111110000000100",
			4293 => "0000000100001101001101",
			4294 => "0000000100001101001101",
			4295 => "0001011000000000000100",
			4296 => "0000000100001101001101",
			4297 => "1111111100001101001101",
			4298 => "0001110001010000000100",
			4299 => "1111111100001101001101",
			4300 => "0010011101101000000100",
			4301 => "0000000100001101001101",
			4302 => "0000011101000000000100",
			4303 => "0000000100001101001101",
			4304 => "0000101101011000000100",
			4305 => "1111111100001101001101",
			4306 => "0000000100001101001101",
			4307 => "0010101000111000101000",
			4308 => "0011111011011100100000",
			4309 => "0001111000111000010100",
			4310 => "0001111111011000000100",
			4311 => "0000000100010000101001",
			4312 => "0011001010100100000100",
			4313 => "0000000100010000101001",
			4314 => "0000011000011000000100",
			4315 => "0000000100010000101001",
			4316 => "0010001111001000000100",
			4317 => "0000000100010000101001",
			4318 => "0000000100010000101001",
			4319 => "0000110110000000001000",
			4320 => "0001010101101100000100",
			4321 => "0000000100010000101001",
			4322 => "0000000100010000101001",
			4323 => "0000000100010000101001",
			4324 => "0011101100011000000100",
			4325 => "0000000100010000101001",
			4326 => "0000000100010000101001",
			4327 => "0010110111011100100000",
			4328 => "0000010001100100011000",
			4329 => "0001011000000100001000",
			4330 => "0000110011100100000100",
			4331 => "0000000100010000101001",
			4332 => "0000000100010000101001",
			4333 => "0000111011111000001000",
			4334 => "0000011000111100000100",
			4335 => "0000000100010000101001",
			4336 => "0000000100010000101001",
			4337 => "0010101001011000000100",
			4338 => "0000000100010000101001",
			4339 => "0000000100010000101001",
			4340 => "0010010101101100000100",
			4341 => "0000000100010000101001",
			4342 => "0000000100010000101001",
			4343 => "0000000101101000011000",
			4344 => "0001111000101000001100",
			4345 => "0001011011000000001000",
			4346 => "0010011010000100000100",
			4347 => "0000000100010000101001",
			4348 => "0000000100010000101001",
			4349 => "0000000100010000101001",
			4350 => "0001011110111000000100",
			4351 => "0000000100010000101001",
			4352 => "0001001101001000000100",
			4353 => "0000000100010000101001",
			4354 => "0000000100010000101001",
			4355 => "0010001010000100000100",
			4356 => "0000000100010000101001",
			4357 => "0000101111001100001000",
			4358 => "0000101101111000000100",
			4359 => "0000000100010000101001",
			4360 => "0000000100010000101001",
			4361 => "0000000100010000101001",
			4362 => "0000010011110001001100",
			4363 => "0001000101010100011000",
			4364 => "0010101111011000001000",
			4365 => "0001100100101000000100",
			4366 => "0000000100010011101101",
			4367 => "0000000100010011101101",
			4368 => "0000011001100000001100",
			4369 => "0010111011101100000100",
			4370 => "0000000100010011101101",
			4371 => "0001001011101100000100",
			4372 => "0000000100010011101101",
			4373 => "0000000100010011101101",
			4374 => "0000000100010011101101",
			4375 => "0000010001110000010100",
			4376 => "0010101100010000001000",
			4377 => "0000011000111100000100",
			4378 => "0000000100010011101101",
			4379 => "0000000100010011101101",
			4380 => "0011011011101100001000",
			4381 => "0010110111011100000100",
			4382 => "0000000100010011101101",
			4383 => "0000000100010011101101",
			4384 => "0000000100010011101101",
			4385 => "0011111000100100011100",
			4386 => "0011100010110000001100",
			4387 => "0000000011001100001000",
			4388 => "0011010011010000000100",
			4389 => "0000000100010011101101",
			4390 => "0000000100010011101101",
			4391 => "0000000100010011101101",
			4392 => "0011011110011000001000",
			4393 => "0011001110011000000100",
			4394 => "0000000100010011101101",
			4395 => "0000000100010011101101",
			4396 => "0000011001100000000100",
			4397 => "0000000100010011101101",
			4398 => "0000000100010011101101",
			4399 => "0000000100010011101101",
			4400 => "0000110011100100001000",
			4401 => "0000001101011100000100",
			4402 => "0000000100010011101101",
			4403 => "0000000100010011101101",
			4404 => "0000101101011000001100",
			4405 => "0001110110101100001000",
			4406 => "0000000010110100000100",
			4407 => "0000000100010011101101",
			4408 => "0000000100010011101101",
			4409 => "0000000100010011101101",
			4410 => "0000000100010011101101",
			4411 => "0011011110011000110000",
			4412 => "0010101000000000010000",
			4413 => "0001111111011000000100",
			4414 => "0000000100010110111001",
			4415 => "0000000100011000000100",
			4416 => "0000000100010110111001",
			4417 => "0010101111011000000100",
			4418 => "0000000100010110111001",
			4419 => "0000000100010110111001",
			4420 => "0000010001100100011100",
			4421 => "0010010101101100010100",
			4422 => "0010111110011000010000",
			4423 => "0001101101010000001000",
			4424 => "0011100110100000000100",
			4425 => "0000000100010110111001",
			4426 => "0000000100010110111001",
			4427 => "0000000101101000000100",
			4428 => "0000000100010110111001",
			4429 => "0000000100010110111001",
			4430 => "0000000100010110111001",
			4431 => "0000111000000000000100",
			4432 => "0000000100010110111001",
			4433 => "0000000100010110111001",
			4434 => "0000000100010110111001",
			4435 => "0000100011111000011000",
			4436 => "0001011100110000000100",
			4437 => "0000000100010110111001",
			4438 => "0001011000101000001000",
			4439 => "0000001011011000000100",
			4440 => "0000000100010110111001",
			4441 => "0000000100010110111001",
			4442 => "0001111000000000001000",
			4443 => "0000001010001000000100",
			4444 => "0000000100010110111001",
			4445 => "0000000100010110111001",
			4446 => "0000000100010110111001",
			4447 => "0000011001100000001000",
			4448 => "0010110111011100000100",
			4449 => "0000000100010110111001",
			4450 => "0000000100010110111001",
			4451 => "0001011101001000000100",
			4452 => "0000000100010110111001",
			4453 => "0001001100000000001000",
			4454 => "0011110101111100000100",
			4455 => "0000000100010110111001",
			4456 => "0000000100010110111001",
			4457 => "0001011011000000000100",
			4458 => "0000000100010110111001",
			4459 => "0011011100101000000100",
			4460 => "0000000100010110111001",
			4461 => "0000000100010110111001",
			4462 => "0011100000110100100100",
			4463 => "0001111000000000011000",
			4464 => "0001000101010100010000",
			4465 => "0000010110010000000100",
			4466 => "0000000100011001110101",
			4467 => "0000110101101100001000",
			4468 => "0000110111011100000100",
			4469 => "0000000100011001110101",
			4470 => "0000000100011001110101",
			4471 => "0000000100011001110101",
			4472 => "0001100000100000000100",
			4473 => "0000000100011001110101",
			4474 => "0000000100011001110101",
			4475 => "0010101010000100001000",
			4476 => "0010100101101100000100",
			4477 => "0000000100011001110101",
			4478 => "0000000100011001110101",
			4479 => "1111111100011001110101",
			4480 => "0010001001001100001100",
			4481 => "0000000110010100000100",
			4482 => "0000000100011001110101",
			4483 => "0000100110010100000100",
			4484 => "0000000100011001110101",
			4485 => "1111111100011001110101",
			4486 => "0000001101110100000100",
			4487 => "1111111100011001110101",
			4488 => "0011101101100000010000",
			4489 => "0001111000101000001100",
			4490 => "0000100011111000000100",
			4491 => "0000000100011001110101",
			4492 => "0011011110011000000100",
			4493 => "0000000100011001110101",
			4494 => "0000001100011001110101",
			4495 => "0000000100011001110101",
			4496 => "0010011101101000001100",
			4497 => "0010101100010000000100",
			4498 => "0000000100011001110101",
			4499 => "0010101001010100000100",
			4500 => "1111111100011001110101",
			4501 => "0000000100011001110101",
			4502 => "0010101011111000001000",
			4503 => "0010010011000000000100",
			4504 => "0000001100011001110101",
			4505 => "0000000100011001110101",
			4506 => "0001001100000000000100",
			4507 => "1111111100011001110101",
			4508 => "0000000100011001110101",
			4509 => "0010101000111000100100",
			4510 => "0001010011001000010000",
			4511 => "0000110011000000001100",
			4512 => "0001111000000100000100",
			4513 => "0000000100011101100001",
			4514 => "0000000101011000000100",
			4515 => "0000000100011101100001",
			4516 => "0000000100011101100001",
			4517 => "0000000100011101100001",
			4518 => "0000110011100100010000",
			4519 => "0000011001100000001100",
			4520 => "0001000110000000001000",
			4521 => "0001101001110000000100",
			4522 => "0000000100011101100001",
			4523 => "0000000100011101100001",
			4524 => "0000000100011101100001",
			4525 => "0000000100011101100001",
			4526 => "0000000100011101100001",
			4527 => "0010110111011100101000",
			4528 => "0000011000011000010100",
			4529 => "0000001011001000001000",
			4530 => "0011110001100000000100",
			4531 => "0000000100011101100001",
			4532 => "0000000100011101100001",
			4533 => "0010110011010000001000",
			4534 => "0000011001100100000100",
			4535 => "0000000100011101100001",
			4536 => "1111111100011101100001",
			4537 => "0000000100011101100001",
			4538 => "0010111110011000000100",
			4539 => "0000000100011101100001",
			4540 => "0011011010100100001000",
			4541 => "0001111000101000000100",
			4542 => "0000000100011101100001",
			4543 => "0000000100011101100001",
			4544 => "0001001001001000000100",
			4545 => "0000000100011101100001",
			4546 => "0000000100011101100001",
			4547 => "0010101011111000011000",
			4548 => "0001011100010000000100",
			4549 => "0000000100011101100001",
			4550 => "0011010101011100001000",
			4551 => "0001100000100000000100",
			4552 => "0000000100011101100001",
			4553 => "0000000100011101100001",
			4554 => "0011110100110100000100",
			4555 => "0000000100011101100001",
			4556 => "0011100111101000000100",
			4557 => "0000000100011101100001",
			4558 => "0000000100011101100001",
			4559 => "0011001001000100001100",
			4560 => "0010000101011100001000",
			4561 => "0000010111110000000100",
			4562 => "0000000100011101100001",
			4563 => "0000000100011101100001",
			4564 => "0000000100011101100001",
			4565 => "0010111001001000000100",
			4566 => "0000000100011101100001",
			4567 => "0000000100011101100001",
			4568 => "0000010011110001010000",
			4569 => "0001000101010100100000",
			4570 => "0010101111011000001000",
			4571 => "0001100100101000000100",
			4572 => "0000000100100000101101",
			4573 => "0000000100100000101101",
			4574 => "0000011001100000010100",
			4575 => "0001010101111000001100",
			4576 => "0011100100010000001000",
			4577 => "0010111010100100000100",
			4578 => "0000000100100000101101",
			4579 => "0000000100100000101101",
			4580 => "0000000100100000101101",
			4581 => "0011111010111100000100",
			4582 => "0000000100100000101101",
			4583 => "0000000100100000101101",
			4584 => "0000000100100000101101",
			4585 => "0000010001110000010100",
			4586 => "0010101100010000001000",
			4587 => "0000011000111100000100",
			4588 => "0000000100100000101101",
			4589 => "0000000100100000101101",
			4590 => "0011011011101100001000",
			4591 => "0010110111011100000100",
			4592 => "0000000100100000101101",
			4593 => "0000000100100000101101",
			4594 => "0000000100100000101101",
			4595 => "0011111000100100011000",
			4596 => "0011100010110000001100",
			4597 => "0000000011001100001000",
			4598 => "0011010011010000000100",
			4599 => "0000000100100000101101",
			4600 => "0000000100100000101101",
			4601 => "0000000100100000101101",
			4602 => "0010101001010100000100",
			4603 => "0000000100100000101101",
			4604 => "0001011001010000000100",
			4605 => "0000000100100000101101",
			4606 => "0000000100100000101101",
			4607 => "0000000100100000101101",
			4608 => "0001000101010100001000",
			4609 => "0001000011010000000100",
			4610 => "0000000100100000101101",
			4611 => "0000000100100000101101",
			4612 => "0000101101011000001100",
			4613 => "0000110011001000001000",
			4614 => "0000110101111000000100",
			4615 => "0000000100100000101101",
			4616 => "0000000100100000101101",
			4617 => "0000000100100000101101",
			4618 => "0000000100100000101101",
			4619 => "0011100100100100010000",
			4620 => "0010001111001000000100",
			4621 => "1111111100100011101001",
			4622 => "0010001010000100001000",
			4623 => "0000001010111100000100",
			4624 => "0000000100100011101001",
			4625 => "0000001100100011101001",
			4626 => "1111111100100011101001",
			4627 => "0000111000000000101100",
			4628 => "0011001010100100010100",
			4629 => "0010101101001000010000",
			4630 => "0011111001111000001100",
			4631 => "0000001001110100001000",
			4632 => "0000000100110100000100",
			4633 => "0000000100100011101001",
			4634 => "0000001100100011101001",
			4635 => "0000000100100011101001",
			4636 => "0000001100100011101001",
			4637 => "1111111100100011101001",
			4638 => "0000001001110100001000",
			4639 => "0001001010100100000100",
			4640 => "0000000100100011101001",
			4641 => "1111111100100011101001",
			4642 => "0011010111011100001100",
			4643 => "0000101011010000000100",
			4644 => "0000001100100011101001",
			4645 => "0001111001010100000100",
			4646 => "1111111100100011101001",
			4647 => "0000000100100011101001",
			4648 => "0000001100100011101001",
			4649 => "0010110011010000001000",
			4650 => "0000001011001000000100",
			4651 => "0000001100100011101001",
			4652 => "1111111100100011101001",
			4653 => "0001111000101000001000",
			4654 => "0001011000100000000100",
			4655 => "0000001100100011101001",
			4656 => "1111111100100011101001",
			4657 => "0010000101101100000100",
			4658 => "0000001100100011101001",
			4659 => "0010111100101000001000",
			4660 => "0010010101111000000100",
			4661 => "1111111100100011101001",
			4662 => "0000000100100011101001",
			4663 => "0010010011001000000100",
			4664 => "0000001100100011101001",
			4665 => "1111111100100011101001",
			4666 => "0011110100001100000100",
			4667 => "1111111100100101011101",
			4668 => "0000011101000000101100",
			4669 => "0010101000100000101000",
			4670 => "0001011011000000100000",
			4671 => "0000111000000000010000",
			4672 => "0011001010100100001000",
			4673 => "0010101101001000000100",
			4674 => "0000001100100101011101",
			4675 => "1111111100100101011101",
			4676 => "0000001001110100000100",
			4677 => "1111111100100101011101",
			4678 => "0000000100100101011101",
			4679 => "0011000101010100001000",
			4680 => "0000001101110100000100",
			4681 => "0000000100100101011101",
			4682 => "1111111100100101011101",
			4683 => "0000011001100000000100",
			4684 => "0000000100100101011101",
			4685 => "0000000100100101011101",
			4686 => "0011000101010100000100",
			4687 => "1111111100100101011101",
			4688 => "0000001100100101011101",
			4689 => "1111111100100101011101",
			4690 => "0011001001001000000100",
			4691 => "1111111100100101011101",
			4692 => "0010010011001000000100",
			4693 => "0000000100100101011101",
			4694 => "1111111100100101011101",
			4695 => "0011010111011101001100",
			4696 => "0010101111011000001100",
			4697 => "0001111000000100000100",
			4698 => "0000000100101000101001",
			4699 => "0000000101011000000100",
			4700 => "0000000100101000101001",
			4701 => "0000000100101000101001",
			4702 => "0011000101011100110100",
			4703 => "0010001111111100011100",
			4704 => "0000111000000000010000",
			4705 => "0010010101011100001000",
			4706 => "0000001011100000000100",
			4707 => "0000000100101000101001",
			4708 => "0000000100101000101001",
			4709 => "0011010110110100000100",
			4710 => "0000000100101000101001",
			4711 => "0000000100101000101001",
			4712 => "0010110111011100000100",
			4713 => "0000000100101000101001",
			4714 => "0001111100110000000100",
			4715 => "0000000100101000101001",
			4716 => "0000000100101000101001",
			4717 => "0000000110111100001100",
			4718 => "0001011000000000000100",
			4719 => "0000000100101000101001",
			4720 => "0001111000101000000100",
			4721 => "0000000100101000101001",
			4722 => "0000000100101000101001",
			4723 => "0011110100110100000100",
			4724 => "0000000100101000101001",
			4725 => "0001101100111100000100",
			4726 => "0000000100101000101001",
			4727 => "0000000100101000101001",
			4728 => "0001011000101000000100",
			4729 => "0000000100101000101001",
			4730 => "0001001000000000000100",
			4731 => "0000000100101000101001",
			4732 => "0000000100101000101001",
			4733 => "0000011111011100010000",
			4734 => "0000001000010000001100",
			4735 => "0001110110101100001000",
			4736 => "0001111100110000000100",
			4737 => "0000000100101000101001",
			4738 => "0000000100101000101001",
			4739 => "0000000100101000101001",
			4740 => "0000000100101000101001",
			4741 => "0000110011001000001000",
			4742 => "0010010101111000000100",
			4743 => "0000000100101000101001",
			4744 => "0000000100101000101001",
			4745 => "0000000100101000101001",
			4746 => "0001001001010000110000",
			4747 => "0000001010111100000100",
			4748 => "1111111100101010001101",
			4749 => "0000010110110100101000",
			4750 => "0010110101011100011100",
			4751 => "0001101110100000001100",
			4752 => "0001111100110000001000",
			4753 => "0001001001000100000100",
			4754 => "0000000100101010001101",
			4755 => "0000001100101010001101",
			4756 => "1111111100101010001101",
			4757 => "0000110011000000001000",
			4758 => "0000001111101100000100",
			4759 => "0000001100101010001101",
			4760 => "0000000100101010001101",
			4761 => "0010010101011100000100",
			4762 => "1111111100101010001101",
			4763 => "0000000100101010001101",
			4764 => "0010101011000000001000",
			4765 => "0011110000001000000100",
			4766 => "0000000100101010001101",
			4767 => "0000001100101010001101",
			4768 => "0000000100101010001101",
			4769 => "1111111100101010001101",
			4770 => "1111111100101010001101",
			4771 => "0001000011000001011100",
			4772 => "0001001001000100111000",
			4773 => "0011010111011100101000",
			4774 => "0011001010100100010100",
			4775 => "0000011001100000010000",
			4776 => "0010010101011100001000",
			4777 => "0000001011010000000100",
			4778 => "0000000100101101101001",
			4779 => "1111111100101101101001",
			4780 => "0010000101101100000100",
			4781 => "0000001100101101101001",
			4782 => "0000000100101101101001",
			4783 => "1111111100101101101001",
			4784 => "0001111100101100010000",
			4785 => "0000110011000000001000",
			4786 => "0011100000110100000100",
			4787 => "0000000100101101101001",
			4788 => "0000001100101101101001",
			4789 => "0000011001100000000100",
			4790 => "1111111100101101101001",
			4791 => "0000000100101101101001",
			4792 => "0000000100101101101001",
			4793 => "0011010101010100001000",
			4794 => "0010001001000100000100",
			4795 => "0000000100101101101001",
			4796 => "0000001100101101101001",
			4797 => "0011001001001000000100",
			4798 => "0000000100101101101001",
			4799 => "0000000100101101101001",
			4800 => "0000101010010100011100",
			4801 => "0010110111011100010000",
			4802 => "0010011001000100001100",
			4803 => "0010101000111000000100",
			4804 => "0000001100101101101001",
			4805 => "0010001001001100000100",
			4806 => "1111111100101101101001",
			4807 => "0000000100101101101001",
			4808 => "1111111100101101101001",
			4809 => "0001110100101100001000",
			4810 => "0010011010000100000100",
			4811 => "0000001100101101101001",
			4812 => "0000000100101101101001",
			4813 => "0000000100101101101001",
			4814 => "0010111001001000000100",
			4815 => "1111111100101101101001",
			4816 => "0000000100101101101001",
			4817 => "0010010110000000000100",
			4818 => "1111111100101101101001",
			4819 => "0010001001000100001000",
			4820 => "0011100010011000000100",
			4821 => "1111111100101101101001",
			4822 => "0000001100101101101001",
			4823 => "0000000010100000000100",
			4824 => "1111111100101101101001",
			4825 => "0000001100101101101001",
			4826 => "0000010011110001100000",
			4827 => "0011011110011000111000",
			4828 => "0000010110010000011100",
			4829 => "0010101111011000001100",
			4830 => "0011100000110100001000",
			4831 => "0001000101010100000100",
			4832 => "0000000100110001010101",
			4833 => "0000000100110001010101",
			4834 => "0000000100110001010101",
			4835 => "0010110111011100001100",
			4836 => "0000101110011100001000",
			4837 => "0000000100110100000100",
			4838 => "0000000100110001010101",
			4839 => "0000000100110001010101",
			4840 => "0000000100110001010101",
			4841 => "0000000100110001010101",
			4842 => "0011100100111000011000",
			4843 => "0001011100010000001100",
			4844 => "0010110011010000001000",
			4845 => "0010010101011100000100",
			4846 => "0000000100110001010101",
			4847 => "0000000100110001010101",
			4848 => "0000000100110001010101",
			4849 => "0000000100010100001000",
			4850 => "0010110011010000000100",
			4851 => "0000000100110001010101",
			4852 => "0000000100110001010101",
			4853 => "0000000100110001010101",
			4854 => "0000000100110001010101",
			4855 => "0000010111100100010000",
			4856 => "0001100001100000001100",
			4857 => "0000001011001000001000",
			4858 => "0000000000011100000100",
			4859 => "0000000100110001010101",
			4860 => "0000000100110001010101",
			4861 => "0000000100110001010101",
			4862 => "0000000100110001010101",
			4863 => "0001001010000100001000",
			4864 => "0010000101101100000100",
			4865 => "0000000100110001010101",
			4866 => "0000000100110001010101",
			4867 => "0000011000011000000100",
			4868 => "0000000100110001010101",
			4869 => "0011100011101100001000",
			4870 => "0001111000101000000100",
			4871 => "0000000100110001010101",
			4872 => "0000000100110001010101",
			4873 => "0000000100110001010101",
			4874 => "0000101101011000010100",
			4875 => "0001000101010100001000",
			4876 => "0001000011010000000100",
			4877 => "0000000100110001010101",
			4878 => "0000000100110001010101",
			4879 => "0000110011001000001000",
			4880 => "0000111111011000000100",
			4881 => "0000000100110001010101",
			4882 => "0000000100110001010101",
			4883 => "0000000100110001010101",
			4884 => "0000000100110001010101",
			4885 => "0011110111100000010100",
			4886 => "0010010110000000010000",
			4887 => "0011001100101000001100",
			4888 => "0011010110001100001000",
			4889 => "0000011000011000000100",
			4890 => "1111111100110100011001",
			4891 => "0000001100110100011001",
			4892 => "1111111100110100011001",
			4893 => "0000001100110100011001",
			4894 => "1111111100110100011001",
			4895 => "0000111000000000101000",
			4896 => "0010110101011100100100",
			4897 => "0011001010100100010000",
			4898 => "0011000110001100000100",
			4899 => "0000000100110100011001",
			4900 => "0010101101001000001000",
			4901 => "0001000101010100000100",
			4902 => "0000001100110100011001",
			4903 => "0000001100110100011001",
			4904 => "1111111100110100011001",
			4905 => "0000001001110100001000",
			4906 => "0001000111011100000100",
			4907 => "0000000100110100011001",
			4908 => "1111111100110100011001",
			4909 => "0010001001001100000100",
			4910 => "0000000100110100011001",
			4911 => "0011111001111000000100",
			4912 => "0000001100110100011001",
			4913 => "0000000100110100011001",
			4914 => "0000001100110100011001",
			4915 => "0001010110101100000100",
			4916 => "1111111100110100011001",
			4917 => "0010001111001000011000",
			4918 => "0001000011000000001100",
			4919 => "0010001001001100000100",
			4920 => "1111111100110100011001",
			4921 => "0011111011110100000100",
			4922 => "0000001100110100011001",
			4923 => "0000001100110100011001",
			4924 => "0010010110000000000100",
			4925 => "1111111100110100011001",
			4926 => "0001111011111000000100",
			4927 => "0000001100110100011001",
			4928 => "0000000100110100011001",
			4929 => "0011001001000100000100",
			4930 => "1111111100110100011001",
			4931 => "0010000011001000000100",
			4932 => "0000001100110100011001",
			4933 => "1111111100110100011001",
			4934 => "0001000110000001001000",
			4935 => "0011010111011100111100",
			4936 => "0011011011101100100100",
			4937 => "0001010011001000010100",
			4938 => "0000110011000000001100",
			4939 => "0001111000000100000100",
			4940 => "0000000100110111111101",
			4941 => "0000001100010100000100",
			4942 => "0000000100110111111101",
			4943 => "0000001100110111111101",
			4944 => "0001011010000100000100",
			4945 => "0000000100110111111101",
			4946 => "1111111100110111111101",
			4947 => "0000111000000000001100",
			4948 => "0001000101010100000100",
			4949 => "0000000100110111111101",
			4950 => "0011001010100100000100",
			4951 => "0000001100110111111101",
			4952 => "0000000100110111111101",
			4953 => "0000000100110111111101",
			4954 => "0001110110101100001100",
			4955 => "0000011001100000001000",
			4956 => "0011000011010000000100",
			4957 => "0000000100110111111101",
			4958 => "0000000100110111111101",
			4959 => "1111111100110111111101",
			4960 => "0010101111101000001000",
			4961 => "0010101000111000000100",
			4962 => "0000000100110111111101",
			4963 => "1111111100110111111101",
			4964 => "0000000100110111111101",
			4965 => "0001011101001000001000",
			4966 => "0000000111101100000100",
			4967 => "0000000100110111111101",
			4968 => "0000001100110111111101",
			4969 => "0000000100110111111101",
			4970 => "0001011100110000000100",
			4971 => "1111111100110111111101",
			4972 => "0001011000101000010000",
			4973 => "0001000011000000001100",
			4974 => "0011111001111000001000",
			4975 => "0001001010000100000100",
			4976 => "0000000100110111111101",
			4977 => "0000001100110111111101",
			4978 => "0000000100110111111101",
			4979 => "0000000100110111111101",
			4980 => "0000111100110000000100",
			4981 => "1111111100110111111101",
			4982 => "0010011001000100000100",
			4983 => "1111111100110111111101",
			4984 => "0011011010100100001000",
			4985 => "0001010001001000000100",
			4986 => "0000001100110111111101",
			4987 => "0000000100110111111101",
			4988 => "0011001001000100000100",
			4989 => "0000000100110111111101",
			4990 => "0000000100110111111101",
			4991 => "0011111011011100111000",
			4992 => "0001111001010100110100",
			4993 => "0001111101001000101000",
			4994 => "0000111100010000011100",
			4995 => "0001011000000000010000",
			4996 => "0001111000111000001000",
			4997 => "0011001010100100000100",
			4998 => "0000000100111011010001",
			4999 => "1111111100111011010001",
			5000 => "0000111001000100000100",
			5001 => "0000000100111011010001",
			5002 => "1111111100111011010001",
			5003 => "0010011001000100001000",
			5004 => "0000000100011000000100",
			5005 => "0000000100111011010001",
			5006 => "0000001100111011010001",
			5007 => "1111111100111011010001",
			5008 => "0000011001100000000100",
			5009 => "1111111100111011010001",
			5010 => "0000001010111100000100",
			5011 => "0000000100111011010001",
			5012 => "0000000100111011010001",
			5013 => "0000011000011000000100",
			5014 => "0000000100111011010001",
			5015 => "0010000000110000000100",
			5016 => "0000001100111011010001",
			5017 => "0000000100111011010001",
			5018 => "1111111100111011010001",
			5019 => "0011010101011100101000",
			5020 => "0011010111011100100000",
			5021 => "0001011011000000011100",
			5022 => "0010000101011100001100",
			5023 => "0000101010010100001000",
			5024 => "0001011101001000000100",
			5025 => "0000001100111011010001",
			5026 => "1111111100111011010001",
			5027 => "1111111100111011010001",
			5028 => "0001000111011100001000",
			5029 => "0001010101111000000100",
			5030 => "0000000100111011010001",
			5031 => "1111111100111011010001",
			5032 => "0000000110111100000100",
			5033 => "0000000100111011010001",
			5034 => "0000000100111011010001",
			5035 => "0000001100111011010001",
			5036 => "0001011000101000000100",
			5037 => "0000001100111011010001",
			5038 => "0000000100111011010001",
			5039 => "0011111110011100000100",
			5040 => "1111111100111011010001",
			5041 => "0001101101001100000100",
			5042 => "0000000100111011010001",
			5043 => "0000000100111011010001",
			5044 => "0011011110011000110000",
			5045 => "0010101000000000010000",
			5046 => "0001111111011000000100",
			5047 => "0000000100111110111101",
			5048 => "0000000100011000000100",
			5049 => "0000000100111110111101",
			5050 => "0010101111011000000100",
			5051 => "0000000100111110111101",
			5052 => "0000000100111110111101",
			5053 => "0000010001100100011100",
			5054 => "0010010101101100010100",
			5055 => "0010111110011000010000",
			5056 => "0001101101010000001000",
			5057 => "0011100110100000000100",
			5058 => "0000000100111110111101",
			5059 => "0000000100111110111101",
			5060 => "0000000101101000000100",
			5061 => "0000000100111110111101",
			5062 => "0000000100111110111101",
			5063 => "0000000100111110111101",
			5064 => "0000111000000000000100",
			5065 => "0000000100111110111101",
			5066 => "0000000100111110111101",
			5067 => "0000000100111110111101",
			5068 => "0010011001001000001000",
			5069 => "0010101101001000000100",
			5070 => "0000000100111110111101",
			5071 => "0000000100111110111101",
			5072 => "0010110011010000010000",
			5073 => "0001011000000000000100",
			5074 => "0000000100111110111101",
			5075 => "0011011010100100001000",
			5076 => "0010101000101000000100",
			5077 => "0000000100111110111101",
			5078 => "0000000100111110111101",
			5079 => "0000000100111110111101",
			5080 => "0011101101100000010100",
			5081 => "0001111000101000001100",
			5082 => "0001010011000100001000",
			5083 => "0011111110000000000100",
			5084 => "0000000100111110111101",
			5085 => "0000000100111110111101",
			5086 => "0000000100111110111101",
			5087 => "0000110011001000000100",
			5088 => "0000000100111110111101",
			5089 => "0000000100111110111101",
			5090 => "0001011011000000010000",
			5091 => "0010110101011100001000",
			5092 => "0010110111011100000100",
			5093 => "0000000100111110111101",
			5094 => "0000000100111110111101",
			5095 => "0000101111001100000100",
			5096 => "0000000100111110111101",
			5097 => "0000000100111110111101",
			5098 => "0000101011100100000100",
			5099 => "0000000100111110111101",
			5100 => "0000101111001100000100",
			5101 => "0000000100111110111101",
			5102 => "0000000100111110111101",
			5103 => "0001111111011000000100",
			5104 => "1111111101000001011001",
			5105 => "0000110011000000001000",
			5106 => "0000000101011000000100",
			5107 => "0000000101000001011001",
			5108 => "0000001101000001011001",
			5109 => "0010110011010000011100",
			5110 => "0001000011000000011000",
			5111 => "0011111010101100001000",
			5112 => "0001001001000100000100",
			5113 => "0000000101000001011001",
			5114 => "0000000101000001011001",
			5115 => "0011110000001000001000",
			5116 => "0011110010000100000100",
			5117 => "0000000101000001011001",
			5118 => "1111111101000001011001",
			5119 => "0000001101110000000100",
			5120 => "0000001101000001011001",
			5121 => "0000000101000001011001",
			5122 => "1111111101000001011001",
			5123 => "0000010111100100001100",
			5124 => "0001011100110000000100",
			5125 => "0000000101000001011001",
			5126 => "0000001100001000000100",
			5127 => "0000000101000001011001",
			5128 => "0000001101000001011001",
			5129 => "0001111000101000001100",
			5130 => "0011011110011000000100",
			5131 => "0000000101000001011001",
			5132 => "0000011000011000000100",
			5133 => "0000000101000001011001",
			5134 => "0000001101000001011001",
			5135 => "0011100001000000001000",
			5136 => "0001011100010000000100",
			5137 => "0000000101000001011001",
			5138 => "1111111101000001011001",
			5139 => "0011100111100000000100",
			5140 => "0000001101000001011001",
			5141 => "0000000101000001011001",
			5142 => "0001111111011000000100",
			5143 => "0000000101000100100111",
			5144 => "0010101000111000100000",
			5145 => "0001000110000000011100",
			5146 => "0001001001000100011000",
			5147 => "0011000011010000001100",
			5148 => "0011111110101100001000",
			5149 => "0010010101011100000100",
			5150 => "0000000101000100100111",
			5151 => "0000000101000100100111",
			5152 => "0000001101000100100111",
			5153 => "0000110011000000001000",
			5154 => "0001010110000000000100",
			5155 => "0000000101000100100111",
			5156 => "0000000101000100100111",
			5157 => "1111111101000100100111",
			5158 => "0000001101000100100111",
			5159 => "0000000101000100100111",
			5160 => "0001011100110000010100",
			5161 => "0011111100111100000100",
			5162 => "1111111101000100100111",
			5163 => "0000010110010000001000",
			5164 => "0010111011101100000100",
			5165 => "0000000101000100100111",
			5166 => "1111111101000100100111",
			5167 => "0001101110000100000100",
			5168 => "0000000101000100100111",
			5169 => "0000000101000100100111",
			5170 => "0010101011111000011100",
			5171 => "0001011011111000010000",
			5172 => "0001000011000000001000",
			5173 => "0011111001111000000100",
			5174 => "0000000101000100100111",
			5175 => "0000000101000100100111",
			5176 => "0010110101011100000100",
			5177 => "1111111101000100100111",
			5178 => "0000000101000100100111",
			5179 => "0011010101010100001000",
			5180 => "0011000101010100000100",
			5181 => "0000000101000100100111",
			5182 => "0000001101000100100111",
			5183 => "0000000101000100100111",
			5184 => "0011001001000100001100",
			5185 => "0001110100101100001000",
			5186 => "0001111001010000000100",
			5187 => "0000000101000100100111",
			5188 => "0000000101000100100111",
			5189 => "1111111101000100100111",
			5190 => "0010011000000100000100",
			5191 => "0000001101000100100111",
			5192 => "0000000101000100100111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1797, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3471, initial_addr_3'length));
	end generate gen_rom_4;

	gen_rom_5: if SELECT_ROM = 5 generate
		bank <= (
			0 => "0001101010001000010000",
			1 => "0011110010110000000100",
			2 => "1111111000000010000101",
			3 => "0000001000100100001000",
			4 => "0001011000000000000100",
			5 => "1111111000000010000101",
			6 => "0000001000000010000101",
			7 => "1111111000000010000101",
			8 => "0000011001100000010000",
			9 => "0011100011101000001000",
			10 => "0001111100010000000100",
			11 => "0000000000000010000101",
			12 => "1111111000000010000101",
			13 => "0000000101101000000100",
			14 => "1111111000000010000101",
			15 => "0000000000000010000101",
			16 => "0001011000100000011000",
			17 => "0001111110001100010100",
			18 => "0000001010111000001100",
			19 => "0011110010000100000100",
			20 => "0000001000000010000101",
			21 => "0010001111001000000100",
			22 => "1111111000000010000101",
			23 => "0000001000000010000101",
			24 => "0010000011001000000100",
			25 => "0000001000000010000101",
			26 => "0000001000000010000101",
			27 => "1111111000000010000101",
			28 => "0010101100001100001000",
			29 => "0001111001011000000100",
			30 => "0000000000000010000101",
			31 => "1111111000000010000101",
			32 => "0000001000000010000101",
			33 => "0000000110101000011000",
			34 => "0011110010110000000100",
			35 => "1111111000000100000001",
			36 => "0001111000101000001000",
			37 => "0010001001000100000100",
			38 => "1111111000000100000001",
			39 => "0000010000000100000001",
			40 => "0000010011010000000100",
			41 => "1111111000000100000001",
			42 => "0000000010101100000100",
			43 => "0000000000000100000001",
			44 => "1111111000000100000001",
			45 => "0010000101101100000100",
			46 => "1111111000000100000001",
			47 => "0011010011000000011100",
			48 => "0010101010011100011000",
			49 => "0001011000100000010000",
			50 => "0001100001111000001000",
			51 => "0001100111101000000100",
			52 => "0000001000000100000001",
			53 => "1111111000000100000001",
			54 => "0011111011110100000100",
			55 => "0000010000000100000001",
			56 => "0000001000000100000001",
			57 => "0001111000100000000100",
			58 => "0000001000000100000001",
			59 => "1111111000000100000001",
			60 => "0000010000000100000001",
			61 => "0000010101010100000100",
			62 => "0000000000000100000001",
			63 => "1111111000000100000001",
			64 => "0011111010101100001100",
			65 => "0011110010110000000100",
			66 => "1111111000000101110101",
			67 => "0011100000010100000100",
			68 => "0000000000000101110101",
			69 => "1111111000000101110101",
			70 => "0000010111100100000100",
			71 => "1111111000000101110101",
			72 => "0001110011110100100100",
			73 => "0000100000000000010100",
			74 => "0000010011110000001000",
			75 => "0000000111110100000100",
			76 => "0000000000000101110101",
			77 => "1111111000000101110101",
			78 => "0001111111101000000100",
			79 => "0000010000000101110101",
			80 => "0000110011000100000100",
			81 => "0000000000000101110101",
			82 => "0000010000000101110101",
			83 => "0011111011010100000100",
			84 => "0000010000000101110101",
			85 => "0011100100111000000100",
			86 => "0000000000000101110101",
			87 => "0001110001011000000100",
			88 => "0000001000000101110101",
			89 => "0000001000000101110101",
			90 => "0001011011000000000100",
			91 => "0000000000000101110101",
			92 => "1111111000000101110101",
			93 => "0000100100010100110100",
			94 => "0011001100101000100000",
			95 => "0001000101111000010000",
			96 => "0001110001010000001100",
			97 => "0000011001100000000100",
			98 => "0000000000001001000001",
			99 => "0000001101001100000100",
			100 => "0000000000001001000001",
			101 => "0000000000001001000001",
			102 => "0000000000001001000001",
			103 => "0001101111110000000100",
			104 => "0000000000001001000001",
			105 => "0000111011111000001000",
			106 => "0010000101101100000100",
			107 => "0000000000001001000001",
			108 => "0000000000001001000001",
			109 => "0000000000001001000001",
			110 => "0000011100101000001100",
			111 => "0000111110001100000100",
			112 => "1111111000001001000001",
			113 => "0010111001001000000100",
			114 => "0000000000001001000001",
			115 => "0000000000001001000001",
			116 => "0011100110111000000100",
			117 => "0000000000001001000001",
			118 => "0000000000001001000001",
			119 => "0000010101011100101000",
			120 => "0000011101000000010000",
			121 => "0010110111011100001100",
			122 => "0000010111100100000100",
			123 => "0000000000001001000001",
			124 => "0010000101101100000100",
			125 => "0000000000001001000001",
			126 => "0000000000001001000001",
			127 => "0000000000001001000001",
			128 => "0001110011110100010000",
			129 => "0000111101001000000100",
			130 => "0000000000001001000001",
			131 => "0001010110011100000100",
			132 => "0000000000001001000001",
			133 => "0001011000100000000100",
			134 => "0000000000001001000001",
			135 => "0000000000001001000001",
			136 => "0001000110101100000100",
			137 => "0000000000001001000001",
			138 => "0000000000001001000001",
			139 => "0000011100101000000100",
			140 => "0000000000001001000001",
			141 => "0011110011111100000100",
			142 => "0000000000001001000001",
			143 => "0000000000001001000001",
			144 => "0011110000001100010100",
			145 => "0011110010110000000100",
			146 => "1111111000001011100101",
			147 => "0011100000010100000100",
			148 => "0000001000001011100101",
			149 => "0000100010101000001000",
			150 => "0000001001111000000100",
			151 => "1111111000001011100101",
			152 => "0000001000001011100101",
			153 => "1111111000001011100101",
			154 => "0011011101101000110100",
			155 => "0000011001100000010000",
			156 => "0000001010111000001000",
			157 => "0001111100101100000100",
			158 => "1111111000001011100101",
			159 => "0000000000001011100101",
			160 => "0010111110011000000100",
			161 => "0000010000001011100101",
			162 => "0000000000001011100101",
			163 => "0000001010111000011000",
			164 => "0011100110111000010000",
			165 => "0000011101000000001000",
			166 => "0011100110110000000100",
			167 => "0000000000001011100101",
			168 => "0000010000001011100101",
			169 => "0010111001001000000100",
			170 => "0000011000001011100101",
			171 => "0000000000001011100101",
			172 => "0000000101101000000100",
			173 => "1111111000001011100101",
			174 => "0000001000001011100101",
			175 => "0001011000100000001000",
			176 => "0011111110011100000100",
			177 => "0000011000001011100101",
			178 => "0000010000001011100101",
			179 => "0000001000001011100101",
			180 => "0000010111011100001000",
			181 => "0011011010000100000100",
			182 => "1111111000001011100101",
			183 => "0000010000001011100101",
			184 => "1111111000001011100101",
			185 => "0011110100010000001100",
			186 => "0010111011101100001000",
			187 => "0001001001000100000100",
			188 => "1111111000001101101001",
			189 => "0000010000001101101001",
			190 => "1111111000001101101001",
			191 => "0000010111100100000100",
			192 => "1111111000001101101001",
			193 => "0010110111011100011000",
			194 => "0001010011001000001000",
			195 => "0010101100010000000100",
			196 => "0000000000001101101001",
			197 => "1111111000001101101001",
			198 => "0001101110010000000100",
			199 => "0000001000001101101001",
			200 => "0000100011111000000100",
			201 => "1111111000001101101001",
			202 => "0010000101101100000100",
			203 => "1111111000001101101001",
			204 => "0000001000001101101001",
			205 => "0011010101010100001100",
			206 => "0010101001000000001000",
			207 => "0001001000000100000100",
			208 => "1111111000001101101001",
			209 => "1111111000001101101001",
			210 => "0000001000001101101001",
			211 => "0011111101010000000100",
			212 => "1111111000001101101001",
			213 => "0011010101111000001000",
			214 => "0000011100101000000100",
			215 => "0000000000001101101001",
			216 => "0000001000001101101001",
			217 => "1111111000001101101001",
			218 => "0000100000000000110100",
			219 => "0011111010101100010100",
			220 => "0011110010110000000100",
			221 => "1111111000010000011101",
			222 => "0011100000010100000100",
			223 => "0000010000010000011101",
			224 => "0010101100010000001000",
			225 => "0000001000001000000100",
			226 => "1111111000010000011101",
			227 => "0000001000010000011101",
			228 => "1111111000010000011101",
			229 => "0000011001100000000100",
			230 => "1111111000010000011101",
			231 => "0010000011100100010000",
			232 => "0001101000110100000100",
			233 => "0000101000010000011101",
			234 => "0000001000010000000100",
			235 => "1111111000010000011101",
			236 => "0000101111101100000100",
			237 => "0000100000010000011101",
			238 => "0000001000010000011101",
			239 => "0001011011000000000100",
			240 => "0000001000010000011101",
			241 => "0001011110010100000100",
			242 => "1111111000010000011101",
			243 => "0000000000010000011101",
			244 => "0001110011110100100000",
			245 => "0000011001100000001000",
			246 => "0000010111100100000100",
			247 => "1111111000010000011101",
			248 => "0000001000010000011101",
			249 => "0001110001011000010000",
			250 => "0010001111001000000100",
			251 => "0000010000010000011101",
			252 => "0000111000101000001000",
			253 => "0000111101001000000100",
			254 => "0000100000010000011101",
			255 => "0000011000010000011101",
			256 => "0000101000010000011101",
			257 => "0001010011000100000100",
			258 => "0000011000010000011101",
			259 => "0000000000010000011101",
			260 => "0000111001010000000100",
			261 => "0000001000010000011101",
			262 => "1111111000010000011101",
			263 => "0011010011000000110000",
			264 => "0010001111111100000100",
			265 => "1111111000010010000001",
			266 => "0011011010000100011100",
			267 => "0011010110000000011000",
			268 => "0001111110111000010000",
			269 => "0011011100101000001000",
			270 => "0010110101010100000100",
			271 => "0000000000010010000001",
			272 => "0000000000010010000001",
			273 => "0000101101111000000100",
			274 => "0000000000010010000001",
			275 => "0000001000010010000001",
			276 => "0000011110011000000100",
			277 => "0000000000010010000001",
			278 => "1111111000010010000001",
			279 => "1111111000010010000001",
			280 => "0000111111101000001000",
			281 => "0001011101101000000100",
			282 => "0000000000010010000001",
			283 => "0000001000010010000001",
			284 => "0010101110010100000100",
			285 => "1111111000010010000001",
			286 => "0000001000010010000001",
			287 => "1111111000010010000001",
			288 => "0000100100010100111000",
			289 => "0011001100101000100100",
			290 => "0001000101111000010000",
			291 => "0001110001010000001100",
			292 => "0000011001100000000100",
			293 => "0000000000010101011101",
			294 => "0000001101001100000100",
			295 => "0000000000010101011101",
			296 => "0000000000010101011101",
			297 => "0000000000010101011101",
			298 => "0010011101101000001100",
			299 => "0000001100111100001000",
			300 => "0000000000010000000100",
			301 => "0000000000010101011101",
			302 => "0000000000010101011101",
			303 => "0000000000010101011101",
			304 => "0001100001101100000100",
			305 => "0000000000010101011101",
			306 => "0000000000010101011101",
			307 => "0000011100101000001100",
			308 => "0000111110001100000100",
			309 => "1111111000010101011101",
			310 => "0010111001001000000100",
			311 => "0000000000010101011101",
			312 => "0000000000010101011101",
			313 => "0011100110111000000100",
			314 => "0000000000010101011101",
			315 => "0000000000010101011101",
			316 => "0000010101011100101100",
			317 => "0010001010000100010100",
			318 => "0000111000000000001000",
			319 => "0010001111111100000100",
			320 => "0000000000010101011101",
			321 => "0000000000010101011101",
			322 => "0001010110011100001000",
			323 => "0011100101000000000100",
			324 => "0000000000010101011101",
			325 => "0000000000010101011101",
			326 => "0000000000010101011101",
			327 => "0001000011000000000100",
			328 => "0000000000010101011101",
			329 => "0010001100110000010000",
			330 => "0010111001001000001000",
			331 => "0010001111011000000100",
			332 => "0000000000010101011101",
			333 => "0000000000010101011101",
			334 => "0000100111111000000100",
			335 => "0000000000010101011101",
			336 => "0000000000010101011101",
			337 => "0000000000010101011101",
			338 => "0000011100101000000100",
			339 => "0000000000010101011101",
			340 => "0011110011111100000100",
			341 => "0000000000010101011101",
			342 => "0000000000010101011101",
			343 => "0011110100010000001100",
			344 => "0011000011010000001000",
			345 => "0000011101000000000100",
			346 => "1111111000010111010001",
			347 => "0000001000010111010001",
			348 => "1111111000010111010001",
			349 => "0000010111100100000100",
			350 => "1111111000010111010001",
			351 => "0001111100110000000100",
			352 => "0000001000010111010001",
			353 => "0011100100101000010100",
			354 => "0010011100000000010000",
			355 => "0000011101000000001000",
			356 => "0001100110000100000100",
			357 => "0000001000010111010001",
			358 => "1111111000010111010001",
			359 => "0001000110000000000100",
			360 => "0000000000010111010001",
			361 => "0000001000010111010001",
			362 => "1111111000010111010001",
			363 => "0011100101100000001100",
			364 => "0000001101011100000100",
			365 => "1111111000010111010001",
			366 => "0000001100100100000100",
			367 => "0000010000010111010001",
			368 => "0000001000010111010001",
			369 => "0000111001010000000100",
			370 => "0000000000010111010001",
			371 => "1111111000010111010001",
			372 => "0011010011000000110100",
			373 => "0011100101100000101100",
			374 => "0011111011011000100000",
			375 => "0001000101010100000100",
			376 => "1111111000011000111101",
			377 => "0000010110001100010000",
			378 => "0001011100101100001000",
			379 => "0010000000110000000100",
			380 => "0000000000011000111101",
			381 => "0000000000011000111101",
			382 => "0000101011001100000100",
			383 => "1111111000011000111101",
			384 => "0000000000011000111101",
			385 => "0001001001001000000100",
			386 => "1111111000011000111101",
			387 => "0011011001001000000100",
			388 => "0000000000011000111101",
			389 => "0000000000011000111101",
			390 => "0011001110011000000100",
			391 => "0000000000011000111101",
			392 => "0011101110010000000100",
			393 => "0000001000011000111101",
			394 => "0000000000011000111101",
			395 => "0011110110001000000100",
			396 => "1111111000011000111101",
			397 => "0000000000011000111101",
			398 => "1111111000011000111101",
			399 => "0011110100010000001100",
			400 => "0011000011010000001000",
			401 => "0000011101000000000100",
			402 => "1111111000011011000001",
			403 => "0000001000011011000001",
			404 => "1111111000011011000001",
			405 => "0000010111100100000100",
			406 => "1111111000011011000001",
			407 => "0010110011010000011100",
			408 => "0001010011001000001000",
			409 => "0011001110011000000100",
			410 => "1111111000011011000001",
			411 => "0000000000011011000001",
			412 => "0010000101101100001000",
			413 => "0011110000001000000100",
			414 => "0000001000011011000001",
			415 => "1111111000011011000001",
			416 => "0011111011010100000100",
			417 => "0000001000011011000001",
			418 => "0000001101011000000100",
			419 => "0000000000011011000001",
			420 => "0000001000011011000001",
			421 => "0000010011110000000100",
			422 => "1111111000011011000001",
			423 => "0000111010011100010000",
			424 => "0001011011000000001000",
			425 => "0001101110000100000100",
			426 => "0000000000011011000001",
			427 => "0000001000011011000001",
			428 => "0001111100011100000100",
			429 => "0000000000011011000001",
			430 => "1111111000011011000001",
			431 => "0000001000011011000001",
			432 => "0001101111110000000100",
			433 => "1111111000011100011101",
			434 => "0010010110101100101000",
			435 => "0000011100101000100000",
			436 => "0010111010000100011100",
			437 => "0010000011100100010000",
			438 => "0001001111011000001000",
			439 => "0000011001100000000100",
			440 => "1111111000011100011101",
			441 => "0000000000011100011101",
			442 => "0001111100101100000100",
			443 => "0000001000011100011101",
			444 => "0000000000011100011101",
			445 => "0000111100110000000100",
			446 => "0000000000011100011101",
			447 => "0010101001011000000100",
			448 => "1111111000011100011101",
			449 => "0000000000011100011101",
			450 => "0000001000011100011101",
			451 => "0000111011111000000100",
			452 => "0000001000011100011101",
			453 => "0000000000011100011101",
			454 => "1111111000011100011101",
			455 => "0011110010110000000100",
			456 => "1111111000011101110001",
			457 => "0010001111111100000100",
			458 => "1111111000011101110001",
			459 => "0001111100110000000100",
			460 => "0000001000011101110001",
			461 => "0010101000111000000100",
			462 => "1111111000011101110001",
			463 => "0000111100010000001100",
			464 => "0000010011010000001000",
			465 => "0011000101010100000100",
			466 => "0000001000011101110001",
			467 => "0000000000011101110001",
			468 => "0000001000011101110001",
			469 => "0001011011111000001000",
			470 => "0010111100101000000100",
			471 => "0000000000011101110001",
			472 => "1111111000011101110001",
			473 => "0000010110001100000100",
			474 => "0000000000011101110001",
			475 => "0000000000011101110001",
			476 => "0001011000000000011000",
			477 => "0001111100010000001000",
			478 => "0000110011001000000100",
			479 => "0000000000100000110101",
			480 => "0000000000100000110101",
			481 => "0000110011000000001000",
			482 => "0000111101101000000100",
			483 => "0000000000100000110101",
			484 => "0000000000100000110101",
			485 => "0011101000110100000100",
			486 => "0000000000100000110101",
			487 => "0000000000100000110101",
			488 => "0000101100001000100100",
			489 => "0011111110101100011100",
			490 => "0001011011000000011000",
			491 => "0010101001010100001100",
			492 => "0001011100010000000100",
			493 => "0000000000100000110101",
			494 => "0001011001010100000100",
			495 => "0000000000100000110101",
			496 => "0000000000100000110101",
			497 => "0010111100101000001000",
			498 => "0010000101101100000100",
			499 => "0000000000100000110101",
			500 => "0000000000100000110101",
			501 => "0000000000100000110101",
			502 => "0000000000100000110101",
			503 => "0001111111101000000100",
			504 => "0000000000100000110101",
			505 => "0000000000100000110101",
			506 => "0011000101010100001000",
			507 => "0000010111100100000100",
			508 => "0000000000100000110101",
			509 => "0000000000100000110101",
			510 => "0010010011000000001000",
			511 => "0010010110000000000100",
			512 => "0000000000100000110101",
			513 => "0000000000100000110101",
			514 => "0001011011111000001000",
			515 => "0000001010111000000100",
			516 => "0000000000100000110101",
			517 => "0000000000100000110101",
			518 => "0001010011000100001000",
			519 => "0010010110101100000100",
			520 => "0000000000100000110101",
			521 => "0000000000100000110101",
			522 => "0010101100001100000100",
			523 => "0000000000100000110101",
			524 => "0000000000100000110101",
			525 => "0000100100010101001100",
			526 => "0011000101101100111000",
			527 => "0001101010001000011100",
			528 => "0000011000011000010000",
			529 => "0010111010100100001100",
			530 => "0000110011001000000100",
			531 => "0000000000100100111001",
			532 => "0000001000100100000100",
			533 => "0000000000100100111001",
			534 => "0000000000100100111001",
			535 => "0000000000100100111001",
			536 => "0000110011000000001000",
			537 => "0000111001000100000100",
			538 => "0000000000100100111001",
			539 => "0000000000100100111001",
			540 => "0000000000100100111001",
			541 => "0001100001100000001100",
			542 => "0011111110101100001000",
			543 => "0000010111100100000100",
			544 => "0000000000100100111001",
			545 => "0000000000100100111001",
			546 => "0000000000100100111001",
			547 => "0000000100010100000100",
			548 => "0000000000100100111001",
			549 => "0001100111101000000100",
			550 => "0000000000100100111001",
			551 => "0011111011000100000100",
			552 => "0000000000100100111001",
			553 => "0000000000100100111001",
			554 => "0000011100101000001100",
			555 => "0010100111010100000100",
			556 => "0000000000100100111001",
			557 => "0001010000110100000100",
			558 => "0000000000100100111001",
			559 => "0000000000100100111001",
			560 => "0011100110111000000100",
			561 => "0000000000100100111001",
			562 => "0000000000100100111001",
			563 => "0001100100100000010100",
			564 => "0001101110001000001000",
			565 => "0000001110110000000100",
			566 => "0000000000100100111001",
			567 => "0000000000100100111001",
			568 => "0011111011010100001000",
			569 => "0000010011110000000100",
			570 => "0000000000100100111001",
			571 => "0000000000100100111001",
			572 => "0000000000100100111001",
			573 => "0000001101011000010000",
			574 => "0011010101101100001000",
			575 => "0000111000101000000100",
			576 => "0000000000100100111001",
			577 => "0000000000100100111001",
			578 => "0001010011000100000100",
			579 => "0000000000100100111001",
			580 => "0000000000100100111001",
			581 => "0000010101010100001100",
			582 => "0000101110101000001000",
			583 => "0010000000110000000100",
			584 => "0000000000100100111001",
			585 => "0000000000100100111001",
			586 => "0000000000100100111001",
			587 => "0000011100101000000100",
			588 => "0000000000100100111001",
			589 => "0000000000100100111001",
			590 => "0010011000000101000000",
			591 => "0011001001001000101100",
			592 => "0011011100101000101000",
			593 => "0010110101010100011100",
			594 => "0000010011110000001100",
			595 => "0010111010100100001000",
			596 => "0010000101101100000100",
			597 => "1111111000101000010101",
			598 => "0000000000101000010101",
			599 => "1111111000101000010101",
			600 => "0011101110100100001000",
			601 => "0000001101001100000100",
			602 => "1111111000101000010101",
			603 => "0000001000101000010101",
			604 => "0000111001010100000100",
			605 => "1111111000101000010101",
			606 => "0000000000101000010101",
			607 => "0010101001011000000100",
			608 => "1111111000101000010101",
			609 => "0010010011000000000100",
			610 => "0000000000101000010101",
			611 => "0000000000101000010101",
			612 => "0000001000101000010101",
			613 => "0010100000111100001000",
			614 => "0000101011001100000100",
			615 => "1111111000101000010101",
			616 => "0000000000101000010101",
			617 => "0011000101101100001000",
			618 => "0010010101111000000100",
			619 => "0000000000101000010101",
			620 => "0000001000101000010101",
			621 => "0000000000101000010101",
			622 => "0001010011000100100000",
			623 => "0000111000000000001100",
			624 => "0011011001001000001000",
			625 => "0011011100101000000100",
			626 => "0000000000101000010101",
			627 => "0000000000101000010101",
			628 => "1111111000101000010101",
			629 => "0010010110101100010000",
			630 => "0011101111010100000100",
			631 => "1111111000101000010101",
			632 => "0001011011111000000100",
			633 => "0000000000101000010101",
			634 => "0000010111011100000100",
			635 => "0000001000101000010101",
			636 => "0000000000101000010101",
			637 => "1111111000101000010101",
			638 => "0000110000111000001000",
			639 => "0010000011001000000100",
			640 => "0000000000101000010101",
			641 => "1111111000101000010101",
			642 => "0001001110010100000100",
			643 => "0000001000101000010101",
			644 => "0000000000101000010101",
			645 => "0010110101010100111000",
			646 => "0000101100001000100000",
			647 => "0011100001000100011100",
			648 => "0011100011010100010000",
			649 => "0011110011101100001000",
			650 => "0001101100100000000100",
			651 => "0000000000101100000001",
			652 => "0000000000101100000001",
			653 => "0001001100000000000100",
			654 => "0000000000101100000001",
			655 => "0000000000101100000001",
			656 => "0000100010101100001000",
			657 => "0000011000011000000100",
			658 => "0000000000101100000001",
			659 => "0000000000101100000001",
			660 => "0000000000101100000001",
			661 => "0000000000101100000001",
			662 => "0000010111100100000100",
			663 => "0000000000101100000001",
			664 => "0011100100101000001100",
			665 => "0001100101100000000100",
			666 => "0000000000101100000001",
			667 => "0011111101001100000100",
			668 => "0000000000101100000001",
			669 => "0000000000101100000001",
			670 => "0011001110011000000100",
			671 => "0000000000101100000001",
			672 => "0000000000101100000001",
			673 => "0011011100101000010000",
			674 => "0000000000000000001100",
			675 => "0000111001010100000100",
			676 => "0000000000101100000001",
			677 => "0000001010000000000100",
			678 => "0000000000101100000001",
			679 => "0000000000101100000001",
			680 => "0000000000101100000001",
			681 => "0000100100010100010100",
			682 => "0000101100010100001000",
			683 => "0000000111011000000100",
			684 => "0000000000101100000001",
			685 => "0000000000101100000001",
			686 => "0000110011000100000100",
			687 => "0000000000101100000001",
			688 => "0000110000111100000100",
			689 => "0000000000101100000001",
			690 => "0000000000101100000001",
			691 => "0011011101101000001100",
			692 => "0001001000000000001000",
			693 => "0001011011111000000100",
			694 => "0000000000101100000001",
			695 => "0000000000101100000001",
			696 => "0000000000101100000001",
			697 => "0001000110101100000100",
			698 => "0000000000101100000001",
			699 => "0010001100110000000100",
			700 => "0000000000101100000001",
			701 => "0001111110001100000100",
			702 => "0000000000101100000001",
			703 => "0000000000101100000001",
			704 => "0011010011000000110100",
			705 => "0011100101001100101100",
			706 => "0000100101010000100100",
			707 => "0000011100101000100000",
			708 => "0001101100111000010000",
			709 => "0000010110001100001000",
			710 => "0001111011111000000100",
			711 => "0000000000101101101101",
			712 => "1111111000101101101101",
			713 => "0000010111011100000100",
			714 => "0000000000101101101101",
			715 => "0000000000101101101101",
			716 => "0011100100101000001000",
			717 => "0011101110100100000100",
			718 => "0000000000101101101101",
			719 => "1111111000101101101101",
			720 => "0001111100011100000100",
			721 => "0000000000101101101101",
			722 => "1111111000101101101101",
			723 => "0000000000101101101101",
			724 => "0001001001000100000100",
			725 => "0000000000101101101101",
			726 => "0000001000101101101101",
			727 => "0000111001010000000100",
			728 => "0000000000101101101101",
			729 => "1111111000101101101101",
			730 => "1111111000101101101101",
			731 => "0010101100001101010000",
			732 => "0001011000100000110100",
			733 => "0010111101101000101000",
			734 => "0010001010000100010000",
			735 => "0011000101011100001100",
			736 => "0010011101101000001000",
			737 => "0010111011101100000100",
			738 => "0000000000110000011001",
			739 => "0000000000110000011001",
			740 => "0000000000110000011001",
			741 => "0000000000110000011001",
			742 => "0000001010111000010000",
			743 => "0011111000001000001000",
			744 => "0001101010111100000100",
			745 => "0000000000110000011001",
			746 => "0000000000110000011001",
			747 => "0000111001010100000100",
			748 => "0000000000110000011001",
			749 => "0000000000110000011001",
			750 => "0011010101101100000100",
			751 => "0000001000110000011001",
			752 => "0000000000110000011001",
			753 => "0000010111011100001000",
			754 => "0010011100110000000100",
			755 => "0000000000110000011001",
			756 => "0000000000110000011001",
			757 => "0000000000110000011001",
			758 => "0010000011001000010100",
			759 => "0011001001001000001100",
			760 => "0011110010111100001000",
			761 => "0000001011001000000100",
			762 => "0000000000110000011001",
			763 => "0000000000110000011001",
			764 => "0000000000110000011001",
			765 => "0010101001000000000100",
			766 => "0000000000110000011001",
			767 => "0000000000110000011001",
			768 => "0000100101101000000100",
			769 => "1111111000110000011001",
			770 => "0000000000110000011001",
			771 => "0000001100100100000100",
			772 => "0000000000110000011001",
			773 => "0000000000110000011001",
			774 => "0001110011110101001100",
			775 => "0011111010101100011000",
			776 => "0000011000011000001100",
			777 => "0010111010100100001000",
			778 => "0000110011001000000100",
			779 => "0000000000110010110101",
			780 => "0000000000110010110101",
			781 => "0000000000110010110101",
			782 => "0000110011000000001000",
			783 => "0000111001000100000100",
			784 => "0000000000110010110101",
			785 => "0000000000110010110101",
			786 => "0000000000110010110101",
			787 => "0011110101100100100000",
			788 => "0000001110110000010100",
			789 => "0000001111001100010000",
			790 => "0011000101101100001000",
			791 => "0000011001100000000100",
			792 => "0000000000110010110101",
			793 => "0000000000110010110101",
			794 => "0011100110111000000100",
			795 => "0000000000110010110101",
			796 => "0000000000110010110101",
			797 => "0000000000110010110101",
			798 => "0000011101000000001000",
			799 => "0011101111010100000100",
			800 => "0000000000110010110101",
			801 => "0000000000110010110101",
			802 => "0000000000110010110101",
			803 => "0000001000110000010000",
			804 => "0001011011111000001100",
			805 => "0000001010111000000100",
			806 => "0000000000110010110101",
			807 => "0001101110000100000100",
			808 => "0000000000110010110101",
			809 => "0000000000110010110101",
			810 => "0000000000110010110101",
			811 => "0000000000110010110101",
			812 => "0000000000110010110101",
			813 => "0001110011110101011000",
			814 => "0000000110101000101000",
			815 => "0011111110101100011100",
			816 => "0011110000001100011000",
			817 => "0001100011011000001100",
			818 => "0011110010110000000100",
			819 => "0000000000110110000001",
			820 => "0011011010100100000100",
			821 => "0000000000110110000001",
			822 => "0000000000110110000001",
			823 => "0000110011001000001000",
			824 => "0010011100101000000100",
			825 => "0000000000110110000001",
			826 => "0000000000110110000001",
			827 => "0000000000110110000001",
			828 => "0000000000110110000001",
			829 => "0001001100101000001000",
			830 => "0001110100101100000100",
			831 => "0000000000110110000001",
			832 => "0000000000110110000001",
			833 => "1111111000110110000001",
			834 => "0011011001000100100000",
			835 => "0001111001011000010100",
			836 => "0000010110001100010000",
			837 => "0001101010101100001000",
			838 => "0000000101010000000100",
			839 => "1111111000110110000001",
			840 => "0000000000110110000001",
			841 => "0011110101100100000100",
			842 => "0000000000110110000001",
			843 => "0000000000110110000001",
			844 => "0000000000110110000001",
			845 => "0001101110000100001000",
			846 => "0000010011010000000100",
			847 => "0000000000110110000001",
			848 => "1111111000110110000001",
			849 => "0000000000110110000001",
			850 => "0000111011111000001000",
			851 => "0010011000111000000100",
			852 => "0000001000110110000001",
			853 => "0000000000110110000001",
			854 => "0001001111101000000100",
			855 => "0000000000110110000001",
			856 => "0000000000110110000001",
			857 => "0011000011000000000100",
			858 => "0000000000110110000001",
			859 => "0000001010010000000100",
			860 => "0000000000110110000001",
			861 => "0000101001101000000100",
			862 => "0000000000110110000001",
			863 => "0000000000110110000001",
			864 => "0011110010110000000100",
			865 => "1111111000110111111101",
			866 => "0011100101001100110100",
			867 => "0000100101010000101000",
			868 => "0000011100101000100000",
			869 => "0011110101100100010000",
			870 => "0011000101101100001000",
			871 => "0010001111001000000100",
			872 => "0000000000110111111101",
			873 => "0000000000110111111101",
			874 => "0011011010000100000100",
			875 => "0000000000110111111101",
			876 => "0000001000110111111101",
			877 => "0001100000000100001000",
			878 => "0000101111001100000100",
			879 => "1111111000110111111101",
			880 => "0000000000110111111101",
			881 => "0001111100011100000100",
			882 => "0000001000110111111101",
			883 => "1111111000110111111101",
			884 => "0010001100110000000100",
			885 => "0000001000110111111101",
			886 => "1111111000110111111101",
			887 => "0001000101111000001000",
			888 => "0000101000001100000100",
			889 => "0000000000110111111101",
			890 => "0000000000110111111101",
			891 => "0000001000110111111101",
			892 => "0000111001010000000100",
			893 => "0000000000110111111101",
			894 => "1111111000110111111101",
			895 => "0001101111110000000100",
			896 => "1111111000111001100001",
			897 => "0010010110101100101100",
			898 => "0000011100101000100100",
			899 => "0010111010000100100000",
			900 => "0010110101011100010000",
			901 => "0000010011110000001000",
			902 => "0010111010100100000100",
			903 => "0000000000111001100001",
			904 => "1111111000111001100001",
			905 => "0011110101100100000100",
			906 => "0000001000111001100001",
			907 => "0000000000111001100001",
			908 => "0000101100001000001000",
			909 => "0010101011000000000100",
			910 => "1111111000111001100001",
			911 => "0000000000111001100001",
			912 => "0001011011111000000100",
			913 => "0000000000111001100001",
			914 => "0000000000111001100001",
			915 => "0000001000111001100001",
			916 => "0000111011111000000100",
			917 => "0000001000111001100001",
			918 => "0000000000111001100001",
			919 => "1111111000111001100001",
			920 => "0010001000000001100100",
			921 => "0001110110011101001000",
			922 => "0011000101010100101000",
			923 => "0001010011001000001100",
			924 => "0000110011000000001000",
			925 => "0000111101101000000100",
			926 => "0000000000111101000101",
			927 => "0000000000111101000101",
			928 => "0000000000111101000101",
			929 => "0001011001010000010000",
			930 => "0011110100010000001000",
			931 => "0000110011000000000100",
			932 => "0000000000111101000101",
			933 => "0000000000111101000101",
			934 => "0010001111111100000100",
			935 => "0000000000111101000101",
			936 => "0000000000111101000101",
			937 => "0001001010000100000100",
			938 => "0000000000111101000101",
			939 => "0011101111010100000100",
			940 => "0000000000111101000101",
			941 => "0000000000111101000101",
			942 => "0010001111011000010000",
			943 => "0001010011000100001000",
			944 => "0001001100000000000100",
			945 => "0000000000111101000101",
			946 => "0000000000111101000101",
			947 => "0001001100110000000100",
			948 => "0000000000111101000101",
			949 => "0000000000111101000101",
			950 => "0011000101101100001000",
			951 => "0000000110101000000100",
			952 => "0000000000111101000101",
			953 => "0000000000111101000101",
			954 => "0001011110111000000100",
			955 => "0000000000111101000101",
			956 => "0000000000111101000101",
			957 => "0010101011000000001100",
			958 => "0011100100111000000100",
			959 => "0000000000111101000101",
			960 => "0010001010000100000100",
			961 => "0000000000111101000101",
			962 => "0000000000111101000101",
			963 => "0000111011000000001000",
			964 => "0010000011001000000100",
			965 => "0000000000111101000101",
			966 => "0000000000111101000101",
			967 => "0011001101101000000100",
			968 => "0000000000111101000101",
			969 => "0000000000111101000101",
			970 => "0000101111001100001000",
			971 => "0010111001000100000100",
			972 => "0000000000111101000101",
			973 => "0000000000111101000101",
			974 => "0000111001010000000100",
			975 => "0000000000111101000101",
			976 => "0000000000111101000101",
			977 => "0010001010000100110000",
			978 => "0000100101010000101100",
			979 => "0001101100000100100000",
			980 => "0011101001011100001100",
			981 => "0010111011101100001000",
			982 => "0010110110001100000100",
			983 => "0000000001000000111001",
			984 => "0000000001000000111001",
			985 => "0000000001000000111001",
			986 => "0001101110010000001100",
			987 => "0010101100010000000100",
			988 => "0000000001000000111001",
			989 => "0010110111011100000100",
			990 => "0000000001000000111001",
			991 => "0000000001000000111001",
			992 => "0011111110000100000100",
			993 => "0000000001000000111001",
			994 => "0000000001000000111001",
			995 => "0001001100000000001000",
			996 => "0001111100110000000100",
			997 => "0000000001000000111001",
			998 => "0000000001000000111001",
			999 => "0000000001000000111001",
			1000 => "0000000001000000111001",
			1001 => "0010111001001000011100",
			1002 => "0000100110010100010000",
			1003 => "0001100100000100001100",
			1004 => "0001001000000100001000",
			1005 => "0001011000000000000100",
			1006 => "0000000001000000111001",
			1007 => "0000000001000000111001",
			1008 => "0000000001000000111001",
			1009 => "0000000001000000111001",
			1010 => "0001011000100000001000",
			1011 => "0011010101011100000100",
			1012 => "0000000001000000111001",
			1013 => "0000000001000000111001",
			1014 => "0000000001000000111001",
			1015 => "0011100110111000010000",
			1016 => "0000111100110000001000",
			1017 => "0010001000000000000100",
			1018 => "0000000001000000111001",
			1019 => "0000000001000000111001",
			1020 => "0010101111100100000100",
			1021 => "0000000001000000111001",
			1022 => "0000000001000000111001",
			1023 => "0011101010001000001000",
			1024 => "0010100011000100000100",
			1025 => "0000000001000000111001",
			1026 => "0000000001000000111001",
			1027 => "0000010111011100001100",
			1028 => "0011000110000000000100",
			1029 => "0000000001000000111001",
			1030 => "0000010011010000000100",
			1031 => "0000000001000000111001",
			1032 => "0000000001000000111001",
			1033 => "0000011100101000000100",
			1034 => "0000000001000000111001",
			1035 => "0010010110101100000100",
			1036 => "0000000001000000111001",
			1037 => "0000000001000000111001",
			1038 => "0000101110000100000100",
			1039 => "1111111001000011010101",
			1040 => "0001011000100000101100",
			1041 => "0001001000111000100100",
			1042 => "0011011101101000011100",
			1043 => "0011011100101000010000",
			1044 => "0011000101010100001000",
			1045 => "0011010110001100000100",
			1046 => "0000000001000011010101",
			1047 => "0000000001000011010101",
			1048 => "0001100100110000000100",
			1049 => "0000000001000011010101",
			1050 => "1111111001000011010101",
			1051 => "0000111000101000001000",
			1052 => "0000111001010100000100",
			1053 => "0000000001000011010101",
			1054 => "0000000001000011010101",
			1055 => "0000001001000011010101",
			1056 => "0010001001010100000100",
			1057 => "1111111001000011010101",
			1058 => "0000000001000011010101",
			1059 => "0001101101010000000100",
			1060 => "0000000001000011010101",
			1061 => "0000001001000011010101",
			1062 => "0010101100001100011000",
			1063 => "0011000101011100001000",
			1064 => "0000001000010000000100",
			1065 => "0000000001000011010101",
			1066 => "0000000001000011010101",
			1067 => "0010101011111000000100",
			1068 => "0000000001000011010101",
			1069 => "0010001111011000001000",
			1070 => "0001001011111000000100",
			1071 => "0000000001000011010101",
			1072 => "0000000001000011010101",
			1073 => "1111111001000011010101",
			1074 => "0000000000101000000100",
			1075 => "0000000001000011010101",
			1076 => "0000001001000011010101",
			1077 => "0000100100010101000000",
			1078 => "0000110100101100110100",
			1079 => "0010101001010100011100",
			1080 => "0010000011100100010100",
			1081 => "0010010101101100010000",
			1082 => "0010111010100100001000",
			1083 => "0011110000001100000100",
			1084 => "0000000001000111000001",
			1085 => "0000000001000111000001",
			1086 => "0001000101010100000100",
			1087 => "0000000001000111000001",
			1088 => "0000000001000111000001",
			1089 => "0000000001000111000001",
			1090 => "0010001000000000000100",
			1091 => "0000000001000111000001",
			1092 => "0000000001000111000001",
			1093 => "0010000011100100010000",
			1094 => "0011100011101000001100",
			1095 => "0000000110111100001000",
			1096 => "0001101111110000000100",
			1097 => "0000000001000111000001",
			1098 => "0000000001000111000001",
			1099 => "0000000001000111000001",
			1100 => "0000000001000111000001",
			1101 => "0010101001011000000100",
			1102 => "0000000001000111000001",
			1103 => "0000000001000111000001",
			1104 => "0000111110001100000100",
			1105 => "0000000001000111000001",
			1106 => "0001011111100000000100",
			1107 => "0000000001000111000001",
			1108 => "0000000001000111000001",
			1109 => "0001101000010100010100",
			1110 => "0001110100101100010000",
			1111 => "0011001010100100000100",
			1112 => "0000000001000111000001",
			1113 => "0001100101100000000100",
			1114 => "0000000001000111000001",
			1115 => "0001011001010100000100",
			1116 => "0000000001000111000001",
			1117 => "0000000001000111000001",
			1118 => "0000000001000111000001",
			1119 => "0000100111111000001000",
			1120 => "0011000101010100000100",
			1121 => "0000000001000111000001",
			1122 => "0000000001000111000001",
			1123 => "0010101101001000000100",
			1124 => "0000000001000111000001",
			1125 => "0000111001010000001000",
			1126 => "0011110100110100000100",
			1127 => "0000000001000111000001",
			1128 => "0000000001000111000001",
			1129 => "0010101001011000001000",
			1130 => "0011001001001000000100",
			1131 => "0000000001000111000001",
			1132 => "0000000001000111000001",
			1133 => "0001100010111100000100",
			1134 => "0000000001000111000001",
			1135 => "0000000001000111000001",
			1136 => "0000010011110000110100",
			1137 => "0010111010100100110000",
			1138 => "0001011000000000010000",
			1139 => "0000110011000000001000",
			1140 => "0011101111110100000100",
			1141 => "0000000001001011000101",
			1142 => "0000000001001011000101",
			1143 => "0011101100000100000100",
			1144 => "0000000001001011000101",
			1145 => "0000000001001011000101",
			1146 => "0010101000101000010000",
			1147 => "0010101101001000001000",
			1148 => "0011101001011100000100",
			1149 => "0000000001001011000101",
			1150 => "0000000001001011000101",
			1151 => "0010001111111100000100",
			1152 => "0000000001001011000101",
			1153 => "0000000001001011000101",
			1154 => "0000111001010100001000",
			1155 => "0001011001010000000100",
			1156 => "0000000001001011000101",
			1157 => "0000000001001011000101",
			1158 => "0000100110111100000100",
			1159 => "0000000001001011000101",
			1160 => "0000000001001011000101",
			1161 => "0000000001001011000101",
			1162 => "0010111001001000101000",
			1163 => "0011011100101000100000",
			1164 => "0010110101010100010100",
			1165 => "0001010011001000000100",
			1166 => "0000000001001011000101",
			1167 => "0000111000000000001000",
			1168 => "0001100101001000000100",
			1169 => "0000000001001011000101",
			1170 => "0000000001001011000101",
			1171 => "0000111001010100000100",
			1172 => "0000000001001011000101",
			1173 => "0000000001001011000101",
			1174 => "0011101100011000001000",
			1175 => "0010010101111000000100",
			1176 => "0000000001001011000101",
			1177 => "0000000001001011000101",
			1178 => "0000000001001011000101",
			1179 => "0000001101111000000100",
			1180 => "0000000001001011000101",
			1181 => "0000000001001011000101",
			1182 => "0011011001000100010000",
			1183 => "0000001010111000001100",
			1184 => "0010001111011000001000",
			1185 => "0010000000110000000100",
			1186 => "0000000001001011000101",
			1187 => "0000000001001011000101",
			1188 => "0000000001001011000101",
			1189 => "0000000001001011000101",
			1190 => "0001101010110000010000",
			1191 => "0011111001111000001000",
			1192 => "0001011111111000000100",
			1193 => "0000000001001011000101",
			1194 => "0000000001001011000101",
			1195 => "0011100100011100000100",
			1196 => "0000000001001011000101",
			1197 => "0000000001001011000101",
			1198 => "0010011100010000000100",
			1199 => "0000000001001011000101",
			1200 => "0000000001001011000101",
			1201 => "0010000101101100000100",
			1202 => "1111111001001101001001",
			1203 => "0011110010110000000100",
			1204 => "1111111001001101001001",
			1205 => "0010110111011100011000",
			1206 => "0001000101010100001000",
			1207 => "0011011110011000000100",
			1208 => "0000000001001101001001",
			1209 => "1111111001001101001001",
			1210 => "0001011001010000001000",
			1211 => "0001111111101000000100",
			1212 => "0000001001001101001001",
			1213 => "0000000001001101001001",
			1214 => "0010101011111000000100",
			1215 => "0000000001001101001001",
			1216 => "0000001001001101001001",
			1217 => "0010000000110000010000",
			1218 => "0010100001011100001100",
			1219 => "0001101110010000001000",
			1220 => "0011100011010100000100",
			1221 => "1111111001001101001001",
			1222 => "0000000001001101001001",
			1223 => "1111111001001101001001",
			1224 => "0000001001001101001001",
			1225 => "0011010101111000010000",
			1226 => "0000001011001100001000",
			1227 => "0000000110100100000100",
			1228 => "0000000001001101001001",
			1229 => "1111111001001101001001",
			1230 => "0000010101011100000100",
			1231 => "0000001001001101001001",
			1232 => "1111111001001101001001",
			1233 => "1111111001001101001001",
			1234 => "0000010011110000110100",
			1235 => "0010111010100100110000",
			1236 => "0001011000000000010000",
			1237 => "0000110011000000001000",
			1238 => "0011101111110100000100",
			1239 => "0000000001010001011101",
			1240 => "0000000001010001011101",
			1241 => "0011101100000100000100",
			1242 => "0000000001010001011101",
			1243 => "0000000001010001011101",
			1244 => "0010101000101000010000",
			1245 => "0010101101001000001000",
			1246 => "0011101001011100000100",
			1247 => "0000000001010001011101",
			1248 => "0000000001010001011101",
			1249 => "0010001111111100000100",
			1250 => "0000000001010001011101",
			1251 => "0000000001010001011101",
			1252 => "0000111001010100001000",
			1253 => "0001011001010000000100",
			1254 => "0000000001010001011101",
			1255 => "0000000001010001011101",
			1256 => "0000100110111100000100",
			1257 => "0000000001010001011101",
			1258 => "0000000001010001011101",
			1259 => "0000000001010001011101",
			1260 => "0010111001001000101000",
			1261 => "0001001000000100011100",
			1262 => "0001000110000000010000",
			1263 => "0011000111011100001000",
			1264 => "0001010011001000000100",
			1265 => "0000000001010001011101",
			1266 => "0000000001010001011101",
			1267 => "0001000111011100000100",
			1268 => "0000000001010001011101",
			1269 => "0000000001010001011101",
			1270 => "0011110000010000000100",
			1271 => "0000000001010001011101",
			1272 => "0011010101010100000100",
			1273 => "0000000001010001011101",
			1274 => "0000000001010001011101",
			1275 => "0000110011000100001000",
			1276 => "0011101100011000000100",
			1277 => "0000000001010001011101",
			1278 => "0000000001010001011101",
			1279 => "0000000001010001011101",
			1280 => "0000111100110000010000",
			1281 => "0011011101101000001100",
			1282 => "0011010101101100001000",
			1283 => "0011011001001000000100",
			1284 => "0000000001010001011101",
			1285 => "0000000001010001011101",
			1286 => "0000000001010001011101",
			1287 => "0000000001010001011101",
			1288 => "0011011010000100010000",
			1289 => "0000001101011000001100",
			1290 => "0010001111011000001000",
			1291 => "0010000000110000000100",
			1292 => "0000000001010001011101",
			1293 => "0000000001010001011101",
			1294 => "0000000001010001011101",
			1295 => "0000000001010001011101",
			1296 => "0000010101011100001100",
			1297 => "0011100100011100001000",
			1298 => "0000101100001000000100",
			1299 => "0000000001010001011101",
			1300 => "0000000001010001011101",
			1301 => "0000000001010001011101",
			1302 => "0000000001010001011101",
			1303 => "0010000101101100001000",
			1304 => "0000010011110000000100",
			1305 => "1111111001010100101001",
			1306 => "0000000001010100101001",
			1307 => "0011000101010100100000",
			1308 => "0001001010000100010100",
			1309 => "0000011101000000010000",
			1310 => "0010111010100100001100",
			1311 => "0000000100010100001000",
			1312 => "0001001001001000000100",
			1313 => "1111111001010100101001",
			1314 => "0000000001010100101001",
			1315 => "0000001001010100101001",
			1316 => "1111111001010100101001",
			1317 => "0000001001010100101001",
			1318 => "0011011110011000000100",
			1319 => "0000000001010100101001",
			1320 => "0001101111110000000100",
			1321 => "0000000001010100101001",
			1322 => "0000001001010100101001",
			1323 => "0000010110001100100100",
			1324 => "0001011100101100010100",
			1325 => "0011011100101000001100",
			1326 => "0010110101010100001000",
			1327 => "0010011101101000000100",
			1328 => "0000000001010100101001",
			1329 => "0000000001010100101001",
			1330 => "1111111001010100101001",
			1331 => "0000111100010000000100",
			1332 => "0000000001010100101001",
			1333 => "0000001001010100101001",
			1334 => "0010011101101000000100",
			1335 => "0000000001010100101001",
			1336 => "0011011001001000000100",
			1337 => "1111111001010100101001",
			1338 => "0011010101101100000100",
			1339 => "0000000001010100101001",
			1340 => "1111111001010100101001",
			1341 => "0001001001000100001100",
			1342 => "0001000011010000001000",
			1343 => "0001001010100100000100",
			1344 => "0000000001010100101001",
			1345 => "0000000001010100101001",
			1346 => "1111111001010100101001",
			1347 => "0011110100001000000100",
			1348 => "1111111001010100101001",
			1349 => "0000111100010000000100",
			1350 => "0000001001010100101001",
			1351 => "0001011011111000000100",
			1352 => "1111111001010100101001",
			1353 => "0000000001010100101001",
			1354 => "0000100101010001100100",
			1355 => "0011110101100101001100",
			1356 => "0011100100101000110000",
			1357 => "0011000101101100011100",
			1358 => "0000011101000000010000",
			1359 => "0010111011101100001000",
			1360 => "0011011011101100000100",
			1361 => "0000000001011000000101",
			1362 => "0000001001011000000101",
			1363 => "0001011100101100000100",
			1364 => "0000000001011000000101",
			1365 => "1111111001011000000101",
			1366 => "0011110101111100001000",
			1367 => "0011111100111000000100",
			1368 => "0000000001011000000101",
			1369 => "0000001001011000000101",
			1370 => "0000000001011000000101",
			1371 => "0000110000111000001100",
			1372 => "0010001111011000001000",
			1373 => "0001111011111000000100",
			1374 => "0000000001011000000101",
			1375 => "0000000001011000000101",
			1376 => "1111111001011000000101",
			1377 => "0001001100110100000100",
			1378 => "0000001001011000000101",
			1379 => "0000000001011000000101",
			1380 => "0001011001010000001000",
			1381 => "0000101011100000000100",
			1382 => "0000000001011000000101",
			1383 => "0000001001011000000101",
			1384 => "0000111000101000000100",
			1385 => "0000000001011000000101",
			1386 => "0000111011111000001000",
			1387 => "0000010111011100000100",
			1388 => "0000001001011000000101",
			1389 => "0000000001011000000101",
			1390 => "0001101000010100000100",
			1391 => "0000000001011000000101",
			1392 => "0000000001011000000101",
			1393 => "0010000000110000001100",
			1394 => "0001111001010000000100",
			1395 => "0000000001011000000101",
			1396 => "0000111001010100000100",
			1397 => "1111111001011000000101",
			1398 => "0000000001011000000101",
			1399 => "0011011101101000001000",
			1400 => "0001011100101100000100",
			1401 => "0000000001011000000101",
			1402 => "0000000001011000000101",
			1403 => "1111111001011000000101",
			1404 => "0001100000100100001000",
			1405 => "0011100101100000000100",
			1406 => "0000001001011000000101",
			1407 => "0000000001011000000101",
			1408 => "0000000001011000000101",
			1409 => "0011110010110000000100",
			1410 => "1111111001011010100001",
			1411 => "0011100101001101000100",
			1412 => "0000001101011000110000",
			1413 => "0011110101100100011100",
			1414 => "0001011100101100001100",
			1415 => "0010001111111100000100",
			1416 => "1111111001011010100001",
			1417 => "0001010011001000000100",
			1418 => "1111111001011010100001",
			1419 => "0000000001011010100001",
			1420 => "0000010110001100001000",
			1421 => "0011000101010100000100",
			1422 => "0000000001011010100001",
			1423 => "1111111001011010100001",
			1424 => "0011000101101100000100",
			1425 => "0000001001011010100001",
			1426 => "0000000001011010100001",
			1427 => "0001101110000100001000",
			1428 => "0011110000101100000100",
			1429 => "1111111001011010100001",
			1430 => "1111111001011010100001",
			1431 => "0001111100011100001000",
			1432 => "0010011001001000000100",
			1433 => "1111111001011010100001",
			1434 => "0000001001011010100001",
			1435 => "1111111001011010100001",
			1436 => "0001111011111000001000",
			1437 => "0000100101010000000100",
			1438 => "1111111001011010100001",
			1439 => "0000001001011010100001",
			1440 => "0011000101111000001000",
			1441 => "0001010110011100000100",
			1442 => "0000001001011010100001",
			1443 => "0000001001011010100001",
			1444 => "1111111001011010100001",
			1445 => "0000101101011000000100",
			1446 => "1111111001011010100001",
			1447 => "0000000001011010100001",
			1448 => "0000010111100100000100",
			1449 => "1111111001011101001101",
			1450 => "0001011001010000100100",
			1451 => "0010001000000000100000",
			1452 => "0000001101001100000100",
			1453 => "0000000001011101001101",
			1454 => "0010001001000100001100",
			1455 => "0000001001101000001000",
			1456 => "0001011000000100000100",
			1457 => "0000000001011101001101",
			1458 => "0000000001011101001101",
			1459 => "0000000001011101001101",
			1460 => "0011111100111100001000",
			1461 => "0011100001000100000100",
			1462 => "0000000001011101001101",
			1463 => "0000000001011101001101",
			1464 => "0000111100010000000100",
			1465 => "0000001001011101001101",
			1466 => "0000000001011101001101",
			1467 => "0000000001011101001101",
			1468 => "0000100110010100010100",
			1469 => "0000101100010100001000",
			1470 => "0000100011011100000100",
			1471 => "0000000001011101001101",
			1472 => "0000000001011101001101",
			1473 => "0010101011000000000100",
			1474 => "1111111001011101001101",
			1475 => "0001001100010000000100",
			1476 => "0000000001011101001101",
			1477 => "0000000001011101001101",
			1478 => "0001000011000000001000",
			1479 => "0001010100101100000100",
			1480 => "0000000001011101001101",
			1481 => "0000001001011101001101",
			1482 => "0000000110100100000100",
			1483 => "0000000001011101001101",
			1484 => "0010001100110000001000",
			1485 => "0011000101011100000100",
			1486 => "0000000001011101001101",
			1487 => "0000000001011101001101",
			1488 => "0000111001010100000100",
			1489 => "0000000001011101001101",
			1490 => "0000000001011101001101",
			1491 => "0011010101111001100100",
			1492 => "0000010110001100111000",
			1493 => "0010111011101100001100",
			1494 => "0001010011001000000100",
			1495 => "0000000001100000011001",
			1496 => "0010001111111100000100",
			1497 => "0000000001100000011001",
			1498 => "0000001001100000011001",
			1499 => "0010001111001000010100",
			1500 => "0000110011001000001100",
			1501 => "0011100101110100000100",
			1502 => "0000000001100000011001",
			1503 => "0001111000101000000100",
			1504 => "0000000001100000011001",
			1505 => "0000000001100000011001",
			1506 => "0001001010100100000100",
			1507 => "0000000001100000011001",
			1508 => "1111111001100000011001",
			1509 => "0011100100101000010000",
			1510 => "0001011001010000001000",
			1511 => "0001011000000000000100",
			1512 => "0000000001100000011001",
			1513 => "0000000001100000011001",
			1514 => "0011011100101000000100",
			1515 => "1111111001100000011001",
			1516 => "0000000001100000011001",
			1517 => "0011000101010100000100",
			1518 => "0000001001100000011001",
			1519 => "0000000001100000011001",
			1520 => "0001111001011000010000",
			1521 => "0010010011000000001000",
			1522 => "0001011001010100000100",
			1523 => "0000000001100000011001",
			1524 => "0000000001100000011001",
			1525 => "0011110100001000000100",
			1526 => "0000000001100000011001",
			1527 => "0000001001100000011001",
			1528 => "0001111000100000000100",
			1529 => "0000000001100000011001",
			1530 => "0001010011000100001100",
			1531 => "0001011011111000000100",
			1532 => "0000000001100000011001",
			1533 => "0000010111011100000100",
			1534 => "0000001001100000011001",
			1535 => "0000000001100000011001",
			1536 => "0000110000111100001000",
			1537 => "0000010101010100000100",
			1538 => "1111111001100000011001",
			1539 => "0000000001100000011001",
			1540 => "0000000001100000011001",
			1541 => "1111111001100000011001",
			1542 => "0000101010010001011100",
			1543 => "0001100111010001001100",
			1544 => "0011000101010100011100",
			1545 => "0010001001000100010000",
			1546 => "0010111011101100001000",
			1547 => "0010011100101000000100",
			1548 => "0000000001100011010101",
			1549 => "0000000001100011010101",
			1550 => "0001111011111000000100",
			1551 => "0000000001100011010101",
			1552 => "0000000001100011010101",
			1553 => "0000001101001100000100",
			1554 => "0000000001100011010101",
			1555 => "0011111011010100000100",
			1556 => "0000000001100011010101",
			1557 => "0000000001100011010101",
			1558 => "0010100000111100100000",
			1559 => "0001111000100000010000",
			1560 => "0000000110111100001000",
			1561 => "0000001111101100000100",
			1562 => "0000000001100011010101",
			1563 => "0000000001100011010101",
			1564 => "0010000011001000000100",
			1565 => "0000000001100011010101",
			1566 => "0000000001100011010101",
			1567 => "0010001000000000001000",
			1568 => "0011100110111000000100",
			1569 => "0000000001100011010101",
			1570 => "0000000001100011010101",
			1571 => "0010001001010100000100",
			1572 => "0000000001100011010101",
			1573 => "0000000001100011010101",
			1574 => "0000000101101000001100",
			1575 => "0011110111010000001000",
			1576 => "0000100010100100000100",
			1577 => "0000000001100011010101",
			1578 => "0000000001100011010101",
			1579 => "0000000001100011010101",
			1580 => "0000000001100011010101",
			1581 => "0011110100110100000100",
			1582 => "0000000001100011010101",
			1583 => "0000011100101000000100",
			1584 => "0000000001100011010101",
			1585 => "0000011111001000000100",
			1586 => "0000000001100011010101",
			1587 => "0000000001100011010101",
			1588 => "0000000001100011010101",
			1589 => "0001011000000000010100",
			1590 => "0001111100010000001000",
			1591 => "0001111000111000000100",
			1592 => "0000000001100111101001",
			1593 => "0000000001100111101001",
			1594 => "0001000110000000001000",
			1595 => "0011101000110100000100",
			1596 => "0000000001100111101001",
			1597 => "0000000001100111101001",
			1598 => "0000000001100111101001",
			1599 => "0011000101010100100100",
			1600 => "0000101100001000011000",
			1601 => "0001111000101000010100",
			1602 => "0010001111001000010000",
			1603 => "0000001100111100001000",
			1604 => "0000101110010000000100",
			1605 => "0000000001100111101001",
			1606 => "0000000001100111101001",
			1607 => "0011100001101100000100",
			1608 => "0000000001100111101001",
			1609 => "0000000001100111101001",
			1610 => "0000000001100111101001",
			1611 => "0000000001100111101001",
			1612 => "0010000101101100000100",
			1613 => "0000000001100111101001",
			1614 => "0001101010101100000100",
			1615 => "0000000001100111101001",
			1616 => "0000000001100111101001",
			1617 => "0011011100101000100000",
			1618 => "0010110011010000001000",
			1619 => "0000110100101100000100",
			1620 => "0000000001100111101001",
			1621 => "0000000001100111101001",
			1622 => "0010101001011000001000",
			1623 => "0010010110000000000100",
			1624 => "0000000001100111101001",
			1625 => "0000000001100111101001",
			1626 => "0010110101010100001000",
			1627 => "0010011101101000000100",
			1628 => "0000000001100111101001",
			1629 => "0000000001100111101001",
			1630 => "0010100001011100000100",
			1631 => "0000000001100111101001",
			1632 => "0000000001100111101001",
			1633 => "0000101111001100100000",
			1634 => "0011111011110100010000",
			1635 => "0011111100111100001000",
			1636 => "0000101100010100000100",
			1637 => "0000000001100111101001",
			1638 => "0000000001100111101001",
			1639 => "0001111110111000000100",
			1640 => "0000000001100111101001",
			1641 => "0000000001100111101001",
			1642 => "0000111111101000001000",
			1643 => "0001100101111100000100",
			1644 => "0000000001100111101001",
			1645 => "0000000001100111101001",
			1646 => "0000001110110000000100",
			1647 => "0000000001100111101001",
			1648 => "0000000001100111101001",
			1649 => "0000010101011100001000",
			1650 => "0001110011110100000100",
			1651 => "0000000001100111101001",
			1652 => "0000000001100111101001",
			1653 => "0011110011100000001000",
			1654 => "0011110011111100000100",
			1655 => "0000000001100111101001",
			1656 => "0000000001100111101001",
			1657 => "0000000001100111101001",
			1658 => "0000010111100100000100",
			1659 => "1111111001101010111111",
			1660 => "0001011001010000100100",
			1661 => "0010001000000000100000",
			1662 => "0000001101001100000100",
			1663 => "0000000001101010111111",
			1664 => "0010001001000100001100",
			1665 => "0001111101001000000100",
			1666 => "0000000001101010111111",
			1667 => "0010101000101000000100",
			1668 => "0000000001101010111111",
			1669 => "0000000001101010111111",
			1670 => "0011111100111100001000",
			1671 => "0011100001000100000100",
			1672 => "0000000001101010111111",
			1673 => "0000000001101010111111",
			1674 => "0000111100010000000100",
			1675 => "0000001001101010111111",
			1676 => "0000000001101010111111",
			1677 => "0000000001101010111111",
			1678 => "0010001010000100010000",
			1679 => "0011000011010000000100",
			1680 => "0000000001101010111111",
			1681 => "0001010011000100000100",
			1682 => "1111111001101010111111",
			1683 => "0001011100110100000100",
			1684 => "0000000001101010111111",
			1685 => "0000000001101010111111",
			1686 => "0000100000101000011100",
			1687 => "0011000101101100001100",
			1688 => "0010001111011000000100",
			1689 => "0000000001101010111111",
			1690 => "0010011111011000000100",
			1691 => "0000000001101010111111",
			1692 => "0000000001101010111111",
			1693 => "0001001010011100001000",
			1694 => "0001111001011000000100",
			1695 => "0000000001101010111111",
			1696 => "1111111001101010111111",
			1697 => "0001000111010100000100",
			1698 => "0000000001101010111111",
			1699 => "0000000001101010111111",
			1700 => "0001110001011000001000",
			1701 => "0010101011000000000100",
			1702 => "0000001001101010111111",
			1703 => "0000000001101010111111",
			1704 => "0001010011000100001000",
			1705 => "0000010101011100000100",
			1706 => "0000000001101010111111",
			1707 => "0000000001101010111111",
			1708 => "0000000010100000000100",
			1709 => "1111111001101010111111",
			1710 => "0000000001101010111111",
			1711 => "0001101010001000010000",
			1712 => "0011110010110000000100",
			1713 => "1111111001101101000001",
			1714 => "0000001000100100001000",
			1715 => "0001011000000000000100",
			1716 => "1111111001101101000001",
			1717 => "0000010001101101000001",
			1718 => "1111111001101101000001",
			1719 => "0000011001100000010000",
			1720 => "0011100011101000001000",
			1721 => "0001111100010000000100",
			1722 => "0000000001101101000001",
			1723 => "1111111001101101000001",
			1724 => "0000000101101000000100",
			1725 => "1111111001101101000001",
			1726 => "0000000001101101000001",
			1727 => "0001011000100000011000",
			1728 => "0010010110101100010100",
			1729 => "0011110010000100000100",
			1730 => "0000010001101101000001",
			1731 => "0000001010111000001000",
			1732 => "0010001111001000000100",
			1733 => "1111111001101101000001",
			1734 => "0000001001101101000001",
			1735 => "0011001001000100000100",
			1736 => "0000001001101101000001",
			1737 => "0000010001101101000001",
			1738 => "1111111001101101000001",
			1739 => "0010101100001100001000",
			1740 => "0001111001011000000100",
			1741 => "0000000001101101000001",
			1742 => "1111111001101101000001",
			1743 => "0000010001101101000001",
			1744 => "0001101010001000010100",
			1745 => "0000011000011000010000",
			1746 => "0011011010100100000100",
			1747 => "0000000001101111010101",
			1748 => "0001011011111000001000",
			1749 => "0000000100001000000100",
			1750 => "0000000001101111010101",
			1751 => "0000000001101111010101",
			1752 => "0000000001101111010101",
			1753 => "1111111001101111010101",
			1754 => "0011111110101100001100",
			1755 => "0010111100101000001000",
			1756 => "0000001011001000000100",
			1757 => "0000000001101111010101",
			1758 => "0000001001101111010101",
			1759 => "0000000001101111010101",
			1760 => "0000001101011100001100",
			1761 => "0001001100101000001000",
			1762 => "0001111111101000000100",
			1763 => "0000000001101111010101",
			1764 => "0000000001101111010101",
			1765 => "1111111001101111010101",
			1766 => "0001111010011100010100",
			1767 => "0010001001000100001000",
			1768 => "0000001111010000000100",
			1769 => "0000000001101111010101",
			1770 => "0000000001101111010101",
			1771 => "0001011001010100000100",
			1772 => "0000000001101111010101",
			1773 => "0001011011111000000100",
			1774 => "0000000001101111010101",
			1775 => "0000000001101111010101",
			1776 => "0001000110101100000100",
			1777 => "0000000001101111010101",
			1778 => "0000001000001100000100",
			1779 => "0000000001101111010101",
			1780 => "0000000001101111010101",
			1781 => "0010001111001000100100",
			1782 => "0011000011010000011000",
			1783 => "0011011011101100001000",
			1784 => "0000011001100000000100",
			1785 => "1111111001110001111001",
			1786 => "0000000001110001111001",
			1787 => "0001111001010000001000",
			1788 => "0000000100011000000100",
			1789 => "0000000001110001111001",
			1790 => "0000001001110001111001",
			1791 => "0011110111001100000100",
			1792 => "1111111001110001111001",
			1793 => "0000000001110001111001",
			1794 => "0010011001001000001000",
			1795 => "0010101101001000000100",
			1796 => "0000000001110001111001",
			1797 => "0000001001110001111001",
			1798 => "1111111001110001111001",
			1799 => "0001011000000000000100",
			1800 => "1111111001110001111001",
			1801 => "0011000101010100001100",
			1802 => "0000001101001100000100",
			1803 => "0000000001110001111001",
			1804 => "0001100100100000000100",
			1805 => "0000001001110001111001",
			1806 => "0000000001110001111001",
			1807 => "0001011011111000001100",
			1808 => "0010111100101000000100",
			1809 => "0000000001110001111001",
			1810 => "0000111101001000000100",
			1811 => "0000000001110001111001",
			1812 => "1111111001110001111001",
			1813 => "0001011100101100000100",
			1814 => "0000001001110001111001",
			1815 => "0000010110001100001000",
			1816 => "0010000011100100000100",
			1817 => "1111111001110001111001",
			1818 => "0000000001110001111001",
			1819 => "0010000011100100000100",
			1820 => "0000000001110001111001",
			1821 => "0000000001110001111001",
			1822 => "0010100000111100101100",
			1823 => "0010100011000100101000",
			1824 => "0011010011000000100100",
			1825 => "0000101110101000011100",
			1826 => "0010101111101000010000",
			1827 => "0011011001001000001000",
			1828 => "0011010011010000000100",
			1829 => "0000000001110011111101",
			1830 => "0000000001110011111101",
			1831 => "0001011100010000000100",
			1832 => "0000000001110011111101",
			1833 => "1111111001110011111101",
			1834 => "0000111100010000000100",
			1835 => "0000001001110011111101",
			1836 => "0000100010100100000100",
			1837 => "0000000001110011111101",
			1838 => "0000000001110011111101",
			1839 => "0001100000100100000100",
			1840 => "0000001001110011111101",
			1841 => "0000000001110011111101",
			1842 => "1111111001110011111101",
			1843 => "1111111001110011111101",
			1844 => "0001011100011100001000",
			1845 => "0011101101100100000100",
			1846 => "0000000001110011111101",
			1847 => "0000001001110011111101",
			1848 => "0010101100001100000100",
			1849 => "1111111001110011111101",
			1850 => "0010111101101000001000",
			1851 => "0010001010000100000100",
			1852 => "0000000001110011111101",
			1853 => "0000000001110011111101",
			1854 => "0000000001110011111101",
			1855 => "0000100000000000110100",
			1856 => "0001101010001000010100",
			1857 => "0011110010110000000100",
			1858 => "1100110001110110100001",
			1859 => "0011100000010100000100",
			1860 => "1101001001110110100001",
			1861 => "0000001011011000001000",
			1862 => "0011101110111100000100",
			1863 => "1100111001110110100001",
			1864 => "1100110001110110100001",
			1865 => "1100110001110110100001",
			1866 => "0000011001100000000100",
			1867 => "1100110001110110100001",
			1868 => "0001100001100000000100",
			1869 => "1101101001110110100001",
			1870 => "0010011000000000010000",
			1871 => "0010011101101000001000",
			1872 => "0001110001010000000100",
			1873 => "1101000001110110100001",
			1874 => "1100110001110110100001",
			1875 => "0001010011000100000100",
			1876 => "1101100001110110100001",
			1877 => "1101000001110110100001",
			1878 => "0000110001001000000100",
			1879 => "1100110001110110100001",
			1880 => "1100111001110110100001",
			1881 => "0001110011110100011000",
			1882 => "0010000101101100000100",
			1883 => "1100110001110110100001",
			1884 => "0000100101101000001100",
			1885 => "0011000101010100000100",
			1886 => "1110010001110110100001",
			1887 => "0000011110011000000100",
			1888 => "1101000001110110100001",
			1889 => "1101110001110110100001",
			1890 => "0001001000000100000100",
			1891 => "1110110001110110100001",
			1892 => "1101110001110110100001",
			1893 => "0001011011000000000100",
			1894 => "1101000001110110100001",
			1895 => "1100110001110110100001",
			1896 => "0000011001100000100000",
			1897 => "0011110011101100001000",
			1898 => "0001100001001100000100",
			1899 => "0000000001111001100101",
			1900 => "0000000001111001100101",
			1901 => "0011101100000100010100",
			1902 => "0000111111011000001100",
			1903 => "0001111101001000001000",
			1904 => "0000111101101000000100",
			1905 => "0000000001111001100101",
			1906 => "0000000001111001100101",
			1907 => "0000000001111001100101",
			1908 => "0001111001011000000100",
			1909 => "0000000001111001100101",
			1910 => "0000000001111001100101",
			1911 => "0000000001111001100101",
			1912 => "0001111100011100110000",
			1913 => "0010100000111100011100",
			1914 => "0001011000100000010100",
			1915 => "0011010011000000010000",
			1916 => "0010001001000100001000",
			1917 => "0010111011101100000100",
			1918 => "0000000001111001100101",
			1919 => "0000000001111001100101",
			1920 => "0001101110000100000100",
			1921 => "0000000001111001100101",
			1922 => "0000000001111001100101",
			1923 => "0000000001111001100101",
			1924 => "0001110001010000000100",
			1925 => "0000000001111001100101",
			1926 => "0000000001111001100101",
			1927 => "0010011100000000001000",
			1928 => "0000010110001100000100",
			1929 => "0000000001111001100101",
			1930 => "0000000001111001100101",
			1931 => "0011000101111000001000",
			1932 => "0001011010110100000100",
			1933 => "0000000001111001100101",
			1934 => "0000000001111001100101",
			1935 => "0000000001111001100101",
			1936 => "0011000011000000001000",
			1937 => "0011110100111100000100",
			1938 => "0000000001111001100101",
			1939 => "0000000001111001100101",
			1940 => "0001101100111100000100",
			1941 => "0000000001111001100101",
			1942 => "0000111111101000000100",
			1943 => "0000000001111001100101",
			1944 => "0000000001111001100101",
			1945 => "0000001110110000111100",
			1946 => "0010001111001000010100",
			1947 => "0010111011101100010000",
			1948 => "0011001011101100000100",
			1949 => "0000000001111100010001",
			1950 => "0010110110001100000100",
			1951 => "0000000001111100010001",
			1952 => "0000010001110000000100",
			1953 => "0000000001111100010001",
			1954 => "0000000001111100010001",
			1955 => "0000000001111100010001",
			1956 => "0011000101101100011000",
			1957 => "0010111001001000010100",
			1958 => "0000000100110100001000",
			1959 => "0000110011000000000100",
			1960 => "0000000001111100010001",
			1961 => "0000000001111100010001",
			1962 => "0001011001011000001000",
			1963 => "0001011101001000000100",
			1964 => "0000000001111100010001",
			1965 => "0000000001111100010001",
			1966 => "0000000001111100010001",
			1967 => "0000000001111100010001",
			1968 => "0000000100010100001000",
			1969 => "0011110101111100000100",
			1970 => "0000000001111100010001",
			1971 => "0000000001111100010001",
			1972 => "0001101010101100000100",
			1973 => "0000000001111100010001",
			1974 => "0000000001111100010001",
			1975 => "0010010110101100011000",
			1976 => "0000010111100100000100",
			1977 => "0000000001111100010001",
			1978 => "0011100101001100010000",
			1979 => "0010001010000100001000",
			1980 => "0011100011101000000100",
			1981 => "0000000001111100010001",
			1982 => "0000000001111100010001",
			1983 => "0000010101011100000100",
			1984 => "0000000001111100010001",
			1985 => "0000000001111100010001",
			1986 => "0000000001111100010001",
			1987 => "0000000001111100010001",
			1988 => "0011111010101100010000",
			1989 => "0011110010110000000100",
			1990 => "1111111001111110010101",
			1991 => "0000001000100100001000",
			1992 => "0011011010100100000100",
			1993 => "1111111001111110010101",
			1994 => "0000001001111110010101",
			1995 => "1111111001111110010101",
			1996 => "0010001111111100000100",
			1997 => "1111111001111110010101",
			1998 => "0011010011000000101000",
			1999 => "0000101111001100010100",
			2000 => "0000101010010100010000",
			2001 => "0010001111001000001000",
			2002 => "0010111011101100000100",
			2003 => "0000010001111110010101",
			2004 => "1111111001111110010101",
			2005 => "0011000101101100000100",
			2006 => "0000001001111110010101",
			2007 => "0000000001111110010101",
			2008 => "0000000001111110010101",
			2009 => "0010000011001000001100",
			2010 => "0011000101011100001000",
			2011 => "0010101111101000000100",
			2012 => "0000001001111110010101",
			2013 => "0000001001111110010101",
			2014 => "0000000001111110010101",
			2015 => "0000111111101000000100",
			2016 => "0000001001111110010101",
			2017 => "0000001001111110010101",
			2018 => "0000010101010100000100",
			2019 => "0000000001111110010101",
			2020 => "1111111001111110010101",
			2021 => "0001011000000000011000",
			2022 => "0001111100010000001000",
			2023 => "0000110011001000000100",
			2024 => "0000000010000001101001",
			2025 => "0000000010000001101001",
			2026 => "0000110011000000001000",
			2027 => "0000111101101000000100",
			2028 => "0000000010000001101001",
			2029 => "0000000010000001101001",
			2030 => "0011101000110100000100",
			2031 => "0000000010000001101001",
			2032 => "0000000010000001101001",
			2033 => "0011000101010100100100",
			2034 => "0000101100001000011000",
			2035 => "0001111000101000010000",
			2036 => "0010001001000100001000",
			2037 => "0000001100111100000100",
			2038 => "0000000010000001101001",
			2039 => "0000000010000001101001",
			2040 => "0001001010000100000100",
			2041 => "0000000010000001101001",
			2042 => "0000000010000001101001",
			2043 => "0001001001000100000100",
			2044 => "0000000010000001101001",
			2045 => "0000000010000001101001",
			2046 => "0000010111100100000100",
			2047 => "0000000010000001101001",
			2048 => "0001101010101100000100",
			2049 => "0000000010000001101001",
			2050 => "0000000010000001101001",
			2051 => "0011011100101000010000",
			2052 => "0000010110001100001000",
			2053 => "0010110011010000000100",
			2054 => "0000000010000001101001",
			2055 => "0000000010000001101001",
			2056 => "0000001010010100000100",
			2057 => "0000000010000001101001",
			2058 => "0000000010000001101001",
			2059 => "0010111001001000001000",
			2060 => "0010100011000100000100",
			2061 => "0000000010000001101001",
			2062 => "0000000010000001101001",
			2063 => "0011000110000000001000",
			2064 => "0000100101101000000100",
			2065 => "0000000010000001101001",
			2066 => "0000000010000001101001",
			2067 => "0000010111011100001000",
			2068 => "0001010011000100000100",
			2069 => "0000000010000001101001",
			2070 => "0000000010000001101001",
			2071 => "0011101010001000000100",
			2072 => "0000000010000001101001",
			2073 => "0000000010000001101001",
			2074 => "0000100100010100110100",
			2075 => "0011110000000100100000",
			2076 => "0011111010101100010000",
			2077 => "0001100011011000001100",
			2078 => "0011110010110000000100",
			2079 => "0000000010000101001101",
			2080 => "0001011100101100000100",
			2081 => "0000000010000101001101",
			2082 => "0000000010000101001101",
			2083 => "0000000010000101001101",
			2084 => "0010111001001000001100",
			2085 => "0000010011110000001000",
			2086 => "0000001010000000000100",
			2087 => "0000000010000101001101",
			2088 => "0000000010000101001101",
			2089 => "0000000010000101001101",
			2090 => "0000000010000101001101",
			2091 => "0010110101101100001100",
			2092 => "0001000101011100001000",
			2093 => "0001110001010000000100",
			2094 => "0000000010000101001101",
			2095 => "0000000010000101001101",
			2096 => "0000000010000101001101",
			2097 => "0000000100010100000100",
			2098 => "0000000010000101001101",
			2099 => "0000000010000101001101",
			2100 => "0011110101100100011100",
			2101 => "0001100001111000001000",
			2102 => "0000000101101000000100",
			2103 => "0000000010000101001101",
			2104 => "0000000010000101001101",
			2105 => "0001000110000000000100",
			2106 => "0000000010000101001101",
			2107 => "0001011100101100000100",
			2108 => "0000000010000101001101",
			2109 => "0000011101000000000100",
			2110 => "0000000010000101001101",
			2111 => "0000010111011100000100",
			2112 => "0000000010000101001101",
			2113 => "0000000010000101001101",
			2114 => "0000101010010000011100",
			2115 => "0001011011111000001100",
			2116 => "0001000101111000001000",
			2117 => "0001111000101000000100",
			2118 => "0000000010000101001101",
			2119 => "0000000010000101001101",
			2120 => "0000000010000101001101",
			2121 => "0011010011000000001100",
			2122 => "0001010011000100000100",
			2123 => "0000000010000101001101",
			2124 => "0010011000000000000100",
			2125 => "0000000010000101001101",
			2126 => "0000000010000101001101",
			2127 => "0000000010000101001101",
			2128 => "0001111001000000000100",
			2129 => "0000000010000101001101",
			2130 => "0000000010000101001101",
			2131 => "0010001111001000101000",
			2132 => "0011000011010000011100",
			2133 => "0001101110010000001100",
			2134 => "0001111000111000000100",
			2135 => "1111111010001000000001",
			2136 => "0001010011001000000100",
			2137 => "0000000010001000000001",
			2138 => "0000001010001000000001",
			2139 => "0000001111010000001100",
			2140 => "0001011111101000001000",
			2141 => "0001111100010000000100",
			2142 => "0000000010001000000001",
			2143 => "1111111010001000000001",
			2144 => "0000000010001000000001",
			2145 => "0000000010001000000001",
			2146 => "0010011001001000001000",
			2147 => "0010101101001000000100",
			2148 => "0000000010001000000001",
			2149 => "0000001010001000000001",
			2150 => "1111111010001000000001",
			2151 => "0001011000000000000100",
			2152 => "1111111010001000000001",
			2153 => "0011000101010100001100",
			2154 => "0000001101001100000100",
			2155 => "0000000010001000000001",
			2156 => "0001100100100000000100",
			2157 => "0000001010001000000001",
			2158 => "0000000010001000000001",
			2159 => "0001011011111000010000",
			2160 => "0000001010111000001100",
			2161 => "0000101100010100000100",
			2162 => "0000001010001000000001",
			2163 => "0000111100010000000100",
			2164 => "0000000010001000000001",
			2165 => "1111111010001000000001",
			2166 => "0000000010001000000001",
			2167 => "0001011100101100000100",
			2168 => "0000001010001000000001",
			2169 => "0000010110001100001000",
			2170 => "0010000011100100000100",
			2171 => "1111111010001000000001",
			2172 => "0000000010001000000001",
			2173 => "0011011001001000000100",
			2174 => "0000001010001000000001",
			2175 => "0000000010001000000001",
			2176 => "0000000110101000100000",
			2177 => "0011110100010000001100",
			2178 => "0011110010110000000100",
			2179 => "1111111010001010100101",
			2180 => "0010000000110000000100",
			2181 => "1111111010001010100101",
			2182 => "0000001010001010100101",
			2183 => "0011110100111000000100",
			2184 => "0000010010001010100101",
			2185 => "0001111000101000001000",
			2186 => "0010011001000100000100",
			2187 => "1111111010001010100101",
			2188 => "0000001010001010100101",
			2189 => "0000010011010000000100",
			2190 => "1111111010001010100101",
			2191 => "0000000010001010100101",
			2192 => "0010000101101100000100",
			2193 => "1111111010001010100101",
			2194 => "0011010011000000101000",
			2195 => "0000001010111000010100",
			2196 => "0000110011000100010000",
			2197 => "0010100011000100001000",
			2198 => "0010001111001000000100",
			2199 => "0000000010001010100101",
			2200 => "0000001010001010100101",
			2201 => "0000010011010000000100",
			2202 => "1111111010001010100101",
			2203 => "0000000010001010100101",
			2204 => "0000010010001010100101",
			2205 => "0011100101001100010000",
			2206 => "0010000011001000001000",
			2207 => "0001010001010000000100",
			2208 => "0000001010001010100101",
			2209 => "0000001010001010100101",
			2210 => "0001011011000000000100",
			2211 => "0000010010001010100101",
			2212 => "0000001010001010100101",
			2213 => "0000000010001010100101",
			2214 => "0000010101010100000100",
			2215 => "0000000010001010100101",
			2216 => "1111111010001010100101",
			2217 => "0011110010110000000100",
			2218 => "1111111010001100000001",
			2219 => "0011010011000000101000",
			2220 => "0011011010000100100000",
			2221 => "0011011101101000011100",
			2222 => "0000010011110000001100",
			2223 => "0010110011010000001000",
			2224 => "0010000101101100000100",
			2225 => "1111111010001100000001",
			2226 => "0000000010001100000001",
			2227 => "1111111010001100000001",
			2228 => "0001000011000000001000",
			2229 => "0001001001001000000100",
			2230 => "0000000010001100000001",
			2231 => "0000001010001100000001",
			2232 => "0001111100101100000100",
			2233 => "0000000010001100000001",
			2234 => "0000000010001100000001",
			2235 => "1111111010001100000001",
			2236 => "0001111001000000000100",
			2237 => "0000000010001100000001",
			2238 => "0000001010001100000001",
			2239 => "1111111010001100000001",
			2240 => "0011111010101100001100",
			2241 => "0011110010110000000100",
			2242 => "1111111010001110001101",
			2243 => "0001111100110000000100",
			2244 => "0000000010001110001101",
			2245 => "1111111010001110001101",
			2246 => "0010000101101100001000",
			2247 => "0011111101010000000100",
			2248 => "0000001010001110001101",
			2249 => "1111111010001110001101",
			2250 => "0001110011110100101100",
			2251 => "0000100100010100010100",
			2252 => "0010001000000000010000",
			2253 => "0000011101000000001000",
			2254 => "0000001100010100000100",
			2255 => "0000010010001110001101",
			2256 => "1111111010001110001101",
			2257 => "0011010101101100000100",
			2258 => "0000010010001110001101",
			2259 => "0000000010001110001101",
			2260 => "1111111010001110001101",
			2261 => "0010001010000100001100",
			2262 => "0010111010100100000100",
			2263 => "0000010010001110001101",
			2264 => "0011010111011100000100",
			2265 => "0000000010001110001101",
			2266 => "1111111010001110001101",
			2267 => "0001101000010100000100",
			2268 => "0000011010001110001101",
			2269 => "0010001000000000000100",
			2270 => "0000010010001110001101",
			2271 => "0000000010001110001101",
			2272 => "0001011011000000000100",
			2273 => "0000000010001110001101",
			2274 => "1111111010001110001101",
			2275 => "0011011100101000111100",
			2276 => "0010110101010100101000",
			2277 => "0000010011110000011000",
			2278 => "0010111010100100010100",
			2279 => "0010000101101100000100",
			2280 => "1111111010010001101001",
			2281 => "0001000101010100001000",
			2282 => "0001100000001100000100",
			2283 => "1111111010010001101001",
			2284 => "0000000010010001101001",
			2285 => "0010101000111000000100",
			2286 => "0000000010010001101001",
			2287 => "0000001010010001101001",
			2288 => "1111111010010001101001",
			2289 => "0011101110100100001000",
			2290 => "0000001101001100000100",
			2291 => "1111111010010001101001",
			2292 => "0000001010010001101001",
			2293 => "0000111001010100000100",
			2294 => "1111111010010001101001",
			2295 => "0000000010010001101001",
			2296 => "0010100001011100001100",
			2297 => "0011111110101100001000",
			2298 => "0011100011010100000100",
			2299 => "1111111010010001101001",
			2300 => "0000000010010001101001",
			2301 => "1111111010010001101001",
			2302 => "0001111011111000000100",
			2303 => "0000000010010001101001",
			2304 => "0000000010010001101001",
			2305 => "0011011001001000001100",
			2306 => "0001010011000100001000",
			2307 => "0010101101001000000100",
			2308 => "0000000010010001101001",
			2309 => "0000001010010001101001",
			2310 => "0000000010010001101001",
			2311 => "0010011000000100001100",
			2312 => "0000111111101000001000",
			2313 => "0001011001010000000100",
			2314 => "0000000010010001101001",
			2315 => "1111111010010001101001",
			2316 => "0000000010010001101001",
			2317 => "0011101111010100000100",
			2318 => "1111111010010001101001",
			2319 => "0000000100010100001000",
			2320 => "0010001000111000000100",
			2321 => "0000001010010001101001",
			2322 => "0000000010010001101001",
			2323 => "0000001011001100001000",
			2324 => "0011110100011000000100",
			2325 => "0000000010010001101001",
			2326 => "1111111010010001101001",
			2327 => "0011110101100100000100",
			2328 => "0000001010010001101001",
			2329 => "0000000010010001101001",
			2330 => "0010100000111100111100",
			2331 => "0001010001001000111000",
			2332 => "0000001010111000101000",
			2333 => "0011110000100100011100",
			2334 => "0001001100000000010000",
			2335 => "0001011100101100001000",
			2336 => "0000100100010100000100",
			2337 => "0000000010010011111101",
			2338 => "0000000010010011111101",
			2339 => "0001101110010000000100",
			2340 => "0000000010010011111101",
			2341 => "1111111010010011111101",
			2342 => "0010000011100100001000",
			2343 => "0001001100110000000100",
			2344 => "0000000010010011111101",
			2345 => "0000000010010011111101",
			2346 => "0000000010010011111101",
			2347 => "0010101111101000000100",
			2348 => "0000000010010011111101",
			2349 => "0000100111111000000100",
			2350 => "0000000010010011111101",
			2351 => "0000000010010011111101",
			2352 => "0011011101101000001100",
			2353 => "0010001010000100001000",
			2354 => "0000100101010000000100",
			2355 => "0000000010010011111101",
			2356 => "0000000010010011111101",
			2357 => "0000001010010011111101",
			2358 => "0000000010010011111101",
			2359 => "0000000010010011111101",
			2360 => "0001101110000100001100",
			2361 => "0000000110111100000100",
			2362 => "0000000010010011111101",
			2363 => "0000010111011100000100",
			2364 => "0000000010010011111101",
			2365 => "0000000010010011111101",
			2366 => "0000000010010011111101",
			2367 => "0011100001100001001100",
			2368 => "0001001100000000101000",
			2369 => "0001000011001000100100",
			2370 => "0011011101101000100000",
			2371 => "0000011001100000010000",
			2372 => "0011110011101100001000",
			2373 => "0000111100010000000100",
			2374 => "0000000010010110111001",
			2375 => "0000000010010110111001",
			2376 => "0011100011101000000100",
			2377 => "0000000010010110111001",
			2378 => "0000000010010110111001",
			2379 => "0011100100101000001000",
			2380 => "0001101100000100000100",
			2381 => "0000000010010110111001",
			2382 => "0000000010010110111001",
			2383 => "0011100010110100000100",
			2384 => "0000000010010110111001",
			2385 => "0000000010010110111001",
			2386 => "0000000010010110111001",
			2387 => "0000000010010110111001",
			2388 => "0010000011100100010100",
			2389 => "0000100010100100001000",
			2390 => "0001011011000000000100",
			2391 => "0000000010010110111001",
			2392 => "0000000010010110111001",
			2393 => "0010010011000000001000",
			2394 => "0000111011111000000100",
			2395 => "0000000010010110111001",
			2396 => "0000000010010110111001",
			2397 => "0000000010010110111001",
			2398 => "0011011010000100000100",
			2399 => "0000000010010110111001",
			2400 => "0010001100110000000100",
			2401 => "0000000010010110111001",
			2402 => "0000001011001100000100",
			2403 => "0000000010010110111001",
			2404 => "0000000010010110111001",
			2405 => "0000011100101000001100",
			2406 => "0011110100110100000100",
			2407 => "0000000010010110111001",
			2408 => "0000101101011000000100",
			2409 => "0000000010010110111001",
			2410 => "0000000010010110111001",
			2411 => "0000111001010000000100",
			2412 => "0000000010010110111001",
			2413 => "0000000010010110111001",
			2414 => "0010101101001000001000",
			2415 => "0000100101101000000100",
			2416 => "0000000010011001101101",
			2417 => "0000000010011001101101",
			2418 => "0001011001010000011100",
			2419 => "0010001001000100010000",
			2420 => "0001011000000000001000",
			2421 => "0011100010110100000100",
			2422 => "0000000010011001101101",
			2423 => "0000000010011001101101",
			2424 => "0000001001101000000100",
			2425 => "0000000010011001101101",
			2426 => "0000000010011001101101",
			2427 => "0000111001010000001000",
			2428 => "0000001011011000000100",
			2429 => "0000000010011001101101",
			2430 => "0000000010011001101101",
			2431 => "0000000010011001101101",
			2432 => "0011011100101000011000",
			2433 => "0000010110001100010000",
			2434 => "0011000101010100001100",
			2435 => "0011111011000100001000",
			2436 => "0011110110011000000100",
			2437 => "0000000010011001101101",
			2438 => "0000000010011001101101",
			2439 => "0000000010011001101101",
			2440 => "0000000010011001101101",
			2441 => "0011101100011000000100",
			2442 => "0000000010011001101101",
			2443 => "0000000010011001101101",
			2444 => "0000010111011100011000",
			2445 => "0001010011000100001000",
			2446 => "0001011011111000000100",
			2447 => "0000000010011001101101",
			2448 => "0000000010011001101101",
			2449 => "0010101100001100001000",
			2450 => "0010000011001000000100",
			2451 => "0000000010011001101101",
			2452 => "0000000010011001101101",
			2453 => "0001110011110100000100",
			2454 => "0000000010011001101101",
			2455 => "0000000010011001101101",
			2456 => "0011011101101000000100",
			2457 => "0000000010011001101101",
			2458 => "0000000010011001101101",
			2459 => "0001110011110101010100",
			2460 => "0001101110001000110000",
			2461 => "0011110000000100011100",
			2462 => "0010111001001000011000",
			2463 => "0001101010001000001100",
			2464 => "0001100011011000001000",
			2465 => "0001111100010000000100",
			2466 => "0000000010011100110001",
			2467 => "0000000010011100110001",
			2468 => "0000000010011100110001",
			2469 => "0000010011110000001000",
			2470 => "0000000111011000000100",
			2471 => "0000000010011100110001",
			2472 => "0000000010011100110001",
			2473 => "0000001010011100110001",
			2474 => "0000000010011100110001",
			2475 => "0011001010100100001000",
			2476 => "0000001011001100000100",
			2477 => "0000000010011100110001",
			2478 => "0000000010011100110001",
			2479 => "0001001001000100000100",
			2480 => "0000000010011100110001",
			2481 => "0001001000111000000100",
			2482 => "1111111010011100110001",
			2483 => "0000000010011100110001",
			2484 => "0001101100111000001000",
			2485 => "0000001101111000000100",
			2486 => "0000000010011100110001",
			2487 => "0000001010011100110001",
			2488 => "0011100100101000001100",
			2489 => "0001101000010100000100",
			2490 => "0000000010011100110001",
			2491 => "0001111001010000000100",
			2492 => "0000000010011100110001",
			2493 => "1111111010011100110001",
			2494 => "0001001101001000001100",
			2495 => "0001001000111000001000",
			2496 => "0001001111011000000100",
			2497 => "0000000010011100110001",
			2498 => "0000000010011100110001",
			2499 => "0000000010011100110001",
			2500 => "0000000010011100110001",
			2501 => "0011000011000000000100",
			2502 => "1111111010011100110001",
			2503 => "0000001010010000000100",
			2504 => "0000000010011100110001",
			2505 => "0000101001101000000100",
			2506 => "0000000010011100110001",
			2507 => "0000000010011100110001",
			2508 => "0000011101000000110100",
			2509 => "0010111010100100100000",
			2510 => "0000001110110000011000",
			2511 => "0001101110010000010000",
			2512 => "0000110011001000000100",
			2513 => "0000000010100000011101",
			2514 => "0000000100011000000100",
			2515 => "0000000010100000011101",
			2516 => "0000010001110000000100",
			2517 => "0000000010100000011101",
			2518 => "0000000010100000011101",
			2519 => "0010001001000100000100",
			2520 => "0000000010100000011101",
			2521 => "0000000010100000011101",
			2522 => "0000010111100100000100",
			2523 => "0000000010100000011101",
			2524 => "0000000010100000011101",
			2525 => "0011100100101000001100",
			2526 => "0011000011010000001000",
			2527 => "0001011100110000000100",
			2528 => "0000000010100000011101",
			2529 => "0000000010100000011101",
			2530 => "1111111010100000011101",
			2531 => "0011000101010100000100",
			2532 => "0000000010100000011101",
			2533 => "0000000010100000011101",
			2534 => "0010111001001000011000",
			2535 => "0011000101101100010100",
			2536 => "0000111001010100001100",
			2537 => "0011110101111100001000",
			2538 => "0001011000000000000100",
			2539 => "0000000010100000011101",
			2540 => "0000000010100000011101",
			2541 => "0000000010100000011101",
			2542 => "0010110101011100000100",
			2543 => "0000000010100000011101",
			2544 => "0000000010100000011101",
			2545 => "0000000010100000011101",
			2546 => "0010011000000100001000",
			2547 => "0001001001000100000100",
			2548 => "0000000010100000011101",
			2549 => "0000000010100000011101",
			2550 => "0011111001111000010000",
			2551 => "0000011010100100001100",
			2552 => "0010001111011000000100",
			2553 => "0000000010100000011101",
			2554 => "0001011111111000000100",
			2555 => "0000000010100000011101",
			2556 => "0000000010100000011101",
			2557 => "0000000010100000011101",
			2558 => "0010010110101100010000",
			2559 => "0001010011000100001000",
			2560 => "0001011011111000000100",
			2561 => "0000000010100000011101",
			2562 => "0000000010100000011101",
			2563 => "0011001101101000000100",
			2564 => "0000000010100000011101",
			2565 => "0000000010100000011101",
			2566 => "0000000010100000011101",
			2567 => "0001110011110101001100",
			2568 => "0011111010101100011000",
			2569 => "0000011000011000001100",
			2570 => "0010111010100100001000",
			2571 => "0000110011001000000100",
			2572 => "0000000010100010111001",
			2573 => "0000000010100010111001",
			2574 => "0000000010100010111001",
			2575 => "0000110011000000001000",
			2576 => "0000111001000100000100",
			2577 => "0000000010100010111001",
			2578 => "0000000010100010111001",
			2579 => "0000000010100010111001",
			2580 => "0011110101100100100000",
			2581 => "0000001110110000010100",
			2582 => "0000001111001100010000",
			2583 => "0011000101101100001000",
			2584 => "0000011001100000000100",
			2585 => "0000000010100010111001",
			2586 => "0000000010100010111001",
			2587 => "0011100110111000000100",
			2588 => "0000000010100010111001",
			2589 => "0000000010100010111001",
			2590 => "0000000010100010111001",
			2591 => "0000011101000000001000",
			2592 => "0011101111010100000100",
			2593 => "0000000010100010111001",
			2594 => "0000000010100010111001",
			2595 => "0000000010100010111001",
			2596 => "0000001000110000010000",
			2597 => "0011110000101100000100",
			2598 => "0000000010100010111001",
			2599 => "0001001001000100000100",
			2600 => "0000000010100010111001",
			2601 => "0010101011111000000100",
			2602 => "0000000010100010111001",
			2603 => "0000000010100010111001",
			2604 => "0000000010100010111001",
			2605 => "0000000010100010111001",
			2606 => "0000101111001101010000",
			2607 => "0011111011110100111000",
			2608 => "0011110110011000101100",
			2609 => "0001101100000100011000",
			2610 => "0001101010001000001100",
			2611 => "0001111100110000001000",
			2612 => "0001111100010000000100",
			2613 => "0000000010100110000101",
			2614 => "0000000010100110000101",
			2615 => "0000000010100110000101",
			2616 => "0011000101101100001000",
			2617 => "0000011001100000000100",
			2618 => "0000000010100110000101",
			2619 => "0000000010100110000101",
			2620 => "0000000010100110000101",
			2621 => "0001010001101000010000",
			2622 => "0011101100011000001000",
			2623 => "0001001111011000000100",
			2624 => "0000000010100110000101",
			2625 => "0000000010100110000101",
			2626 => "0001111011111000000100",
			2627 => "0000000010100110000101",
			2628 => "1111111010100110000101",
			2629 => "0000000010100110000101",
			2630 => "0001001010000100000100",
			2631 => "0000000010100110000101",
			2632 => "0011100011101000000100",
			2633 => "0000000010100110000101",
			2634 => "0000000010100110000101",
			2635 => "0000100000000000000100",
			2636 => "1111111010100110000101",
			2637 => "0010000011100100001100",
			2638 => "0000001001101000001000",
			2639 => "0001101101010000000100",
			2640 => "0000000010100110000101",
			2641 => "0000000010100110000101",
			2642 => "0000000010100110000101",
			2643 => "0001100111010000000100",
			2644 => "0000000010100110000101",
			2645 => "0000000010100110000101",
			2646 => "0011000101111000010100",
			2647 => "0010000000110000001100",
			2648 => "0010010101101100001000",
			2649 => "0010001111111100000100",
			2650 => "0000000010100110000101",
			2651 => "0000000010100110000101",
			2652 => "0000000010100110000101",
			2653 => "0001110011110100000100",
			2654 => "0000000010100110000101",
			2655 => "0000000010100110000101",
			2656 => "0000000010100110000101",
			2657 => "0010001000000001011100",
			2658 => "0010001111001000100100",
			2659 => "0000101011001100011000",
			2660 => "0011110011101100001000",
			2661 => "0001101110111100000100",
			2662 => "0000000010101001101001",
			2663 => "0000000010101001101001",
			2664 => "0010101100010000001100",
			2665 => "0001101010001000000100",
			2666 => "0000000010101001101001",
			2667 => "0001100001100000000100",
			2668 => "0000000010101001101001",
			2669 => "0000000010101001101001",
			2670 => "0000000010101001101001",
			2671 => "0011101110010000001000",
			2672 => "0000010111100100000100",
			2673 => "0000000010101001101001",
			2674 => "0000000010101001101001",
			2675 => "0000000010101001101001",
			2676 => "0011000101010100001100",
			2677 => "0001011000000100000100",
			2678 => "0000000010101001101001",
			2679 => "0011110010110000000100",
			2680 => "0000000010101001101001",
			2681 => "0000000010101001101001",
			2682 => "0010001111011000011000",
			2683 => "0001001100000000010000",
			2684 => "0011011001001000001000",
			2685 => "0001100111101000000100",
			2686 => "0000000010101001101001",
			2687 => "0000000010101001101001",
			2688 => "0011011001000100000100",
			2689 => "0000000010101001101001",
			2690 => "0000000010101001101001",
			2691 => "0000000110010100000100",
			2692 => "0000000010101001101001",
			2693 => "0000000010101001101001",
			2694 => "0011111101010000000100",
			2695 => "0000000010101001101001",
			2696 => "0010111001001000001000",
			2697 => "0001111001011000000100",
			2698 => "0000000010101001101001",
			2699 => "0000000010101001101001",
			2700 => "0001101101010000000100",
			2701 => "0000000010101001101001",
			2702 => "0000000010101001101001",
			2703 => "0001000011000000001000",
			2704 => "0010001100110000000100",
			2705 => "0000000010101001101001",
			2706 => "0000000010101001101001",
			2707 => "0010001001010100001000",
			2708 => "0000111010100000000100",
			2709 => "0000000010101001101001",
			2710 => "0000000010101001101001",
			2711 => "0011101010001000000100",
			2712 => "0000000010101001101001",
			2713 => "0000000010101001101001",
			2714 => "0001010011001000000100",
			2715 => "1111111010101011111101",
			2716 => "0010111011101100001100",
			2717 => "0010001111111100000100",
			2718 => "0000000010101011111101",
			2719 => "0001100010000100000100",
			2720 => "0000001010101011111101",
			2721 => "0000000010101011111101",
			2722 => "0010001111001000011000",
			2723 => "0011110100110100010000",
			2724 => "0001011000111000001100",
			2725 => "0001100101000000001000",
			2726 => "0000000101100100000100",
			2727 => "0000000010101011111101",
			2728 => "0000000010101011111101",
			2729 => "0000000010101011111101",
			2730 => "1111111010101011111101",
			2731 => "0011100001100000000100",
			2732 => "0000000010101011111101",
			2733 => "0000000010101011111101",
			2734 => "0011000101010100001100",
			2735 => "0010101000101000001000",
			2736 => "0000110011100100000100",
			2737 => "0000001010101011111101",
			2738 => "0000000010101011111101",
			2739 => "0000001010101011111101",
			2740 => "0010100000111100001100",
			2741 => "0010100011000100001000",
			2742 => "0011111100111100000100",
			2743 => "0000000010101011111101",
			2744 => "0000000010101011111101",
			2745 => "1111111010101011111101",
			2746 => "0011101110010000001000",
			2747 => "0000001100100100000100",
			2748 => "0000000010101011111101",
			2749 => "0000001010101011111101",
			2750 => "0000000010101011111101",
			2751 => "0010001000000001100100",
			2752 => "0001110110011101001000",
			2753 => "0011000101010100101000",
			2754 => "0001010011001000001100",
			2755 => "0000110011000000001000",
			2756 => "0000111101101000000100",
			2757 => "0000000010101111100001",
			2758 => "0000000010101111100001",
			2759 => "0000000010101111100001",
			2760 => "0001011001010000010000",
			2761 => "0011110100010000001000",
			2762 => "0000110011000000000100",
			2763 => "0000000010101111100001",
			2764 => "0000000010101111100001",
			2765 => "0010001111111100000100",
			2766 => "0000000010101111100001",
			2767 => "0000000010101111100001",
			2768 => "0001001010000100000100",
			2769 => "0000000010101111100001",
			2770 => "0011101111010100000100",
			2771 => "0000000010101111100001",
			2772 => "0000000010101111100001",
			2773 => "0010001111011000010000",
			2774 => "0001010011000100001000",
			2775 => "0001001100000000000100",
			2776 => "0000000010101111100001",
			2777 => "0000000010101111100001",
			2778 => "0001001100110000000100",
			2779 => "0000000010101111100001",
			2780 => "0000000010101111100001",
			2781 => "0010010011001000001000",
			2782 => "0010010101111000000100",
			2783 => "0000000010101111100001",
			2784 => "0000000010101111100001",
			2785 => "0010100000111100000100",
			2786 => "0000000010101111100001",
			2787 => "0000000010101111100001",
			2788 => "0010101011000000001100",
			2789 => "0011100100111000000100",
			2790 => "0000000010101111100001",
			2791 => "0000001110101000000100",
			2792 => "0000000010101111100001",
			2793 => "0000000010101111100001",
			2794 => "0000111011000000001000",
			2795 => "0010000011001000000100",
			2796 => "0000000010101111100001",
			2797 => "0000000010101111100001",
			2798 => "0011001101101000000100",
			2799 => "0000000010101111100001",
			2800 => "0000000010101111100001",
			2801 => "0000101111001100001000",
			2802 => "0010111001000100000100",
			2803 => "0000000010101111100001",
			2804 => "0000000010101111100001",
			2805 => "0000111001010000000100",
			2806 => "0000000010101111100001",
			2807 => "0000000010101111100001",
			2808 => "0010000101101100000100",
			2809 => "1111111010110001101101",
			2810 => "0000001101011000110100",
			2811 => "0010100000111100100100",
			2812 => "0010100011000100100000",
			2813 => "0011111011010100010000",
			2814 => "0011100001000000001000",
			2815 => "0011010101101100000100",
			2816 => "0000000010110001101101",
			2817 => "1111111010110001101101",
			2818 => "0000001101011100000100",
			2819 => "0000000010110001101101",
			2820 => "0000001010110001101101",
			2821 => "0011010101101100001000",
			2822 => "0001101110000100000100",
			2823 => "1111111010110001101101",
			2824 => "0000000010110001101101",
			2825 => "0001001000000000000100",
			2826 => "0000000010110001101101",
			2827 => "1111111010110001101101",
			2828 => "1111111010110001101101",
			2829 => "0000001100100100000100",
			2830 => "1111111010110001101101",
			2831 => "0000001110110000001000",
			2832 => "0001101010101100000100",
			2833 => "0000001010110001101101",
			2834 => "1111111010110001101101",
			2835 => "0000001010110001101101",
			2836 => "0001111110001100001100",
			2837 => "0010101011000000001000",
			2838 => "0010101111101000000100",
			2839 => "0000000010110001101101",
			2840 => "0000001010110001101101",
			2841 => "0000000010110001101101",
			2842 => "1111111010110001101101",
			2843 => "0010101101001000011100",
			2844 => "0000000100110100000100",
			2845 => "1111111010110100111001",
			2846 => "0001101110010000001000",
			2847 => "0011011011101100000100",
			2848 => "0000000010110100111001",
			2849 => "0000000010110100111001",
			2850 => "0001000111011100001100",
			2851 => "0001111001010000001000",
			2852 => "0001001011101100000100",
			2853 => "0000000010110100111001",
			2854 => "0000000010110100111001",
			2855 => "0000000010110100111001",
			2856 => "1111111010110100111001",
			2857 => "0000111100110000011100",
			2858 => "0000010011010000011000",
			2859 => "0000001010111000010100",
			2860 => "0001110001010000010000",
			2861 => "0000001100100100001000",
			2862 => "0001101111110000000100",
			2863 => "0000000010110100111001",
			2864 => "0000000010110100111001",
			2865 => "0001011100110000000100",
			2866 => "0000000010110100111001",
			2867 => "0000000010110100111001",
			2868 => "1111111010110100111001",
			2869 => "0000001010110100111001",
			2870 => "0000001010110100111001",
			2871 => "0001011011111000010100",
			2872 => "0010110101010100010000",
			2873 => "0011110101100100001000",
			2874 => "0011011110011000000100",
			2875 => "0000000010110100111001",
			2876 => "0000000010110100111001",
			2877 => "0001111100101100000100",
			2878 => "0000000010110100111001",
			2879 => "0000000010110100111001",
			2880 => "1111111010110100111001",
			2881 => "0001011100101100000100",
			2882 => "0000000010110100111001",
			2883 => "0000010110001100001100",
			2884 => "0011100001000000001000",
			2885 => "0010111010100100000100",
			2886 => "0000000010110100111001",
			2887 => "1111111010110100111001",
			2888 => "0000000010110100111001",
			2889 => "0000101001101000001000",
			2890 => "0001010011000100000100",
			2891 => "0000000010110100111001",
			2892 => "0000000010110100111001",
			2893 => "1111111010110100111001",
			2894 => "0001110011110101100100",
			2895 => "0000011101000000110100",
			2896 => "0010111010100100011100",
			2897 => "0000001110110000010100",
			2898 => "0010111011101100001100",
			2899 => "0011100110111000001000",
			2900 => "0000000100011000000100",
			2901 => "0000000010111000011101",
			2902 => "0000001010111000011101",
			2903 => "0000000010111000011101",
			2904 => "0010011001000100000100",
			2905 => "1111111010111000011101",
			2906 => "0000000010111000011101",
			2907 => "0000010111100100000100",
			2908 => "0000000010111000011101",
			2909 => "0000001010111000011101",
			2910 => "0010000000110000001100",
			2911 => "0001011100000000001000",
			2912 => "0001010011001000000100",
			2913 => "0000000010111000011101",
			2914 => "0000000010111000011101",
			2915 => "1111111010111000011101",
			2916 => "0001011100101100001000",
			2917 => "0000010011110000000100",
			2918 => "0000000010111000011101",
			2919 => "0000001010111000011101",
			2920 => "1111111010111000011101",
			2921 => "0001001001001000010000",
			2922 => "0011000111011100000100",
			2923 => "0000000010111000011101",
			2924 => "0001000011010000001000",
			2925 => "0001001010100100000100",
			2926 => "0000000010111000011101",
			2927 => "0000000010111000011101",
			2928 => "1111111010111000011101",
			2929 => "0011110000001100001000",
			2930 => "0010000000110000000100",
			2931 => "0000000010111000011101",
			2932 => "1111111010111000011101",
			2933 => "0000111101001000001000",
			2934 => "0010000011001000000100",
			2935 => "0000000010111000011101",
			2936 => "0000001010111000011101",
			2937 => "0000000110100100001000",
			2938 => "0010000011100100000100",
			2939 => "0000001010111000011101",
			2940 => "0000000010111000011101",
			2941 => "0000100100010100000100",
			2942 => "1111111010111000011101",
			2943 => "0000000010111000011101",
			2944 => "0011000011000000000100",
			2945 => "1111111010111000011101",
			2946 => "0000001010010000000100",
			2947 => "0000000010111000011101",
			2948 => "0000001111010000000100",
			2949 => "0000001010111000011101",
			2950 => "0000000010111000011101",
			2951 => "0000101111001101011000",
			2952 => "0011110101100101001000",
			2953 => "0001011100101100100100",
			2954 => "0010001111001000010100",
			2955 => "0010111011101100001000",
			2956 => "0010001111111100000100",
			2957 => "0000000010111100000001",
			2958 => "0000000010111100000001",
			2959 => "0000010011110000000100",
			2960 => "0000000010111100000001",
			2961 => "0011011010100100000100",
			2962 => "0000000010111100000001",
			2963 => "0000000010111100000001",
			2964 => "0001011000000000000100",
			2965 => "0000000010111100000001",
			2966 => "0011110010110000000100",
			2967 => "0000000010111100000001",
			2968 => "0010110101011100000100",
			2969 => "0000000010111100000001",
			2970 => "0000000010111100000001",
			2971 => "0010100000111100011000",
			2972 => "0001111001000000010000",
			2973 => "0001111111101000001000",
			2974 => "0011100100001100000100",
			2975 => "0000000010111100000001",
			2976 => "0000000010111100000001",
			2977 => "0001111000100000000100",
			2978 => "0000000010111100000001",
			2979 => "0000000010111100000001",
			2980 => "0011111011110100000100",
			2981 => "0000000010111100000001",
			2982 => "0000000010111100000001",
			2983 => "0000001100100100000100",
			2984 => "0000000010111100000001",
			2985 => "0000010111011100000100",
			2986 => "0000000010111100000001",
			2987 => "0000000010111100000001",
			2988 => "0011101110010000000100",
			2989 => "0000000010111100000001",
			2990 => "0001100100011000001000",
			2991 => "0001010011000100000100",
			2992 => "0000000010111100000001",
			2993 => "0000000010111100000001",
			2994 => "0000000010111100000001",
			2995 => "0001001101001000011000",
			2996 => "0010001010000100001100",
			2997 => "0010111010100100001000",
			2998 => "0000010111100100000100",
			2999 => "0000000010111100000001",
			3000 => "0000000010111100000001",
			3001 => "0000000010111100000001",
			3002 => "0010110011000000001000",
			3003 => "0001110011110100000100",
			3004 => "0000000010111100000001",
			3005 => "0000000010111100000001",
			3006 => "0000000010111100000001",
			3007 => "0000000010111100000001",
			3008 => "0010101101001000011100",
			3009 => "0000000100110100000100",
			3010 => "1111111010111111010101",
			3011 => "0001101110010000001000",
			3012 => "0011111100111000000100",
			3013 => "0000000010111111010101",
			3014 => "0000001010111111010101",
			3015 => "0001000111011100001100",
			3016 => "0001111001010000001000",
			3017 => "0001001011101100000100",
			3018 => "0000000010111111010101",
			3019 => "0000000010111111010101",
			3020 => "0000000010111111010101",
			3021 => "1111111010111111010101",
			3022 => "0000111100110000011100",
			3023 => "0000010011010000011000",
			3024 => "0000001010111000010100",
			3025 => "0001110001010000010000",
			3026 => "0000001100100100001000",
			3027 => "0001101111110000000100",
			3028 => "0000000010111111010101",
			3029 => "0000000010111111010101",
			3030 => "0001011100110000000100",
			3031 => "0000000010111111010101",
			3032 => "0000000010111111010101",
			3033 => "1111111010111111010101",
			3034 => "0000001010111111010101",
			3035 => "0000001010111111010101",
			3036 => "0001011011111000010100",
			3037 => "0010110101010100010000",
			3038 => "0011110101100100001000",
			3039 => "0011011110011000000100",
			3040 => "0000000010111111010101",
			3041 => "0000000010111111010101",
			3042 => "0001111100101100000100",
			3043 => "0000000010111111010101",
			3044 => "0000000010111111010101",
			3045 => "1111111010111111010101",
			3046 => "0001011100101100000100",
			3047 => "0000001010111111010101",
			3048 => "0000010110001100010000",
			3049 => "0010110011010000001000",
			3050 => "0010101011111000000100",
			3051 => "0000000010111111010101",
			3052 => "0000000010111111010101",
			3053 => "0010010110000000000100",
			3054 => "0000000010111111010101",
			3055 => "1111111010111111010101",
			3056 => "0000101001101000001000",
			3057 => "0001010011000100000100",
			3058 => "0000000010111111010101",
			3059 => "0000000010111111010101",
			3060 => "1111111010111111010101",
			3061 => "0001110011110101100000",
			3062 => "0011011100101000110000",
			3063 => "0010110101010100101000",
			3064 => "0001001100000000011100",
			3065 => "0001011001010000010000",
			3066 => "0000100101011000001000",
			3067 => "0010111010100100000100",
			3068 => "1111111011000010110001",
			3069 => "0000000011000010110001",
			3070 => "0011010110001100000100",
			3071 => "0000000011000010110001",
			3072 => "0000000011000010110001",
			3073 => "0000111000101000001000",
			3074 => "0011101111111000000100",
			3075 => "0000000011000010110001",
			3076 => "1111111011000010110001",
			3077 => "0000000011000010110001",
			3078 => "0011101001011100000100",
			3079 => "0000000011000010110001",
			3080 => "0000010111100100000100",
			3081 => "0000000011000010110001",
			3082 => "0000001011000010110001",
			3083 => "0000010110001100000100",
			3084 => "1111111011000010110001",
			3085 => "0000000011000010110001",
			3086 => "0010111001001000001100",
			3087 => "0001101110010000000100",
			3088 => "0000000011000010110001",
			3089 => "0011111011110100000100",
			3090 => "0000001011000010110001",
			3091 => "0000000011000010110001",
			3092 => "0000111100110000001100",
			3093 => "0000010011010000001000",
			3094 => "0011011001001000000100",
			3095 => "0000000011000010110001",
			3096 => "0000000011000010110001",
			3097 => "0000001011000010110001",
			3098 => "0011011010000100001100",
			3099 => "0001011011111000000100",
			3100 => "1111111011000010110001",
			3101 => "0001100010010000000100",
			3102 => "0000000011000010110001",
			3103 => "0000000011000010110001",
			3104 => "0000010101011100001000",
			3105 => "0001111001000000000100",
			3106 => "0000000011000010110001",
			3107 => "0000001011000010110001",
			3108 => "0000000011000010110001",
			3109 => "0011000011000000000100",
			3110 => "1111111011000010110001",
			3111 => "0000001010010000000100",
			3112 => "0000000011000010110001",
			3113 => "0000101001101000000100",
			3114 => "0000000011000010110001",
			3115 => "0000000011000010110001",
			3116 => "0000100100010101000100",
			3117 => "0000110100101100111000",
			3118 => "0010101001010100011100",
			3119 => "0010000011100100010100",
			3120 => "0010010101101100010000",
			3121 => "0010111010100100001000",
			3122 => "0011110000001100000100",
			3123 => "0000000011000110101101",
			3124 => "0000000011000110101101",
			3125 => "0001000101010100000100",
			3126 => "0000000011000110101101",
			3127 => "0000000011000110101101",
			3128 => "0000000011000110101101",
			3129 => "0010001000000000000100",
			3130 => "0000000011000110101101",
			3131 => "0000000011000110101101",
			3132 => "0010010011001000010000",
			3133 => "0011100110111000001100",
			3134 => "0001101111110000000100",
			3135 => "0000000011000110101101",
			3136 => "0000000110111100000100",
			3137 => "0000000011000110101101",
			3138 => "0000000011000110101101",
			3139 => "0000000011000110101101",
			3140 => "0011011010000100000100",
			3141 => "0000000011000110101101",
			3142 => "0001001100010000000100",
			3143 => "0000000011000110101101",
			3144 => "0000000011000110101101",
			3145 => "0000111110001100000100",
			3146 => "0000000011000110101101",
			3147 => "0001011111100000000100",
			3148 => "0000000011000110101101",
			3149 => "0000000011000110101101",
			3150 => "0001101000010100010100",
			3151 => "0001110100101100010000",
			3152 => "0011001010100100000100",
			3153 => "0000000011000110101101",
			3154 => "0001100101100000000100",
			3155 => "0000000011000110101101",
			3156 => "0001011001010100000100",
			3157 => "0000000011000110101101",
			3158 => "0000000011000110101101",
			3159 => "0000000011000110101101",
			3160 => "0000100111111000001000",
			3161 => "0011000101010100000100",
			3162 => "0000000011000110101101",
			3163 => "0000000011000110101101",
			3164 => "0010101101001000000100",
			3165 => "0000000011000110101101",
			3166 => "0000111001010000001100",
			3167 => "0011110100110100000100",
			3168 => "0000000011000110101101",
			3169 => "0000010111011100000100",
			3170 => "0000000011000110101101",
			3171 => "0000000011000110101101",
			3172 => "0010101001011000001000",
			3173 => "0011001001001000000100",
			3174 => "0000000011000110101101",
			3175 => "0000000011000110101101",
			3176 => "0001100010111100000100",
			3177 => "0000000011000110101101",
			3178 => "0000000011000110101101",
			3179 => "0000010111100100000100",
			3180 => "0000000011001001011001",
			3181 => "0000101111001100111100",
			3182 => "0010001000000000101100",
			3183 => "0010001111001000010000",
			3184 => "0000010011110000000100",
			3185 => "1111111011001001011001",
			3186 => "0011001010100100000100",
			3187 => "0000000011001001011001",
			3188 => "0000110011001000000100",
			3189 => "0000000011001001011001",
			3190 => "0000000011001001011001",
			3191 => "0011011001001000010000",
			3192 => "0000010110001100001000",
			3193 => "0001011100101100000100",
			3194 => "0000000011001001011001",
			3195 => "1111111011001001011001",
			3196 => "0010010011000000000100",
			3197 => "0000000011001001011001",
			3198 => "0000001011001001011001",
			3199 => "0000000100010100001000",
			3200 => "0011110100001000000100",
			3201 => "0000000011001001011001",
			3202 => "0000000011001001011001",
			3203 => "0000000011001001011001",
			3204 => "0010100000111100001000",
			3205 => "0001100101111100000100",
			3206 => "1111111011001001011001",
			3207 => "0000000011001001011001",
			3208 => "0000100110100100000100",
			3209 => "0000000011001001011001",
			3210 => "0000000011001001011001",
			3211 => "0011000101111000010100",
			3212 => "0011100101001100010000",
			3213 => "0010001010000100001000",
			3214 => "0010111010100100000100",
			3215 => "0000001011001001011001",
			3216 => "0000000011001001011001",
			3217 => "0000111111101000000100",
			3218 => "0000001011001001011001",
			3219 => "0000000011001001011001",
			3220 => "0000000011001001011001",
			3221 => "0000000011001001011001",
			3222 => "0010111101101001101000",
			3223 => "0000011101000001000000",
			3224 => "0010111010100100100100",
			3225 => "0001001100101000010100",
			3226 => "0011011110011000010000",
			3227 => "0011001011101100001000",
			3228 => "0000011000011000000100",
			3229 => "0000000011001101000101",
			3230 => "0000000011001101000101",
			3231 => "0000000100010100000100",
			3232 => "0000000011001101000101",
			3233 => "0000000011001101000101",
			3234 => "0000000011001101000101",
			3235 => "0000000100011000000100",
			3236 => "0000000011001101000101",
			3237 => "0010001111111100000100",
			3238 => "0000000011001101000101",
			3239 => "0011011011101100000100",
			3240 => "0000000011001101000101",
			3241 => "0000000011001101000101",
			3242 => "0011100001000000010100",
			3243 => "0011011100101000001100",
			3244 => "0001011100000000001000",
			3245 => "0010101000111000000100",
			3246 => "0000000011001101000101",
			3247 => "0000000011001101000101",
			3248 => "1111111011001101000101",
			3249 => "0010011111011000000100",
			3250 => "0000000011001101000101",
			3251 => "0000000011001101000101",
			3252 => "0011000101010100000100",
			3253 => "0000000011001101000101",
			3254 => "0000000011001101000101",
			3255 => "0011000101011100001100",
			3256 => "0010001001000100000100",
			3257 => "0000000011001101000101",
			3258 => "0001101110111100000100",
			3259 => "0000000011001101000101",
			3260 => "0000000011001101000101",
			3261 => "0010010101111000000100",
			3262 => "0000000011001101000101",
			3263 => "0000000110101000001100",
			3264 => "0000101100010100001000",
			3265 => "0001001101101000000100",
			3266 => "0000000011001101000101",
			3267 => "0000000011001101000101",
			3268 => "0000000011001101000101",
			3269 => "0001111010011100001000",
			3270 => "0001011000100000000100",
			3271 => "0000000011001101000101",
			3272 => "0000000011001101000101",
			3273 => "0000000011001101000101",
			3274 => "0001000110101100000100",
			3275 => "1111111011001101000101",
			3276 => "0000010111011100001000",
			3277 => "0011011010000100000100",
			3278 => "0000000011001101000101",
			3279 => "0000000011001101000101",
			3280 => "0000000011001101000101",
			3281 => "0011110010110000000100",
			3282 => "1111111011001110111001",
			3283 => "0010001111111100000100",
			3284 => "1111111011001110111001",
			3285 => "0001111100110000000100",
			3286 => "0000001011001110111001",
			3287 => "0000100100010100010100",
			3288 => "0010001000000000010000",
			3289 => "0000001100100100001000",
			3290 => "0011111100111000000100",
			3291 => "0000000011001110111001",
			3292 => "0000000011001110111001",
			3293 => "0011010111011100000100",
			3294 => "0000000011001110111001",
			3295 => "1111111011001110111001",
			3296 => "1111111011001110111001",
			3297 => "0010101111101000001100",
			3298 => "0011110101100100000100",
			3299 => "0000001011001110111001",
			3300 => "0011110100110100000100",
			3301 => "1111111011001110111001",
			3302 => "0000000011001110111001",
			3303 => "0001000011000000001000",
			3304 => "0010001010000100000100",
			3305 => "0000000011001110111001",
			3306 => "0000001011001110111001",
			3307 => "0010001100110000000100",
			3308 => "0000000011001110111001",
			3309 => "0000001011001110111001",
			3310 => "0000001000110001101100",
			3311 => "0000010110001101000000",
			3312 => "0010111011101100010000",
			3313 => "0001100100001000001100",
			3314 => "0000000100011000000100",
			3315 => "0000000011010010011101",
			3316 => "0011010110001100000100",
			3317 => "0000000011010010011101",
			3318 => "0000001011010010011101",
			3319 => "0000000011010010011101",
			3320 => "0011011100101000011000",
			3321 => "0011000101010100001100",
			3322 => "0010001010000100001000",
			3323 => "0000011101000000000100",
			3324 => "0000000011010010011101",
			3325 => "0000000011010010011101",
			3326 => "0000000011010010011101",
			3327 => "0010110011010000000100",
			3328 => "0000000011010010011101",
			3329 => "0001001010000100000100",
			3330 => "0000000011010010011101",
			3331 => "1111111011010010011101",
			3332 => "0001011100101100001100",
			3333 => "0010001111011000000100",
			3334 => "0000000011010010011101",
			3335 => "0001101100010000000100",
			3336 => "0000000011010010011101",
			3337 => "0000001011010010011101",
			3338 => "0010000000110000000100",
			3339 => "1111111011010010011101",
			3340 => "0000011101000000000100",
			3341 => "0000000011010010011101",
			3342 => "0000000011010010011101",
			3343 => "0001001001001000001100",
			3344 => "0001000011010000001000",
			3345 => "0010001111011000000100",
			3346 => "0000000011010010011101",
			3347 => "0000000011010010011101",
			3348 => "1111111011010010011101",
			3349 => "0010111001001000001100",
			3350 => "0010010011000000000100",
			3351 => "0000000011010010011101",
			3352 => "0010011111011000000100",
			3353 => "0000001011010010011101",
			3354 => "0000000011010010011101",
			3355 => "0011111001111000000100",
			3356 => "1111111011010010011101",
			3357 => "0000111001010000001000",
			3358 => "0001001111011000000100",
			3359 => "0000001011010010011101",
			3360 => "0000000011010010011101",
			3361 => "0010101001011000000100",
			3362 => "1111111011010010011101",
			3363 => "0000000011010010011101",
			3364 => "0001100000100100000100",
			3365 => "0000001011010010011101",
			3366 => "0000000011010010011101",
			3367 => "0000001000110001011100",
			3368 => "0011110101100101000000",
			3369 => "0000001110110000110000",
			3370 => "0001011100101100100000",
			3371 => "0000100101011000010000",
			3372 => "0010101001010100001000",
			3373 => "0011010011010000000100",
			3374 => "1111111011010101100001",
			3375 => "0000000011010101100001",
			3376 => "0001111100110000000100",
			3377 => "0000001011010101100001",
			3378 => "0000000011010101100001",
			3379 => "0010101000101000001000",
			3380 => "0000011001100000000100",
			3381 => "0000000011010101100001",
			3382 => "0000001011010101100001",
			3383 => "0010101111101000000100",
			3384 => "1111111011010101100001",
			3385 => "0000000011010101100001",
			3386 => "0000010110001100000100",
			3387 => "1111111011010101100001",
			3388 => "0011000101101100000100",
			3389 => "0000000011010101100001",
			3390 => "0001111001000000000100",
			3391 => "1111111011010101100001",
			3392 => "0000000011010101100001",
			3393 => "0000010011010000001100",
			3394 => "0001001000000100001000",
			3395 => "0000011001100000000100",
			3396 => "0000000011010101100001",
			3397 => "0000000011010101100001",
			3398 => "0000000011010101100001",
			3399 => "0000001011010101100001",
			3400 => "0011110000101100000100",
			3401 => "1111111011010101100001",
			3402 => "0011100101100000010100",
			3403 => "0011000101111000010000",
			3404 => "0001011011111000001000",
			3405 => "0000001010111000000100",
			3406 => "1111111011010101100001",
			3407 => "0000000011010101100001",
			3408 => "0001010011000100000100",
			3409 => "0000000011010101100001",
			3410 => "0000000011010101100001",
			3411 => "1111111011010101100001",
			3412 => "1111111011010101100001",
			3413 => "0001100000100100000100",
			3414 => "0000001011010101100001",
			3415 => "0000000011010101100001",
			3416 => "0000101010010001001100",
			3417 => "0000110000111001000100",
			3418 => "0001010001001000111100",
			3419 => "0010001010000100100000",
			3420 => "0010111011101100010000",
			3421 => "0010010101011100001000",
			3422 => "0001001010000100000100",
			3423 => "0000000011010111111111",
			3424 => "0000000011010111111111",
			3425 => "0001001100101000000100",
			3426 => "0000000011010111111111",
			3427 => "0000000011010111111111",
			3428 => "0001101010110000001000",
			3429 => "0001001100000000000100",
			3430 => "0000000011010111111111",
			3431 => "0000000011010111111111",
			3432 => "0001100111010000000100",
			3433 => "0000000011010111111111",
			3434 => "0000000011010111111111",
			3435 => "0010110101010100001100",
			3436 => "0000001101001100000100",
			3437 => "0000000011010111111111",
			3438 => "0000001000010000000100",
			3439 => "0000000011010111111111",
			3440 => "0000000011010111111111",
			3441 => "0010011000000100001000",
			3442 => "0001110110011100000100",
			3443 => "0000000011010111111111",
			3444 => "0000000011010111111111",
			3445 => "0010110101101100000100",
			3446 => "0000000011010111111111",
			3447 => "0000000011010111111111",
			3448 => "0001001000000000000100",
			3449 => "0000000011010111111111",
			3450 => "1111111011010111111111",
			3451 => "0011111000101100000100",
			3452 => "0000000011010111111111",
			3453 => "0000000011010111111111",
			3454 => "0000000011010111111111",
			3455 => "0010100000111100100100",
			3456 => "0010100011000100100000",
			3457 => "0000111100101100011100",
			3458 => "0010101001011000010100",
			3459 => "0000011100101000001100",
			3460 => "0000010101011100001000",
			3461 => "0000100101010000000100",
			3462 => "0000000011011001101001",
			3463 => "0000000011011001101001",
			3464 => "1111111011011001101001",
			3465 => "0000011001000100000100",
			3466 => "0000001011011001101001",
			3467 => "1111111011011001101001",
			3468 => "0000010110001100000100",
			3469 => "0000000011011001101001",
			3470 => "0000001011011001101001",
			3471 => "1111111011011001101001",
			3472 => "1111111011011001101001",
			3473 => "0000001100100100000100",
			3474 => "1111111011011001101001",
			3475 => "0001101110000100001100",
			3476 => "0000000101101000001000",
			3477 => "0001101010101100000100",
			3478 => "0000001011011001101001",
			3479 => "1111111011011001101001",
			3480 => "0000001011011001101001",
			3481 => "1111111011011001101001",
			3482 => "0000101110000100000100",
			3483 => "1111111011011011010101",
			3484 => "0001111100110000010000",
			3485 => "0011011011101100001000",
			3486 => "0001110011001000000100",
			3487 => "0000000011011011010101",
			3488 => "0000000011011011010101",
			3489 => "0001101110111100000100",
			3490 => "0000000011011011010101",
			3491 => "0000001011011011010101",
			3492 => "0011111010101100000100",
			3493 => "1111111011011011010101",
			3494 => "0011111110101100001000",
			3495 => "0010111100101000000100",
			3496 => "0000001011011011010101",
			3497 => "0000000011011011010101",
			3498 => "0000001101011100001000",
			3499 => "0001110001010000000100",
			3500 => "0000000011011011010101",
			3501 => "1111111011011011010101",
			3502 => "0010001010000100001000",
			3503 => "0010111010100100000100",
			3504 => "0000000011011011010101",
			3505 => "1111111011011011010101",
			3506 => "0010110101010100000100",
			3507 => "0000001011011011010101",
			3508 => "0000000011011011010101",
			3509 => "0000011101000000101100",
			3510 => "0010111010100100011100",
			3511 => "0000100111111000010100",
			3512 => "0001001111011000001100",
			3513 => "0010101000000000001000",
			3514 => "0000011001100000000100",
			3515 => "0000000011011110101001",
			3516 => "0000000011011110101001",
			3517 => "0000000011011110101001",
			3518 => "0010101111101000000100",
			3519 => "0000000011011110101001",
			3520 => "0000000011011110101001",
			3521 => "0000010111100100000100",
			3522 => "0000000011011110101001",
			3523 => "0000000011011110101001",
			3524 => "0011000011010000001000",
			3525 => "0000111000101000000100",
			3526 => "0000000011011110101001",
			3527 => "0000000011011110101001",
			3528 => "0010000011001000000100",
			3529 => "0000000011011110101001",
			3530 => "0000000011011110101001",
			3531 => "0001111001011000011000",
			3532 => "0010111001001000001100",
			3533 => "0011111100111000001000",
			3534 => "0001001001000100000100",
			3535 => "0000000011011110101001",
			3536 => "0000000011011110101001",
			3537 => "0000000011011110101001",
			3538 => "0010011000000100000100",
			3539 => "0000000011011110101001",
			3540 => "0001011011000000000100",
			3541 => "0000000011011110101001",
			3542 => "0000000011011110101001",
			3543 => "0000010011010000001100",
			3544 => "0010101100001100001000",
			3545 => "0001101110000100000100",
			3546 => "0000000011011110101001",
			3547 => "0000000011011110101001",
			3548 => "0000000011011110101001",
			3549 => "0000111001010000001100",
			3550 => "0011010011000000001000",
			3551 => "0000001111001100000100",
			3552 => "0000000011011110101001",
			3553 => "0000000011011110101001",
			3554 => "0000000011011110101001",
			3555 => "0001001100010000000100",
			3556 => "0000000011011110101001",
			3557 => "0001010001001000000100",
			3558 => "0000000011011110101001",
			3559 => "0000110000111000000100",
			3560 => "0000000011011110101001",
			3561 => "0000000011011110101001",
			3562 => "0011110100010000001100",
			3563 => "0011000011010000001000",
			3564 => "0010001111001000000100",
			3565 => "1111111011100000010101",
			3566 => "0000001011100000010101",
			3567 => "1111111011100000010101",
			3568 => "0000010111100100000100",
			3569 => "1111111011100000010101",
			3570 => "0011010011000000100100",
			3571 => "0010101100001100011100",
			3572 => "0010110011010000010000",
			3573 => "0001010011001000001000",
			3574 => "0011001110011000000100",
			3575 => "1111111011100000010101",
			3576 => "0000000011100000010101",
			3577 => "0010001111111100000100",
			3578 => "1111111011100000010101",
			3579 => "0000001011100000010101",
			3580 => "0000010011110000000100",
			3581 => "1111111011100000010101",
			3582 => "0000111001010000000100",
			3583 => "0000001011100000010101",
			3584 => "0000000011100000010101",
			3585 => "0000001010101000000100",
			3586 => "1111111011100000010101",
			3587 => "0000001011100000010101",
			3588 => "1111111011100000010101",
			3589 => "0000011101000000101100",
			3590 => "0010111010100100011100",
			3591 => "0000100111111000010100",
			3592 => "0001001111011000001100",
			3593 => "0010101000000000001000",
			3594 => "0000000010101100000100",
			3595 => "0000000011100011101001",
			3596 => "0000000011100011101001",
			3597 => "0000000011100011101001",
			3598 => "0010101111101000000100",
			3599 => "0000000011100011101001",
			3600 => "0000000011100011101001",
			3601 => "0000010111100100000100",
			3602 => "0000000011100011101001",
			3603 => "0000000011100011101001",
			3604 => "0011000011010000001000",
			3605 => "0000111000101000000100",
			3606 => "0000000011100011101001",
			3607 => "0000000011100011101001",
			3608 => "0010000011001000000100",
			3609 => "0000000011100011101001",
			3610 => "0000000011100011101001",
			3611 => "0001111001011000010100",
			3612 => "0011111100111000001100",
			3613 => "0000110011000000001000",
			3614 => "0001111100000000000100",
			3615 => "0000000011100011101001",
			3616 => "0000000011100011101001",
			3617 => "0000000011100011101001",
			3618 => "0000010110001100000100",
			3619 => "0000000011100011101001",
			3620 => "0000000011100011101001",
			3621 => "0001000011000000001000",
			3622 => "0011011101101000000100",
			3623 => "0000000011100011101001",
			3624 => "0000000011100011101001",
			3625 => "0001001100010000001100",
			3626 => "0010001001010100001000",
			3627 => "0000111100110000000100",
			3628 => "0000000011100011101001",
			3629 => "0000000011100011101001",
			3630 => "0000000011100011101001",
			3631 => "0011011010000100001100",
			3632 => "0000110000111100001000",
			3633 => "0000010101010100000100",
			3634 => "0000000011100011101001",
			3635 => "0000000011100011101001",
			3636 => "0000000011100011101001",
			3637 => "0000010111011100001000",
			3638 => "0000011110011000000100",
			3639 => "0000000011100011101001",
			3640 => "0000000011100011101001",
			3641 => "0000000011100011101001",
			3642 => "0000011001100000100000",
			3643 => "0011110011101100001000",
			3644 => "0001100001001100000100",
			3645 => "0000000011100110101101",
			3646 => "0000000011100110101101",
			3647 => "0011101100000100010100",
			3648 => "0000111111011000001100",
			3649 => "0001111101001000001000",
			3650 => "0000111101101000000100",
			3651 => "0000000011100110101101",
			3652 => "0000000011100110101101",
			3653 => "0000000011100110101101",
			3654 => "0001111001011000000100",
			3655 => "0000000011100110101101",
			3656 => "0000000011100110101101",
			3657 => "0000000011100110101101",
			3658 => "0001111100011100110000",
			3659 => "0010100000111100011100",
			3660 => "0001011000100000010100",
			3661 => "0011010011000000010000",
			3662 => "0000101111001100001000",
			3663 => "0011110000100100000100",
			3664 => "0000000011100110101101",
			3665 => "0000000011100110101101",
			3666 => "0001101011011100000100",
			3667 => "0000000011100110101101",
			3668 => "0000000011100110101101",
			3669 => "0000000011100110101101",
			3670 => "0001110001010000000100",
			3671 => "0000000011100110101101",
			3672 => "0000000011100110101101",
			3673 => "0010011100000000001000",
			3674 => "0000010110001100000100",
			3675 => "0000000011100110101101",
			3676 => "0000000011100110101101",
			3677 => "0011000101111000001000",
			3678 => "0001011010110100000100",
			3679 => "0000000011100110101101",
			3680 => "0000000011100110101101",
			3681 => "0000000011100110101101",
			3682 => "0011000011000000001000",
			3683 => "0011110100111100000100",
			3684 => "0000000011100110101101",
			3685 => "0000000011100110101101",
			3686 => "0000001010010000000100",
			3687 => "0000000011100110101101",
			3688 => "0000101001101000000100",
			3689 => "0000000011100110101101",
			3690 => "0000000011100110101101",
			3691 => "0011110000001100010100",
			3692 => "0011110010110000000100",
			3693 => "1111111011101001010001",
			3694 => "0011100000010100000100",
			3695 => "0000001011101001010001",
			3696 => "0001100011011000001000",
			3697 => "0011001100101000000100",
			3698 => "0000001011101001010001",
			3699 => "1111111011101001010001",
			3700 => "1111111011101001010001",
			3701 => "0011011101101000110100",
			3702 => "0000011001100000010000",
			3703 => "0010000101101100000100",
			3704 => "1111111011101001010001",
			3705 => "0010111010100100001000",
			3706 => "0011111101001100000100",
			3707 => "1111111011101001010001",
			3708 => "0000010011101001010001",
			3709 => "1111111011101001010001",
			3710 => "0000001010111000011000",
			3711 => "0010000011100100010000",
			3712 => "0010001111001000001000",
			3713 => "0011001010100100000100",
			3714 => "0000010011101001010001",
			3715 => "1111111011101001010001",
			3716 => "0011110111000000000100",
			3717 => "0000011011101001010001",
			3718 => "0000001011101001010001",
			3719 => "0001010110011100000100",
			3720 => "0000000011101001010001",
			3721 => "1111111011101001010001",
			3722 => "0001011000100000001000",
			3723 => "0010001010000100000100",
			3724 => "0000010011101001010001",
			3725 => "0000010011101001010001",
			3726 => "0000001011101001010001",
			3727 => "0000010111011100001000",
			3728 => "0011011010000100000100",
			3729 => "1111111011101001010001",
			3730 => "0000001011101001010001",
			3731 => "1111111011101001010001",
			3732 => "0010001010000100110100",
			3733 => "0010111011101100001100",
			3734 => "0001010011001000000100",
			3735 => "1111111011101100101101",
			3736 => "0010001111111100000100",
			3737 => "0000000011101100101101",
			3738 => "0000001011101100101101",
			3739 => "0001011001010000011000",
			3740 => "0000011101000000010000",
			3741 => "0011111000100100001100",
			3742 => "0001001010000100000100",
			3743 => "1111111011101100101101",
			3744 => "0001111001010100000100",
			3745 => "1111111011101100101101",
			3746 => "0000000011101100101101",
			3747 => "0000000011101100101101",
			3748 => "0011000101011100000100",
			3749 => "0000001011101100101101",
			3750 => "0000000011101100101101",
			3751 => "0001010011000100001000",
			3752 => "0010011001001000000100",
			3753 => "0000000011101100101101",
			3754 => "1111111011101100101101",
			3755 => "0001010001001000000100",
			3756 => "0000000011101100101101",
			3757 => "1111111011101100101101",
			3758 => "0010110101011100010000",
			3759 => "0001011011000000001100",
			3760 => "0001000101111000001000",
			3761 => "0001011100110000000100",
			3762 => "0000001011101100101101",
			3763 => "0000000011101100101101",
			3764 => "0000001011101100101101",
			3765 => "0000000011101100101101",
			3766 => "0000010110001100010000",
			3767 => "0010101011111000001000",
			3768 => "0001111100101100000100",
			3769 => "1111111011101100101101",
			3770 => "0000000011101100101101",
			3771 => "0010000011100100000100",
			3772 => "1111111011101100101101",
			3773 => "0000000011101100101101",
			3774 => "0001001001000100001100",
			3775 => "0000011110011000001000",
			3776 => "0001001010100100000100",
			3777 => "0000000011101100101101",
			3778 => "0000000011101100101101",
			3779 => "1111111011101100101101",
			3780 => "0011011001001000000100",
			3781 => "0000001011101100101101",
			3782 => "0000111100010000000100",
			3783 => "0000001011101100101101",
			3784 => "0001011011111000000100",
			3785 => "1111111011101100101101",
			3786 => "0000000011101100101101",
			3787 => "0011110100010000001100",
			3788 => "0011000011010000001000",
			3789 => "0011011010100100000100",
			3790 => "1111111011101110100001",
			3791 => "0000010011101110100001",
			3792 => "1111111011101110100001",
			3793 => "0000010111100100000100",
			3794 => "1111111011101110100001",
			3795 => "0011010101111000101000",
			3796 => "0000001010111000011000",
			3797 => "0010001111001000001000",
			3798 => "0010111011101100000100",
			3799 => "0000001011101110100001",
			3800 => "1111111011101110100001",
			3801 => "0010110101011100001000",
			3802 => "0010011001000100000100",
			3803 => "0000000011101110100001",
			3804 => "0000001011101110100001",
			3805 => "0000010110001100000100",
			3806 => "1111111011101110100001",
			3807 => "0000000011101110100001",
			3808 => "0011100101001100001100",
			3809 => "0010001010000100000100",
			3810 => "0000000011101110100001",
			3811 => "0001011100101100000100",
			3812 => "0000001011101110100001",
			3813 => "0000001011101110100001",
			3814 => "0000000011101110100001",
			3815 => "1111111011101110100001",
			3816 => "0011110100010000001100",
			3817 => "0010111011101100001000",
			3818 => "0000001010001000000100",
			3819 => "1111111011110000001101",
			3820 => "0000010011110000001101",
			3821 => "1111111011110000001101",
			3822 => "0000010111100100000100",
			3823 => "1111111011110000001101",
			3824 => "0001111100110000000100",
			3825 => "0000001011110000001101",
			3826 => "0001111110001100100000",
			3827 => "0000011101000000010000",
			3828 => "0010111010100100001000",
			3829 => "0001011000000000000100",
			3830 => "0000000011110000001101",
			3831 => "0000001011110000001101",
			3832 => "0000010011110000000100",
			3833 => "1111111011110000001101",
			3834 => "0000000011110000001101",
			3835 => "0011000101011100001000",
			3836 => "0001001010000100000100",
			3837 => "0000000011110000001101",
			3838 => "0000001011110000001101",
			3839 => "0000000110101000000100",
			3840 => "1111111011110000001101",
			3841 => "0000000011110000001101",
			3842 => "1111111011110000001101",
			3843 => "0010100000111101001000",
			3844 => "0000001010111000110000",
			3845 => "0011110000100100100000",
			3846 => "0010100011000100011100",
			3847 => "0001001100000000010000",
			3848 => "0001000011000000001000",
			3849 => "0000100100010100000100",
			3850 => "0000000011110010111001",
			3851 => "0000000011110010111001",
			3852 => "0011111110000100000100",
			3853 => "0000000011110010111001",
			3854 => "0000000011110010111001",
			3855 => "0010000011100100001000",
			3856 => "0000111100101100000100",
			3857 => "0000001011110010111001",
			3858 => "0000000011110010111001",
			3859 => "0000000011110010111001",
			3860 => "0000000011110010111001",
			3861 => "0010101001011000001100",
			3862 => "0001000110000000001000",
			3863 => "0010101111101000000100",
			3864 => "0000000011110010111001",
			3865 => "0000000011110010111001",
			3866 => "0000000011110010111001",
			3867 => "0000000011110010111001",
			3868 => "0011011101101000010000",
			3869 => "0010001010000100001100",
			3870 => "0010111010100100001000",
			3871 => "0011011011101100000100",
			3872 => "0000000011110010111001",
			3873 => "0000000011110010111001",
			3874 => "0000000011110010111001",
			3875 => "0000000011110010111001",
			3876 => "0001001000000000000100",
			3877 => "0000000011110010111001",
			3878 => "0000000011110010111001",
			3879 => "0001101110000100001100",
			3880 => "0000000110111100000100",
			3881 => "0000000011110010111001",
			3882 => "0000010111011100000100",
			3883 => "0000001011110010111001",
			3884 => "0000000011110010111001",
			3885 => "0000000011110010111001",
			3886 => "0010100000111100111100",
			3887 => "0001010001001000111000",
			3888 => "0010000011100100100100",
			3889 => "0001001100000000010100",
			3890 => "0001000011001000010000",
			3891 => "0000000111111000001000",
			3892 => "0011110010000100000100",
			3893 => "0000000011110101011101",
			3894 => "1111111011110101011101",
			3895 => "0010000000110000000100",
			3896 => "0000000011110101011101",
			3897 => "0000000011110101011101",
			3898 => "1111111011110101011101",
			3899 => "0000111111101000001100",
			3900 => "0000100010100100001000",
			3901 => "0000011001100000000100",
			3902 => "0000000011110101011101",
			3903 => "0000000011110101011101",
			3904 => "0000001011110101011101",
			3905 => "0000000011110101011101",
			3906 => "0000101111001100001100",
			3907 => "0001111011111000000100",
			3908 => "0000000011110101011101",
			3909 => "0001100101111100000100",
			3910 => "1111111011110101011101",
			3911 => "0000000011110101011101",
			3912 => "0000111001010000000100",
			3913 => "0000000011110101011101",
			3914 => "0000000011110101011101",
			3915 => "1111111011110101011101",
			3916 => "0001011100011100001000",
			3917 => "0011101101100100000100",
			3918 => "0000000011110101011101",
			3919 => "0000001011110101011101",
			3920 => "0010101100001100000100",
			3921 => "0000000011110101011101",
			3922 => "0010111101101000001000",
			3923 => "0010001010000100000100",
			3924 => "0000000011110101011101",
			3925 => "0000000011110101011101",
			3926 => "0000000011110101011101",
			3927 => "0010001000000001010100",
			3928 => "0010001111001000100000",
			3929 => "0000101011001100010100",
			3930 => "0011110011101100001000",
			3931 => "0001101110111100000100",
			3932 => "0000000011111000110001",
			3933 => "0000000011111000110001",
			3934 => "0010101100010000001000",
			3935 => "0010101000000100000100",
			3936 => "0000000011111000110001",
			3937 => "0000000011111000110001",
			3938 => "0000000011111000110001",
			3939 => "0011101110010000001000",
			3940 => "0000010111100100000100",
			3941 => "0000000011111000110001",
			3942 => "0000000011111000110001",
			3943 => "0000000011111000110001",
			3944 => "0011000101010100001100",
			3945 => "0001011000000100000100",
			3946 => "0000000011111000110001",
			3947 => "0011110010110000000100",
			3948 => "0000000011111000110001",
			3949 => "0000000011111000110001",
			3950 => "0010001111011000011000",
			3951 => "0001001100000000010000",
			3952 => "0011011001001000001000",
			3953 => "0001100111101000000100",
			3954 => "0000000011111000110001",
			3955 => "0000000011111000110001",
			3956 => "0011011001000100000100",
			3957 => "0000000011111000110001",
			3958 => "0000000011111000110001",
			3959 => "0000000110010100000100",
			3960 => "0000000011111000110001",
			3961 => "0000000011111000110001",
			3962 => "0011111101010000000100",
			3963 => "0000000011111000110001",
			3964 => "0011001101101000001000",
			3965 => "0000011110011000000100",
			3966 => "0000000011111000110001",
			3967 => "0000000011111000110001",
			3968 => "0000000011111000110001",
			3969 => "0001000011000000001000",
			3970 => "0010001100110000000100",
			3971 => "0000000011111000110001",
			3972 => "0000000011111000110001",
			3973 => "0010001001010100001000",
			3974 => "0000111010100000000100",
			3975 => "0000000011111000110001",
			3976 => "0000000011111000110001",
			3977 => "0011101010001000000100",
			3978 => "0000000011111000110001",
			3979 => "0000000011111000110001",
			3980 => "0011110100010000001100",
			3981 => "0011000011010000001000",
			3982 => "0000011101000000000100",
			3983 => "1111111011111010111101",
			3984 => "0000001011111010111101",
			3985 => "1111111011111010111101",
			3986 => "0000010111100100000100",
			3987 => "1111111011111010111101",
			3988 => "0011000101010100011000",
			3989 => "0001010011001000001000",
			3990 => "0000110011001000000100",
			3991 => "0000000011111010111101",
			3992 => "1111111011111010111101",
			3993 => "0010011101101000001100",
			3994 => "0001110110101100000100",
			3995 => "0000001011111010111101",
			3996 => "0010110011010000000100",
			3997 => "0000000011111010111101",
			3998 => "1111111011111010111101",
			3999 => "0000001011111010111101",
			4000 => "0000010110001100001100",
			4001 => "0011011100101000001000",
			4002 => "0010110101010100000100",
			4003 => "0000000011111010111101",
			4004 => "1111111011111010111101",
			4005 => "0000001011111010111101",
			4006 => "0000111000000000000100",
			4007 => "1111111011111010111101",
			4008 => "0000111001010000001000",
			4009 => "0000100000101000000100",
			4010 => "0000000011111010111101",
			4011 => "0000001011111010111101",
			4012 => "0010111001001000000100",
			4013 => "0000001011111010111101",
			4014 => "0000000011111010111101",
			4015 => "0011110010110000000100",
			4016 => "1111111011111101000001",
			4017 => "0010000101101100001100",
			4018 => "0010101000000000001000",
			4019 => "0010011100101000000100",
			4020 => "1111111011111101000001",
			4021 => "0000001011111101000001",
			4022 => "1111111011111101000001",
			4023 => "0011000111011100010100",
			4024 => "0001010011001000000100",
			4025 => "0000000011111101000001",
			4026 => "0001110001010000001000",
			4027 => "0011000011010000000100",
			4028 => "0000001011111101000001",
			4029 => "0000001011111101000001",
			4030 => "0000000000101000000100",
			4031 => "1111111011111101000001",
			4032 => "0000001011111101000001",
			4033 => "0001000110000000001000",
			4034 => "0011111000001000000100",
			4035 => "1111111011111101000001",
			4036 => "0000000011111101000001",
			4037 => "0010001111001000001000",
			4038 => "0010011010000100000100",
			4039 => "1111111011111101000001",
			4040 => "0000000011111101000001",
			4041 => "0011000101011100001000",
			4042 => "0001001111011000000100",
			4043 => "0000000011111101000001",
			4044 => "0000001011111101000001",
			4045 => "0010010011000000000100",
			4046 => "1111111011111101000001",
			4047 => "0000000011111101000001",
			4048 => "0001101010001000010100",
			4049 => "0000011000011000010000",
			4050 => "0010111010100100001100",
			4051 => "0001001111011000000100",
			4052 => "0000000011111111101101",
			4053 => "0000010001110000000100",
			4054 => "0000000011111111101101",
			4055 => "0000000011111111101101",
			4056 => "0000000011111111101101",
			4057 => "1111111011111111101101",
			4058 => "0011111110101100001100",
			4059 => "0010111100101000001000",
			4060 => "0000001011001000000100",
			4061 => "0000000011111111101101",
			4062 => "0000000011111111101101",
			4063 => "0000000011111111101101",
			4064 => "0000001101011100001100",
			4065 => "0001001100101000001000",
			4066 => "0001111111101000000100",
			4067 => "0000000011111111101101",
			4068 => "0000000011111111101101",
			4069 => "1111111011111111101101",
			4070 => "0001110011110100100000",
			4071 => "0001101110001000010000",
			4072 => "0001001100000000001000",
			4073 => "0000101101110000000100",
			4074 => "1111111011111111101101",
			4075 => "0000000011111111101101",
			4076 => "0000000110100100000100",
			4077 => "0000000011111111101101",
			4078 => "0000000011111111101101",
			4079 => "0001101010101100001000",
			4080 => "0011101110100000000100",
			4081 => "0000000011111111101101",
			4082 => "0000001011111111101101",
			4083 => "0010111100101000000100",
			4084 => "0000000011111111101101",
			4085 => "0000000011111111101101",
			4086 => "0011000011000000000100",
			4087 => "0000000011111111101101",
			4088 => "0011010011000000000100",
			4089 => "0000000011111111101101",
			4090 => "0000000011111111101101",
			4091 => "0000001110110001000100",
			4092 => "0010001111001000010100",
			4093 => "0010111011101100010000",
			4094 => "0011001011101100000100",
			4095 => "0000000100000010101001",
			4096 => "0010110110001100000100",
			4097 => "0000000100000010101001",
			4098 => "0000010001110000000100",
			4099 => "0000000100000010101001",
			4100 => "0000000100000010101001",
			4101 => "0000000100000010101001",
			4102 => "0011000101101100011000",
			4103 => "0010111001001000010100",
			4104 => "0000000100110100001000",
			4105 => "0000110011000000000100",
			4106 => "0000000100000010101001",
			4107 => "0000000100000010101001",
			4108 => "0001011001011000001000",
			4109 => "0001011101001000000100",
			4110 => "0000000100000010101001",
			4111 => "0000000100000010101001",
			4112 => "0000000100000010101001",
			4113 => "0000000100000010101001",
			4114 => "0000000100010100001000",
			4115 => "0011110101111100000100",
			4116 => "0000000100000010101001",
			4117 => "0000000100000010101001",
			4118 => "0000111001000000001100",
			4119 => "0010001000000000000100",
			4120 => "0000000100000010101001",
			4121 => "0001101010101100000100",
			4122 => "0000000100000010101001",
			4123 => "0000000100000010101001",
			4124 => "0000000100000010101001",
			4125 => "0010010110101100011000",
			4126 => "0000010111100100000100",
			4127 => "0000000100000010101001",
			4128 => "0011100101001100010000",
			4129 => "0010001010000100001000",
			4130 => "0010111010100100000100",
			4131 => "0000000100000010101001",
			4132 => "0000000100000010101001",
			4133 => "0000010101011100000100",
			4134 => "0000000100000010101001",
			4135 => "0000000100000010101001",
			4136 => "0000000100000010101001",
			4137 => "0000000100000010101001",
			4138 => "0000100100010101010000",
			4139 => "0011000101101100111100",
			4140 => "0001101010001000011100",
			4141 => "0000011000011000010000",
			4142 => "0010111010100100001100",
			4143 => "0000110011001000000100",
			4144 => "0000000100000110110101",
			4145 => "0000001000100100000100",
			4146 => "0000000100000110110101",
			4147 => "0000000100000110110101",
			4148 => "0000000100000110110101",
			4149 => "0000110011000000001000",
			4150 => "0000111001000100000100",
			4151 => "0000000100000110110101",
			4152 => "0000000100000110110101",
			4153 => "0000000100000110110101",
			4154 => "0001100001100000001100",
			4155 => "0011111110101100001000",
			4156 => "0000010111100100000100",
			4157 => "0000000100000110110101",
			4158 => "0000000100000110110101",
			4159 => "0000000100000110110101",
			4160 => "0000000100010100001000",
			4161 => "0001001100101000000100",
			4162 => "0000000100000110110101",
			4163 => "0000000100000110110101",
			4164 => "0001100111101000000100",
			4165 => "0000000100000110110101",
			4166 => "0011111011000100000100",
			4167 => "0000000100000110110101",
			4168 => "0000000100000110110101",
			4169 => "0000011100101000001100",
			4170 => "0010100111010100000100",
			4171 => "0000000100000110110101",
			4172 => "0001010000110100000100",
			4173 => "0000000100000110110101",
			4174 => "0000000100000110110101",
			4175 => "0011100110111000000100",
			4176 => "0000000100000110110101",
			4177 => "0000000100000110110101",
			4178 => "0001100100100000010100",
			4179 => "0001101110001000001000",
			4180 => "0000001110110000000100",
			4181 => "0000000100000110110101",
			4182 => "0000000100000110110101",
			4183 => "0011111011010100001000",
			4184 => "0000010011110000000100",
			4185 => "0000000100000110110101",
			4186 => "0000000100000110110101",
			4187 => "0000000100000110110101",
			4188 => "0000001101011000010000",
			4189 => "0011010101101100001000",
			4190 => "0000111000101000000100",
			4191 => "0000000100000110110101",
			4192 => "0000000100000110110101",
			4193 => "0001010011000100000100",
			4194 => "0000000100000110110101",
			4195 => "0000000100000110110101",
			4196 => "0000010101010100001100",
			4197 => "0000101110101000001000",
			4198 => "0010000000110000000100",
			4199 => "0000000100000110110101",
			4200 => "0000000100000110110101",
			4201 => "0000000100000110110101",
			4202 => "0000011100101000000100",
			4203 => "0000000100000110110101",
			4204 => "0000000100000110110101",
			4205 => "0000001101111000111100",
			4206 => "0000011011101100110000",
			4207 => "0001001100000000100100",
			4208 => "0001111111101000010100",
			4209 => "0000100101011000001100",
			4210 => "0011110011101100001000",
			4211 => "0000010110110100000100",
			4212 => "0000000100001001111001",
			4213 => "0000000100001001111001",
			4214 => "0000000100001001111001",
			4215 => "0000011001100000000100",
			4216 => "0000000100001001111001",
			4217 => "0000000100001001111001",
			4218 => "0001110110011100001100",
			4219 => "0000001010000000001000",
			4220 => "0001100001100000000100",
			4221 => "0000000100001001111001",
			4222 => "0000000100001001111001",
			4223 => "0000000100001001111001",
			4224 => "0000000100001001111001",
			4225 => "0000000010100100001000",
			4226 => "0010101000101000000100",
			4227 => "0000000100001001111001",
			4228 => "0000000100001001111001",
			4229 => "0000000100001001111001",
			4230 => "0000101100010100001000",
			4231 => "0010110101101100000100",
			4232 => "0000000100001001111001",
			4233 => "0000000100001001111001",
			4234 => "0000000100001001111001",
			4235 => "0001011000100000100000",
			4236 => "0010010110101100011100",
			4237 => "0001101010111100001000",
			4238 => "0000001110110000000100",
			4239 => "0000000100001001111001",
			4240 => "0000000100001001111001",
			4241 => "0000010111100100000100",
			4242 => "0000000100001001111001",
			4243 => "0001011011000000001000",
			4244 => "0000001010111000000100",
			4245 => "0000000100001001111001",
			4246 => "0000000100001001111001",
			4247 => "0011011001000100000100",
			4248 => "0000000100001001111001",
			4249 => "0000000100001001111001",
			4250 => "0000000100001001111001",
			4251 => "0000110001001000000100",
			4252 => "0000000100001001111001",
			4253 => "0000000100001001111001",
			4254 => "0010000101101100000100",
			4255 => "1111111100001100010101",
			4256 => "0000001101011000110100",
			4257 => "0010100000111100100100",
			4258 => "0000000110111100010100",
			4259 => "0000011100101000010000",
			4260 => "0011101110100100001000",
			4261 => "0011000101101100000100",
			4262 => "0000000100001100010101",
			4263 => "1111111100001100010101",
			4264 => "0000101011010000000100",
			4265 => "1111111100001100010101",
			4266 => "0000000100001100010101",
			4267 => "0000001100001100010101",
			4268 => "0011111100111100000100",
			4269 => "1111111100001100010101",
			4270 => "0001100100100000000100",
			4271 => "0000000100001100010101",
			4272 => "0011010101101100000100",
			4273 => "1111111100001100010101",
			4274 => "0000000100001100010101",
			4275 => "0000001100100100000100",
			4276 => "1111111100001100010101",
			4277 => "0000001110110000001000",
			4278 => "0001101010101100000100",
			4279 => "0000001100001100010101",
			4280 => "1111111100001100010101",
			4281 => "0000001100001100010101",
			4282 => "0010101011000000001100",
			4283 => "0000010101010100001000",
			4284 => "0000010011110000000100",
			4285 => "0000000100001100010101",
			4286 => "0000001100001100010101",
			4287 => "0000000100001100010101",
			4288 => "0000111011111000000100",
			4289 => "1111111100001100010101",
			4290 => "0001001101001000000100",
			4291 => "0000001100001100010101",
			4292 => "0000000100001100010101",
			4293 => "0010101101001000001000",
			4294 => "0000100101101000000100",
			4295 => "0000000100001111000001",
			4296 => "0000000100001111000001",
			4297 => "0001011001010000011100",
			4298 => "0010001001000100010000",
			4299 => "0001011000000000001000",
			4300 => "0011100010110100000100",
			4301 => "0000000100001111000001",
			4302 => "0000000100001111000001",
			4303 => "0000001001101000000100",
			4304 => "0000000100001111000001",
			4305 => "0000000100001111000001",
			4306 => "0000111001010000001000",
			4307 => "0000001011011000000100",
			4308 => "0000000100001111000001",
			4309 => "0000000100001111000001",
			4310 => "0000000100001111000001",
			4311 => "0000010111011100101100",
			4312 => "0011011100101000010100",
			4313 => "0000010110001100010000",
			4314 => "0011000011010000001000",
			4315 => "0000010111100100000100",
			4316 => "0000000100001111000001",
			4317 => "0000000100001111000001",
			4318 => "0011100100101000000100",
			4319 => "0000000100001111000001",
			4320 => "0000000100001111000001",
			4321 => "0000000100001111000001",
			4322 => "0010111001001000001000",
			4323 => "0001001000000100000100",
			4324 => "0000000100001111000001",
			4325 => "0000000100001111000001",
			4326 => "0011000110000000001000",
			4327 => "0011100100101000000100",
			4328 => "0000000100001111000001",
			4329 => "0000000100001111000001",
			4330 => "0001010011000100000100",
			4331 => "0000000100001111000001",
			4332 => "0000000100001111000001",
			4333 => "0011011101101000000100",
			4334 => "0000000100001111000001",
			4335 => "0000000100001111000001",
			4336 => "0010011000000101000100",
			4337 => "0010111001001000111000",
			4338 => "0000101110101000110000",
			4339 => "0011110010101000011100",
			4340 => "0001101010111100010000",
			4341 => "0001100101100000001000",
			4342 => "0000010011110000000100",
			4343 => "0000000100010010011101",
			4344 => "0000000100010010011101",
			4345 => "0000101011100100000100",
			4346 => "1111111100010010011101",
			4347 => "0000000100010010011101",
			4348 => "0000000100010100000100",
			4349 => "1111111100010010011101",
			4350 => "0010101011000000000100",
			4351 => "0000001100010010011101",
			4352 => "0000000100010010011101",
			4353 => "0000001101011000001100",
			4354 => "0011101000101100000100",
			4355 => "1111111100010010011101",
			4356 => "0011110011111100000100",
			4357 => "0000000100010010011101",
			4358 => "1111111100010010011101",
			4359 => "0000111001010100000100",
			4360 => "0000000100010010011101",
			4361 => "0000000100010010011101",
			4362 => "0001101011000100000100",
			4363 => "0000001100010010011101",
			4364 => "0000000100010010011101",
			4365 => "0001011001010000001000",
			4366 => "0001010110000000000100",
			4367 => "0000000100010010011101",
			4368 => "0000000100010010011101",
			4369 => "1111111100010010011101",
			4370 => "0001010011000100011100",
			4371 => "0001111110001100011000",
			4372 => "0000111000000000001100",
			4373 => "0011011001001000001000",
			4374 => "0010000000110000000100",
			4375 => "0000000100010010011101",
			4376 => "0000000100010010011101",
			4377 => "1111111100010010011101",
			4378 => "0011101111010100000100",
			4379 => "0000000100010010011101",
			4380 => "0001011011111000000100",
			4381 => "0000000100010010011101",
			4382 => "0000001100010010011101",
			4383 => "1111111100010010011101",
			4384 => "0000110000111000001000",
			4385 => "0000001111010000000100",
			4386 => "1111111100010010011101",
			4387 => "0000000100010010011101",
			4388 => "0000001101110100000100",
			4389 => "0000000100010010011101",
			4390 => "0000001100010010011101",
			4391 => "0000011101000000110100",
			4392 => "0010110111011100101100",
			4393 => "0011100100010000100000",
			4394 => "0010111110011000001100",
			4395 => "0011011011101100000100",
			4396 => "0000000100010110010001",
			4397 => "0000000100011000000100",
			4398 => "0000000100010110010001",
			4399 => "0000000100010110010001",
			4400 => "0011001110011000000100",
			4401 => "0000000100010110010001",
			4402 => "0001001100000000001000",
			4403 => "0001011100000000000100",
			4404 => "0000000100010110010001",
			4405 => "0000000100010110010001",
			4406 => "0010011101101000000100",
			4407 => "0000000100010110010001",
			4408 => "0000000100010110010001",
			4409 => "0010000101101100000100",
			4410 => "0000000100010110010001",
			4411 => "0000000100010100000100",
			4412 => "0000000100010110010001",
			4413 => "0000000100010110010001",
			4414 => "0010000011001000000100",
			4415 => "0000000100010110010001",
			4416 => "0000000100010110010001",
			4417 => "0010111001001000011000",
			4418 => "0011000101101100010100",
			4419 => "0000111001010100001100",
			4420 => "0011110101111100001000",
			4421 => "0001011000000000000100",
			4422 => "0000000100010110010001",
			4423 => "0000000100010110010001",
			4424 => "0000000100010110010001",
			4425 => "0010110101011100000100",
			4426 => "0000000100010110010001",
			4427 => "0000000100010110010001",
			4428 => "0000000100010110010001",
			4429 => "0011100110111000010100",
			4430 => "0000111100110000001000",
			4431 => "0000010011010000000100",
			4432 => "0000000100010110010001",
			4433 => "0000000100010110010001",
			4434 => "0000011011101100001000",
			4435 => "0000010110001100000100",
			4436 => "0000000100010110010001",
			4437 => "0000000100010110010001",
			4438 => "0000000100010110010001",
			4439 => "0011101010001000001000",
			4440 => "0010100011000100000100",
			4441 => "0000000100010110010001",
			4442 => "0000000100010110010001",
			4443 => "0000010111011100001000",
			4444 => "0001010011000100000100",
			4445 => "0000000100010110010001",
			4446 => "0000000100010110010001",
			4447 => "0000011100101000000100",
			4448 => "0000000100010110010001",
			4449 => "0011110011111100000100",
			4450 => "0000000100010110010001",
			4451 => "0000000100010110010001",
			4452 => "0011100001100001010000",
			4453 => "0001001100000000101000",
			4454 => "0001000011001000100100",
			4455 => "0011011101101000100000",
			4456 => "0000011001100000010000",
			4457 => "0011110011101100001000",
			4458 => "0000111100010000000100",
			4459 => "0000000100011001010101",
			4460 => "0000000100011001010101",
			4461 => "0011100011101000000100",
			4462 => "0000000100011001010101",
			4463 => "0000000100011001010101",
			4464 => "0011100100101000001000",
			4465 => "0001101100000100000100",
			4466 => "0000000100011001010101",
			4467 => "0000000100011001010101",
			4468 => "0011100010110100000100",
			4469 => "0000000100011001010101",
			4470 => "0000000100011001010101",
			4471 => "0000000100011001010101",
			4472 => "0000000100011001010101",
			4473 => "0010000011100100011000",
			4474 => "0011001101101000010100",
			4475 => "0000000010100100001000",
			4476 => "0001011011000000000100",
			4477 => "0000000100011001010101",
			4478 => "0000000100011001010101",
			4479 => "0010010011000000001000",
			4480 => "0000111011111000000100",
			4481 => "0000000100011001010101",
			4482 => "0000000100011001010101",
			4483 => "0000001100011001010101",
			4484 => "0000000100011001010101",
			4485 => "0011011010000100000100",
			4486 => "0000000100011001010101",
			4487 => "0010001100110000000100",
			4488 => "0000000100011001010101",
			4489 => "0000001011001100000100",
			4490 => "0000000100011001010101",
			4491 => "0000000100011001010101",
			4492 => "0000011100101000001100",
			4493 => "0011110100110100000100",
			4494 => "0000000100011001010101",
			4495 => "0000101101011000000100",
			4496 => "0000000100011001010101",
			4497 => "0000000100011001010101",
			4498 => "0000111001010000000100",
			4499 => "0000000100011001010101",
			4500 => "0000000100011001010101",
			4501 => "0010001010000100110000",
			4502 => "0000100101010000101100",
			4503 => "0001101100000100100000",
			4504 => "0011101001011100001100",
			4505 => "0010111011101100001000",
			4506 => "0010110110001100000100",
			4507 => "0000000100011101001001",
			4508 => "0000000100011101001001",
			4509 => "0000000100011101001001",
			4510 => "0001101110010000001100",
			4511 => "0010101100010000000100",
			4512 => "0000000100011101001001",
			4513 => "0010110111011100000100",
			4514 => "0000000100011101001001",
			4515 => "0000000100011101001001",
			4516 => "0011111110000100000100",
			4517 => "0000000100011101001001",
			4518 => "0000000100011101001001",
			4519 => "0001001100000000001000",
			4520 => "0001111100110000000100",
			4521 => "0000000100011101001001",
			4522 => "0000000100011101001001",
			4523 => "0000000100011101001001",
			4524 => "0000000100011101001001",
			4525 => "0010111001001000011100",
			4526 => "0000100110010100010000",
			4527 => "0001100100000100001100",
			4528 => "0001001000000100001000",
			4529 => "0001011101001000000100",
			4530 => "0000000100011101001001",
			4531 => "0000000100011101001001",
			4532 => "0000000100011101001001",
			4533 => "0000000100011101001001",
			4534 => "0001011000100000001000",
			4535 => "0011010101011100000100",
			4536 => "0000000100011101001001",
			4537 => "0000000100011101001001",
			4538 => "0000000100011101001001",
			4539 => "0011100110111000010000",
			4540 => "0000111100110000001000",
			4541 => "0010001000000000000100",
			4542 => "0000000100011101001001",
			4543 => "0000000100011101001001",
			4544 => "0010101111100100000100",
			4545 => "0000000100011101001001",
			4546 => "0000000100011101001001",
			4547 => "0011101010001000001000",
			4548 => "0010100011000100000100",
			4549 => "0000000100011101001001",
			4550 => "0000000100011101001001",
			4551 => "0000010111011100001100",
			4552 => "0011000110000000000100",
			4553 => "0000000100011101001001",
			4554 => "0000010011010000000100",
			4555 => "0000000100011101001001",
			4556 => "0000000100011101001001",
			4557 => "0000011100101000000100",
			4558 => "0000000100011101001001",
			4559 => "0010010110101100000100",
			4560 => "0000000100011101001001",
			4561 => "0000000100011101001001",
			4562 => "0010000101101100000100",
			4563 => "1111111100011111100101",
			4564 => "0011000101010100100000",
			4565 => "0000011101000000011000",
			4566 => "0001001010000100010000",
			4567 => "0010111010100100001100",
			4568 => "0000000100010100001000",
			4569 => "0000111100010000000100",
			4570 => "1111111100011111100101",
			4571 => "0000000100011111100101",
			4572 => "0000001100011111100101",
			4573 => "1111111100011111100101",
			4574 => "0001101000101100000100",
			4575 => "0000001100011111100101",
			4576 => "0000000100011111100101",
			4577 => "0000001101001100000100",
			4578 => "1111111100011111100101",
			4579 => "0000001100011111100101",
			4580 => "0011011100101000010100",
			4581 => "0000010110001100010000",
			4582 => "0001100010000100001100",
			4583 => "0000111000000000001000",
			4584 => "0010110101010100000100",
			4585 => "0000000100011111100101",
			4586 => "1111111100011111100101",
			4587 => "1111111100011111100101",
			4588 => "0000000100011111100101",
			4589 => "0000000100011111100101",
			4590 => "0011001111011000010100",
			4591 => "0001001001000100000100",
			4592 => "1111111100011111100101",
			4593 => "0001000011000000001000",
			4594 => "0001111000100000000100",
			4595 => "0000000100011111100101",
			4596 => "0000001100011111100101",
			4597 => "0010000011001000000100",
			4598 => "0000001100011111100101",
			4599 => "0000000100011111100101",
			4600 => "1111111100011111100101",
			4601 => "0000011101000000101000",
			4602 => "0001111100110000001100",
			4603 => "0011100011010100001000",
			4604 => "0001111100010000000100",
			4605 => "0000000100100010110001",
			4606 => "0000000100100010110001",
			4607 => "0000000100100010110001",
			4608 => "0010000011001000011000",
			4609 => "0011011100101000010000",
			4610 => "0001100011011000000100",
			4611 => "0000000100100010110001",
			4612 => "0000110011000000000100",
			4613 => "0000000100100010110001",
			4614 => "0011100100110000000100",
			4615 => "0000000100100010110001",
			4616 => "0000000100100010110001",
			4617 => "0000111011111000000100",
			4618 => "0000000100100010110001",
			4619 => "0000000100100010110001",
			4620 => "0000000100100010110001",
			4621 => "0011000101011100001100",
			4622 => "0010111010100100001000",
			4623 => "0001011000111000000100",
			4624 => "0000000100100010110001",
			4625 => "0000000100100010110001",
			4626 => "0000000100100010110001",
			4627 => "0010010101111000000100",
			4628 => "0000000100100010110001",
			4629 => "0010000011100100010100",
			4630 => "0001110001011000001100",
			4631 => "0000001000010000001000",
			4632 => "0001001101101000000100",
			4633 => "0000000100100010110001",
			4634 => "0000000100100010110001",
			4635 => "0000000100100010110001",
			4636 => "0000001100100100000100",
			4637 => "0000000100100010110001",
			4638 => "0000000100100010110001",
			4639 => "0000111001010000001100",
			4640 => "0000101111001100001000",
			4641 => "0010101001010100000100",
			4642 => "0000000100100010110001",
			4643 => "0000000100100010110001",
			4644 => "0000000100100010110001",
			4645 => "0010100000111100001000",
			4646 => "0000100010101100000100",
			4647 => "0000000100100010110001",
			4648 => "0000000100100010110001",
			4649 => "0001101110000100000100",
			4650 => "0000000100100010110001",
			4651 => "0000000100100010110001",
			4652 => "0001011000000000010100",
			4653 => "0001111100010000001000",
			4654 => "0001111000111000000100",
			4655 => "0000000100100110001101",
			4656 => "0000000100100110001101",
			4657 => "0001000110000000001000",
			4658 => "0011101000110100000100",
			4659 => "0000000100100110001101",
			4660 => "0000000100100110001101",
			4661 => "0000000100100110001101",
			4662 => "0010110111011100100000",
			4663 => "0000110100101100011100",
			4664 => "0010001001000100010000",
			4665 => "0000001010111000001100",
			4666 => "0000001011110100001000",
			4667 => "0000000011101000000100",
			4668 => "0000000100100110001101",
			4669 => "0000000100100110001101",
			4670 => "0000000100100110001101",
			4671 => "0000000100100110001101",
			4672 => "0000001101001100000100",
			4673 => "0000000100100110001101",
			4674 => "0011100101000000000100",
			4675 => "0000000100100110001101",
			4676 => "0000000100100110001101",
			4677 => "0000000100100110001101",
			4678 => "0010000000110000010000",
			4679 => "0001011100110000000100",
			4680 => "0000000100100110001101",
			4681 => "0001001000111000000100",
			4682 => "0000000100100110001101",
			4683 => "0010010101111000000100",
			4684 => "0000000100100110001101",
			4685 => "0000000100100110001101",
			4686 => "0000101111001100011100",
			4687 => "0010100000111100010000",
			4688 => "0001000011000000001000",
			4689 => "0011101111010100000100",
			4690 => "0000000100100110001101",
			4691 => "0000000100100110001101",
			4692 => "0010000011001000000100",
			4693 => "0000000100100110001101",
			4694 => "0000000100100110001101",
			4695 => "0000001100100100000100",
			4696 => "0000000100100110001101",
			4697 => "0001111100011100000100",
			4698 => "0000000100100110001101",
			4699 => "0000000100100110001101",
			4700 => "0000010101011100001000",
			4701 => "0000111111101000000100",
			4702 => "0000000100100110001101",
			4703 => "0000000100100110001101",
			4704 => "0011110011100000000100",
			4705 => "0000000100100110001101",
			4706 => "0000000100100110001101",
			4707 => "0010001010000101001000",
			4708 => "0010111011101100010100",
			4709 => "0011010110110100000100",
			4710 => "1111111100101010001001",
			4711 => "0011100110111000001100",
			4712 => "0010001111111100000100",
			4713 => "0000000100101010001001",
			4714 => "0001100001010100000100",
			4715 => "0000000100101010001001",
			4716 => "0000001100101010001001",
			4717 => "0000000100101010001001",
			4718 => "0001011001010000011000",
			4719 => "0010011101101000010000",
			4720 => "0000001101011000001100",
			4721 => "0000010011110000000100",
			4722 => "1111111100101010001001",
			4723 => "0001101000110100000100",
			4724 => "0000001100101010001001",
			4725 => "1111111100101010001001",
			4726 => "0000000100101010001001",
			4727 => "0001000110000000000100",
			4728 => "0000000100101010001001",
			4729 => "0000001100101010001001",
			4730 => "0001110110011100010100",
			4731 => "0001010011000100001000",
			4732 => "0010011001001000000100",
			4733 => "0000000100101010001001",
			4734 => "1111111100101010001001",
			4735 => "0010111010100100001000",
			4736 => "0010101001011000000100",
			4737 => "0000000100101010001001",
			4738 => "0000000100101010001001",
			4739 => "1111111100101010001001",
			4740 => "0001110011000100000100",
			4741 => "0000000100101010001001",
			4742 => "1111111100101010001001",
			4743 => "0001111011000000011000",
			4744 => "0011000101101100010100",
			4745 => "0000100110111100010000",
			4746 => "0001001100000000001100",
			4747 => "0001111100110000001000",
			4748 => "0000000100111000000100",
			4749 => "0000000100101010001001",
			4750 => "0000001100101010001001",
			4751 => "0000000100101010001001",
			4752 => "0000001100101010001001",
			4753 => "0000001100101010001001",
			4754 => "1111111100101010001001",
			4755 => "0000111100010000001000",
			4756 => "0000010011010000000100",
			4757 => "0000000100101010001001",
			4758 => "0000001100101010001001",
			4759 => "0001011011111000000100",
			4760 => "1111111100101010001001",
			4761 => "0000101011010000000100",
			4762 => "1111111100101010001001",
			4763 => "0010011000000100001000",
			4764 => "0000111011111000000100",
			4765 => "0000000100101010001001",
			4766 => "0000000100101010001001",
			4767 => "0001010011000100000100",
			4768 => "0000001100101010001001",
			4769 => "0000000100101010001001",
			4770 => "0000010111100100000100",
			4771 => "1111111100101100100101",
			4772 => "0000100101010001000000",
			4773 => "0010001111001000010100",
			4774 => "0011001010100100001100",
			4775 => "0001111101001000001000",
			4776 => "0011011011101100000100",
			4777 => "0000000100101100100101",
			4778 => "0000000100101100100101",
			4779 => "0000000100101100100101",
			4780 => "0000011101000000000100",
			4781 => "1111111100101100100101",
			4782 => "0000000100101100100101",
			4783 => "0010001000000000011100",
			4784 => "0001011001010000001100",
			4785 => "0001011000000000000100",
			4786 => "0000000100101100100101",
			4787 => "0011010011010000000100",
			4788 => "0000000100101100100101",
			4789 => "0000000100101100100101",
			4790 => "0000111000101000001000",
			4791 => "0011110101111100000100",
			4792 => "0000000100101100100101",
			4793 => "0000000100101100100101",
			4794 => "0000010110001100000100",
			4795 => "0000000100101100100101",
			4796 => "0000000100101100100101",
			4797 => "0000001110110000000100",
			4798 => "1111111100101100100101",
			4799 => "0011001010000100000100",
			4800 => "0000000100101100100101",
			4801 => "0010010110101100000100",
			4802 => "0000000100101100100101",
			4803 => "0000000100101100100101",
			4804 => "0011010011000000001000",
			4805 => "0011100001111000000100",
			4806 => "0000001100101100100101",
			4807 => "0000000100101100100101",
			4808 => "0000000100101100100101",
			4809 => "0001010011001000000100",
			4810 => "1111111100101111011001",
			4811 => "0001011001010000100000",
			4812 => "0010001001000100001100",
			4813 => "0000010011110000001000",
			4814 => "0000001010111000000100",
			4815 => "1111111100101111011001",
			4816 => "0000000100101111011001",
			4817 => "0000000100101111011001",
			4818 => "0000111100110000010000",
			4819 => "0010101000111000001000",
			4820 => "0011010111011100000100",
			4821 => "0000000100101111011001",
			4822 => "1111111100101111011001",
			4823 => "0011111011110100000100",
			4824 => "0000000100101111011001",
			4825 => "0000001100101111011001",
			4826 => "0000000100101111011001",
			4827 => "0010001010000100011000",
			4828 => "0010111011101100000100",
			4829 => "0000000100101111011001",
			4830 => "0001110110011100001100",
			4831 => "0001010011000100000100",
			4832 => "1111111100101111011001",
			4833 => "0001001100110000000100",
			4834 => "0000000100101111011001",
			4835 => "0000000100101111011001",
			4836 => "0001110011000100000100",
			4837 => "0000000100101111011001",
			4838 => "0000000100101111011001",
			4839 => "0010110101010100001000",
			4840 => "0000001000010000000100",
			4841 => "0000000100101111011001",
			4842 => "0000001100101111011001",
			4843 => "0011011100101000001000",
			4844 => "0001101110001000000100",
			4845 => "1111111100101111011001",
			4846 => "0000000100101111011001",
			4847 => "0001011011111000001000",
			4848 => "0000111001010000000100",
			4849 => "0000000100101111011001",
			4850 => "1111111100101111011001",
			4851 => "0001011100101100000100",
			4852 => "0000001100101111011001",
			4853 => "0000000100101111011001",
			4854 => "0010000101101100000100",
			4855 => "1111111100110001011101",
			4856 => "0011110010110000000100",
			4857 => "1111111100110001011101",
			4858 => "0010110111011100011000",
			4859 => "0001000101010100001000",
			4860 => "0011011110011000000100",
			4861 => "0000000100110001011101",
			4862 => "1111111100110001011101",
			4863 => "0010001001000100000100",
			4864 => "0000000100110001011101",
			4865 => "0011010111011100001000",
			4866 => "0011011010100100000100",
			4867 => "0000001100110001011101",
			4868 => "0000001100110001011101",
			4869 => "0000000100110001011101",
			4870 => "0010000000110000010000",
			4871 => "0010100001011100001100",
			4872 => "0001101110010000001000",
			4873 => "0011100011010100000100",
			4874 => "1111111100110001011101",
			4875 => "0000000100110001011101",
			4876 => "1111111100110001011101",
			4877 => "0000001100110001011101",
			4878 => "0011010101111000010000",
			4879 => "0000101111001100001000",
			4880 => "0010100000111100000100",
			4881 => "0000000100110001011101",
			4882 => "0000001100110001011101",
			4883 => "0001011000100000000100",
			4884 => "0000001100110001011101",
			4885 => "0000000100110001011101",
			4886 => "1111111100110001011101",
			4887 => "0001110011110101100100",
			4888 => "0010001010000100110000",
			4889 => "0011000101010100101000",
			4890 => "0001001111011000011100",
			4891 => "0000010011110000010000",
			4892 => "0011111000100100001000",
			4893 => "0010111011101100000100",
			4894 => "0000000100110101000001",
			4895 => "1111111100110101000001",
			4896 => "0010010101011100000100",
			4897 => "0000000100110101000001",
			4898 => "0000000100110101000001",
			4899 => "0001101010001000000100",
			4900 => "0000000100110101000001",
			4901 => "0011100001100000000100",
			4902 => "0000000100110101000001",
			4903 => "0000000100110101000001",
			4904 => "0001101111110000000100",
			4905 => "0000000100110101000001",
			4906 => "0001011000100000000100",
			4907 => "0000000100110101000001",
			4908 => "0000000100110101000001",
			4909 => "0010110011010000000100",
			4910 => "0000000100110101000001",
			4911 => "1111111100110101000001",
			4912 => "0000000110101000011100",
			4913 => "0000101100010100010100",
			4914 => "0010101001010100001100",
			4915 => "0000110011000000001000",
			4916 => "0001001100101000000100",
			4917 => "0000000100110101000001",
			4918 => "0000000100110101000001",
			4919 => "0000000100110101000001",
			4920 => "0001011100101100000100",
			4921 => "0000000100110101000001",
			4922 => "0000000100110101000001",
			4923 => "0010101011000000000100",
			4924 => "0000000100110101000001",
			4925 => "0000000100110101000001",
			4926 => "0001001010000100000100",
			4927 => "0000000100110101000001",
			4928 => "0001000011000000000100",
			4929 => "0000001100110101000001",
			4930 => "0001111001011000001000",
			4931 => "0000001010010100000100",
			4932 => "0000000100110101000001",
			4933 => "0000000100110101000001",
			4934 => "0010110110000000000100",
			4935 => "0000000100110101000001",
			4936 => "0000000100110101000001",
			4937 => "0011000011000000000100",
			4938 => "0000000100110101000001",
			4939 => "0000001010010000000100",
			4940 => "0000000100110101000001",
			4941 => "0000101001101000000100",
			4942 => "0000000100110101000001",
			4943 => "0000000100110101000001",
			4944 => "0010001111111100000100",
			4945 => "1111111100110111101101",
			4946 => "0010111011101100001100",
			4947 => "0001010011001000000100",
			4948 => "1111111100110111101101",
			4949 => "0001110110101100000100",
			4950 => "0000001100110111101101",
			4951 => "0000000100110111101101",
			4952 => "0010001010000100100100",
			4953 => "0001011001010000010100",
			4954 => "0001001001000100001000",
			4955 => "0011111000100100000100",
			4956 => "1111111100110111101101",
			4957 => "0000000100110111101101",
			4958 => "0000010011110000001000",
			4959 => "0010111010100100000100",
			4960 => "0000000100110111101101",
			4961 => "1111111100110111101101",
			4962 => "0000001100110111101101",
			4963 => "0001110110011100001000",
			4964 => "0010010101101100000100",
			4965 => "0000000100110111101101",
			4966 => "1111111100110111101101",
			4967 => "0001110011000100000100",
			4968 => "0000000100110111101101",
			4969 => "1111111100110111101101",
			4970 => "0011000101010100001000",
			4971 => "0000001101001100000100",
			4972 => "0000000100110111101101",
			4973 => "0000001100110111101101",
			4974 => "0001001001000100001100",
			4975 => "0001000011010000001000",
			4976 => "0011010101011100000100",
			4977 => "0000000100110111101101",
			4978 => "0000000100110111101101",
			4979 => "1111111100110111101101",
			4980 => "0001000011000000001000",
			4981 => "0011101111010100000100",
			4982 => "1111111100110111101101",
			4983 => "0000001100110111101101",
			4984 => "0001111100101100000100",
			4985 => "0000001100110111101101",
			4986 => "0000000100110111101101",
			4987 => "0011110010110000000100",
			4988 => "1111111100111001100001",
			4989 => "0010001111111100000100",
			4990 => "1111111100111001100001",
			4991 => "0001111100110000000100",
			4992 => "0000001100111001100001",
			4993 => "0000100100010100010100",
			4994 => "0010001000000000010000",
			4995 => "0001101000110100001000",
			4996 => "0011111100111000000100",
			4997 => "0000000100111001100001",
			4998 => "0000001100111001100001",
			4999 => "0001001100000000000100",
			5000 => "1111111100111001100001",
			5001 => "0000000100111001100001",
			5002 => "1111111100111001100001",
			5003 => "0010101111101000001100",
			5004 => "0000111100110000001000",
			5005 => "0001000110000000000100",
			5006 => "0000000100111001100001",
			5007 => "0000001100111001100001",
			5008 => "1111111100111001100001",
			5009 => "0001000011000000001000",
			5010 => "0010001010000100000100",
			5011 => "0000000100111001100001",
			5012 => "0000001100111001100001",
			5013 => "0010001100110000000100",
			5014 => "0000000100111001100001",
			5015 => "0000001100111001100001",
			5016 => "0000101010010001011100",
			5017 => "0001100111010001001100",
			5018 => "0011000101010100011100",
			5019 => "0010001001000100010000",
			5020 => "0010111011101100001000",
			5021 => "0010011100101000000100",
			5022 => "0000000100111100011101",
			5023 => "0000000100111100011101",
			5024 => "0001111011111000000100",
			5025 => "0000000100111100011101",
			5026 => "0000000100111100011101",
			5027 => "0000001101001100000100",
			5028 => "0000000100111100011101",
			5029 => "0011111011010100000100",
			5030 => "0000000100111100011101",
			5031 => "0000000100111100011101",
			5032 => "0010100000111100100000",
			5033 => "0001111000100000010000",
			5034 => "0000000110111100001000",
			5035 => "0000001111101100000100",
			5036 => "0000000100111100011101",
			5037 => "0000000100111100011101",
			5038 => "0010000011001000000100",
			5039 => "0000000100111100011101",
			5040 => "0000000100111100011101",
			5041 => "0010001000000000001000",
			5042 => "0011100110111000000100",
			5043 => "0000000100111100011101",
			5044 => "0000000100111100011101",
			5045 => "0010001001010100000100",
			5046 => "0000000100111100011101",
			5047 => "0000000100111100011101",
			5048 => "0000000101101000001100",
			5049 => "0011110111010000001000",
			5050 => "0000100010100100000100",
			5051 => "0000000100111100011101",
			5052 => "0000000100111100011101",
			5053 => "0000000100111100011101",
			5054 => "0000000100111100011101",
			5055 => "0011110100110100000100",
			5056 => "0000000100111100011101",
			5057 => "0000011100101000000100",
			5058 => "0000000100111100011101",
			5059 => "0000011111001000000100",
			5060 => "0000000100111100011101",
			5061 => "0000000100111100011101",
			5062 => "0000000100111100011101",
			5063 => "0011010101111001101100",
			5064 => "0000010110001101000000",
			5065 => "0011000101010100100100",
			5066 => "0000011101000000100000",
			5067 => "0010111110011000010000",
			5068 => "0011010110001100001000",
			5069 => "0001011000111000000100",
			5070 => "0000000100111111111001",
			5071 => "0000000100111111111001",
			5072 => "0000000100011000000100",
			5073 => "0000000100111111111001",
			5074 => "0000000100111111111001",
			5075 => "0011100100101000001000",
			5076 => "0000110011100100000100",
			5077 => "0000000100111111111001",
			5078 => "1111111100111111111001",
			5079 => "0011011010100100000100",
			5080 => "0000000100111111111001",
			5081 => "0000001100111111111001",
			5082 => "0000000100111111111001",
			5083 => "0011011100101000001100",
			5084 => "0011110101000100001000",
			5085 => "0010110011010000000100",
			5086 => "0000000100111111111001",
			5087 => "1111111100111111111001",
			5088 => "0000000100111111111001",
			5089 => "0010010011001000001000",
			5090 => "0000111000000000000100",
			5091 => "0000000100111111111001",
			5092 => "0000001100111111111001",
			5093 => "0001111100011100000100",
			5094 => "0000000100111111111001",
			5095 => "0000000100111111111001",
			5096 => "0001111001011000010000",
			5097 => "0010010011000000001000",
			5098 => "0001011001010100000100",
			5099 => "0000000100111111111001",
			5100 => "0000000100111111111001",
			5101 => "0011110100001000000100",
			5102 => "0000000100111111111001",
			5103 => "0000001100111111111001",
			5104 => "0001010011000100010000",
			5105 => "0001010110011100001100",
			5106 => "0000001110101000001000",
			5107 => "0001001111011000000100",
			5108 => "0000000100111111111001",
			5109 => "1111111100111111111001",
			5110 => "0000000100111111111001",
			5111 => "0000001100111111111001",
			5112 => "0000110000111100001000",
			5113 => "0000001101011000000100",
			5114 => "1111111100111111111001",
			5115 => "0000000100111111111001",
			5116 => "0000000100111111111001",
			5117 => "1111111100111111111001",
			5118 => "0010000101101100000100",
			5119 => "1111111101000011011111",
			5120 => "0011000101010100100100",
			5121 => "0001010011001000001000",
			5122 => "0010001001000100000100",
			5123 => "0000000101000011011111",
			5124 => "1111111101000011011111",
			5125 => "0000011101000000010100",
			5126 => "0010111110011000001000",
			5127 => "0001000101101100000100",
			5128 => "0000000101000011011111",
			5129 => "0000001101000011011111",
			5130 => "0011100100101000001000",
			5131 => "0000110011100100000100",
			5132 => "0000000101000011011111",
			5133 => "1111111101000011011111",
			5134 => "0000001101000011011111",
			5135 => "0000001101001100000100",
			5136 => "0000000101000011011111",
			5137 => "0000001101000011011111",
			5138 => "0010000000110000011100",
			5139 => "0010010110000000001000",
			5140 => "0010001001000100000100",
			5141 => "1111111101000011011111",
			5142 => "0000000101000011011111",
			5143 => "0010100001011100001100",
			5144 => "0000111000000000001000",
			5145 => "0000110011001000000100",
			5146 => "1111111101000011011111",
			5147 => "0000000101000011011111",
			5148 => "1111111101000011011111",
			5149 => "0001111011000000000100",
			5150 => "0000001101000011011111",
			5151 => "0000000101000011011111",
			5152 => "0001001001000100010000",
			5153 => "0001000011010000001100",
			5154 => "0001001010100100000100",
			5155 => "0000000101000011011111",
			5156 => "0000010110001100000100",
			5157 => "0000000101000011011111",
			5158 => "0000000101000011011111",
			5159 => "1111111101000011011111",
			5160 => "0001011001011000010000",
			5161 => "0011111100111100001000",
			5162 => "0011111110101100000100",
			5163 => "0000001101000011011111",
			5164 => "0000000101000011011111",
			5165 => "0001011011111000000100",
			5166 => "0000000101000011011111",
			5167 => "0000001101000011011111",
			5168 => "0010100000111100001000",
			5169 => "0000001101011000000100",
			5170 => "1111111101000011011111",
			5171 => "0000000101000011011111",
			5172 => "0001110011000100000100",
			5173 => "0000001101000011011111",
			5174 => "0000000101000011011111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1711, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3455, initial_addr_3'length));
	end generate gen_rom_5;

	gen_rom_6: if SELECT_ROM = 6 generate
		bank <= (
			0 => "0011100111100000001100",
			1 => "0011011101000000001000",
			2 => "0011011111011100000100",
			3 => "0000000000000000111101",
			4 => "0000000000000000111101",
			5 => "0000000000000000111101",
			6 => "0011101100000100001000",
			7 => "0001011100110000000100",
			8 => "0000000000000000111101",
			9 => "0000000000000000111101",
			10 => "0001111100101100000100",
			11 => "0000000000000000111101",
			12 => "0001110011000100000100",
			13 => "0000000000000000111101",
			14 => "0000000000000000111101",
			15 => "0011100101000000010000",
			16 => "0011001011101100001000",
			17 => "0001001001001000000100",
			18 => "0000000000000010000001",
			19 => "0000000000000010000001",
			20 => "0001001110011000000100",
			21 => "0000000000000010000001",
			22 => "0000000000000010000001",
			23 => "0010001001000100001000",
			24 => "0001100000100100000100",
			25 => "0000000000000010000001",
			26 => "0000000000000010000001",
			27 => "0010100100101100000100",
			28 => "0000000000000010000001",
			29 => "0001001111011000000100",
			30 => "0000000000000010000001",
			31 => "0000000000000010000001",
			32 => "0011100111100000001100",
			33 => "0011001011101100001000",
			34 => "0011000110001100000100",
			35 => "0000000000000010111101",
			36 => "0000000000000010111101",
			37 => "0000000000000010111101",
			38 => "0000010111100100000100",
			39 => "0000000000000010111101",
			40 => "0001110011000100001100",
			41 => "0001011001010000001000",
			42 => "0001111011111000000100",
			43 => "0000000000000010111101",
			44 => "0000000000000010111101",
			45 => "0000000000000010111101",
			46 => "0000000000000010111101",
			47 => "0011100111100000001100",
			48 => "0011001011101100001000",
			49 => "0011000110001100000100",
			50 => "0000000000000100000001",
			51 => "0000000000000100000001",
			52 => "0000000000000100000001",
			53 => "0011100101100000010000",
			54 => "0000111000101000001100",
			55 => "0001110110011100001000",
			56 => "0001001001000100000100",
			57 => "0000000000000100000001",
			58 => "0000000000000100000001",
			59 => "0000000000000100000001",
			60 => "0000000000000100000001",
			61 => "0000111001010000000100",
			62 => "0000000000000100000001",
			63 => "0000000000000100000001",
			64 => "0011100110111000000100",
			65 => "1111111000000100111101",
			66 => "0011100010110100001000",
			67 => "0001011100010000000100",
			68 => "0000001000000100111101",
			69 => "0000000000000100111101",
			70 => "0000111100110000001000",
			71 => "0000111000000000000100",
			72 => "0000000000000100111101",
			73 => "0000000000000100111101",
			74 => "0011001010100100000100",
			75 => "0000000000000100111101",
			76 => "0001011001010000000100",
			77 => "0000001000000100111101",
			78 => "0000000000000100111101",
			79 => "0000010111100100010100",
			80 => "0001001110011000001100",
			81 => "0010001001000100001000",
			82 => "0001111100110000000100",
			83 => "0000000000000110010001",
			84 => "0000000000000110010001",
			85 => "0000000000000110010001",
			86 => "0001011101101000000100",
			87 => "0000000000000110010001",
			88 => "0000000000000110010001",
			89 => "0000110011100100001000",
			90 => "0011001011101100000100",
			91 => "0000000000000110010001",
			92 => "0000000000000110010001",
			93 => "0001011001010000001100",
			94 => "0011100101100000001000",
			95 => "0011110000001000000100",
			96 => "0000000000000110010001",
			97 => "0000000000000110010001",
			98 => "0000000000000110010001",
			99 => "0000000000000110010001",
			100 => "0001100010000100001100",
			101 => "0001100100100000000100",
			102 => "1111111000000111011101",
			103 => "0010101000101000000100",
			104 => "0000010000000111011101",
			105 => "1111111000000111011101",
			106 => "0001011001010100010100",
			107 => "0010010101010100000100",
			108 => "0000011000000111011101",
			109 => "0000001010010000001100",
			110 => "0001100111010000000100",
			111 => "0000011000000111011101",
			112 => "0011100101100000000100",
			113 => "0000010000000111011101",
			114 => "0000001000000111011101",
			115 => "1111111000000111011101",
			116 => "0000101111101100000100",
			117 => "0000000000000111011101",
			118 => "1111111000000111011101",
			119 => "0011110000100100010000",
			120 => "0001011000000100001100",
			121 => "0001000101010100000100",
			122 => "0000000000001000110001",
			123 => "0010001111111100000100",
			124 => "0000000000001000110001",
			125 => "0000000000001000110001",
			126 => "0000000000001000110001",
			127 => "0011110011100000010100",
			128 => "0000101101110000010000",
			129 => "0011011010100100001000",
			130 => "0001011000000100000100",
			131 => "0000000000001000110001",
			132 => "0000000000001000110001",
			133 => "0000111001010000000100",
			134 => "0000000000001000110001",
			135 => "0000000000001000110001",
			136 => "0000000000001000110001",
			137 => "0000111001010000000100",
			138 => "0000000000001000110001",
			139 => "0000000000001000110001",
			140 => "0010111011101100010000",
			141 => "0000000010100100000100",
			142 => "0000000000001010001101",
			143 => "0000010001110000000100",
			144 => "0000000000001010001101",
			145 => "0011001110011000000100",
			146 => "0000000000001010001101",
			147 => "0000000000001010001101",
			148 => "0000101010101000010000",
			149 => "0001000101010100001000",
			150 => "0000010110010000000100",
			151 => "0000000000001010001101",
			152 => "0000000000001010001101",
			153 => "0011110101111100000100",
			154 => "0000000000001010001101",
			155 => "0000000000001010001101",
			156 => "0000111001010000000100",
			157 => "0000000000001010001101",
			158 => "0010001001000100000100",
			159 => "0000000000001010001101",
			160 => "0000111000101000000100",
			161 => "0000000000001010001101",
			162 => "0000000000001010001101",
			163 => "0011100110111000000100",
			164 => "1111111000001011001001",
			165 => "0001110011000100011000",
			166 => "0001111011111000001100",
			167 => "0010111011101100000100",
			168 => "0000000000001011001001",
			169 => "0001011000000000000100",
			170 => "1111111000001011001001",
			171 => "0000000000001011001001",
			172 => "0001011001010000001000",
			173 => "0011011110011000000100",
			174 => "0000001000001011001001",
			175 => "0000000000001011001001",
			176 => "1111111000001011001001",
			177 => "1111111000001011001001",
			178 => "0010111011101100010000",
			179 => "0000000010100100000100",
			180 => "0000000000001100100101",
			181 => "0000010001110000000100",
			182 => "0000000000001100100101",
			183 => "0011100110111000000100",
			184 => "0000000000001100100101",
			185 => "0000000000001100100101",
			186 => "0000101010101000001100",
			187 => "0010000101101100000100",
			188 => "0000000000001100100101",
			189 => "0011110101111100000100",
			190 => "0000000000001100100101",
			191 => "0000000000001100100101",
			192 => "0001000111011100000100",
			193 => "0000000000001100100101",
			194 => "0000010110001100001000",
			195 => "0010101011000000000100",
			196 => "0000000000001100100101",
			197 => "0000000000001100100101",
			198 => "0010001111011000000100",
			199 => "0000000000001100100101",
			200 => "0000000000001100100101",
			201 => "0011110011111100100100",
			202 => "0001110100101100010100",
			203 => "0011011110011000001100",
			204 => "0011010110110100001000",
			205 => "0011011111011100000100",
			206 => "0000000000001110001001",
			207 => "0000000000001110001001",
			208 => "0000000000001110001001",
			209 => "0010010101101100000100",
			210 => "0000000000001110001001",
			211 => "0000000000001110001001",
			212 => "0011011110011000000100",
			213 => "0000000000001110001001",
			214 => "0010100100101100000100",
			215 => "0000000000001110001001",
			216 => "0001001010000100000100",
			217 => "0000000000001110001001",
			218 => "0000000000001110001001",
			219 => "0000101101011000001000",
			220 => "0001100000100100000100",
			221 => "0000000000001110001001",
			222 => "0000000000001110001001",
			223 => "0001100010101000000100",
			224 => "0000000000001110001001",
			225 => "0000000000001110001001",
			226 => "0001100000010000000100",
			227 => "1111111000001111000101",
			228 => "0001011001010000011000",
			229 => "0010111011101100001000",
			230 => "0001111000101000000100",
			231 => "0000010000001111000101",
			232 => "0000001000001111000101",
			233 => "0000110011100100000100",
			234 => "1111111000001111000101",
			235 => "0001110100101100000100",
			236 => "0000000000001111000101",
			237 => "0011011010100100000100",
			238 => "0000010000001111000101",
			239 => "0000000000001111000101",
			240 => "1111111000001111000101",
			241 => "0000111100110000100100",
			242 => "0010111011101100010100",
			243 => "0011111000100100010000",
			244 => "0011010110110100001000",
			245 => "0000010111100100000100",
			246 => "0000000000010000101001",
			247 => "0000000000010000101001",
			248 => "0010010101010100000100",
			249 => "0000000000010000101001",
			250 => "0000000000010000101001",
			251 => "0000000000010000101001",
			252 => "0000101010000000001100",
			253 => "0011011110011000001000",
			254 => "0010001001000100000100",
			255 => "0000000000010000101001",
			256 => "0000000000010000101001",
			257 => "0000000000010000101001",
			258 => "0000000000010000101001",
			259 => "0000100011011100000100",
			260 => "0000000000010000101001",
			261 => "0001011001010000001000",
			262 => "0011100110110000000100",
			263 => "0000000000010000101001",
			264 => "0000000000010000101001",
			265 => "0000000000010000101001",
			266 => "0000100011011100000100",
			267 => "0000000000010001110101",
			268 => "0000111100110000011100",
			269 => "0001111000101000001100",
			270 => "0010010101011100001000",
			271 => "0001011000000000000100",
			272 => "0000000000010001110101",
			273 => "0000000000010001110101",
			274 => "0000000000010001110101",
			275 => "0001101101010100001000",
			276 => "0000000100010100000100",
			277 => "0000000000010001110101",
			278 => "0000000000010001110101",
			279 => "0001001001000100000100",
			280 => "0000000000010001110101",
			281 => "0000000000010001110101",
			282 => "0001011001010100000100",
			283 => "0000000000010001110101",
			284 => "0000000000010001110101",
			285 => "0001100000010000000100",
			286 => "1111111000010011001001",
			287 => "0000000111111000010000",
			288 => "0001110011000100001100",
			289 => "0001001100101000001000",
			290 => "0001101101010100000100",
			291 => "0000001000010011001001",
			292 => "0000000000010011001001",
			293 => "0000001000010011001001",
			294 => "1111111000010011001001",
			295 => "0001110001010000001100",
			296 => "0010010101011100000100",
			297 => "0000001000010011001001",
			298 => "0000001110101000000100",
			299 => "0000000000010011001001",
			300 => "1111111000010011001001",
			301 => "0011101000010100001000",
			302 => "0001101011110100000100",
			303 => "1111111000010011001001",
			304 => "1111111000010011001001",
			305 => "0000000000010011001001",
			306 => "0001100100011000101100",
			307 => "0010000101101100011000",
			308 => "0010010101010100001000",
			309 => "0011010110110100000100",
			310 => "0000000000010100111101",
			311 => "0000000000010100111101",
			312 => "0011010110110100001000",
			313 => "0001000101010100000100",
			314 => "0000000000010100111101",
			315 => "0000000000010100111101",
			316 => "0010101011111000000100",
			317 => "0000000000010100111101",
			318 => "0000000000010100111101",
			319 => "0000011000011000001000",
			320 => "0011110000001000000100",
			321 => "0000000000010100111101",
			322 => "0000000000010100111101",
			323 => "0001011100010000000100",
			324 => "0000000000010100111101",
			325 => "0001010110101100000100",
			326 => "0000000000010100111101",
			327 => "0000000000010100111101",
			328 => "0010111011101100000100",
			329 => "0000000000010100111101",
			330 => "0011110111101100001000",
			331 => "0001011001010000000100",
			332 => "0000000000010100111101",
			333 => "0000000000010100111101",
			334 => "0000000000010100111101",
			335 => "0001100000010000000100",
			336 => "1111111000010110000001",
			337 => "0011000111011100011100",
			338 => "0000111100110000010000",
			339 => "0010111011101100000100",
			340 => "0000001000010110000001",
			341 => "0011111011011000001000",
			342 => "0010101001010100000100",
			343 => "1111111000010110000001",
			344 => "0000001000010110000001",
			345 => "1111111000010110000001",
			346 => "0011100110000100000100",
			347 => "0000011000010110000001",
			348 => "0001111100101100000100",
			349 => "0000000000010110000001",
			350 => "0000001000010110000001",
			351 => "1111111000010110000001",
			352 => "0001100000010000000100",
			353 => "1111111000010111011101",
			354 => "0000000111111000010100",
			355 => "0000111100110000001000",
			356 => "0011011110011000000100",
			357 => "0000001000010111011101",
			358 => "1111111000010111011101",
			359 => "0011011010100100000100",
			360 => "0000001000010111011101",
			361 => "0011111101001100000100",
			362 => "1111111000010111011101",
			363 => "0000000000010111011101",
			364 => "0001110001010000001100",
			365 => "0010010101011100000100",
			366 => "0000001000010111011101",
			367 => "0000001110101000000100",
			368 => "0000000000010111011101",
			369 => "1111111000010111011101",
			370 => "0011101000010100001000",
			371 => "0001101011110100000100",
			372 => "1111111000010111011101",
			373 => "1111111000010111011101",
			374 => "0000000000010111011101",
			375 => "0011000011010000100000",
			376 => "0001110100101100011000",
			377 => "0000101010101000000100",
			378 => "0000000000011001000001",
			379 => "0011110011100000010000",
			380 => "0011001110011000001100",
			381 => "0010001001001100000100",
			382 => "0000000000011001000001",
			383 => "0011100110110000000100",
			384 => "0000000000011001000001",
			385 => "0000000000011001000001",
			386 => "0000000000011001000001",
			387 => "0000000000011001000001",
			388 => "0010101000101000000100",
			389 => "0000000000011001000001",
			390 => "0000000000011001000001",
			391 => "0000111001010000000100",
			392 => "0000000000011001000001",
			393 => "0000111111101000001000",
			394 => "0011100010110100000100",
			395 => "0000000000011001000001",
			396 => "0000000000011001000001",
			397 => "0001101001111000000100",
			398 => "0000000000011001000001",
			399 => "0000000000011001000001",
			400 => "0000100011011100000100",
			401 => "1111111000011010011101",
			402 => "0000000111111000011100",
			403 => "0011011010100100010000",
			404 => "0000110011001000000100",
			405 => "1111111000011010011101",
			406 => "0001011001010100001000",
			407 => "0001100000010000000100",
			408 => "0000000000011010011101",
			409 => "0000001000011010011101",
			410 => "0000000000011010011101",
			411 => "0010100100101100000100",
			412 => "1111111000011010011101",
			413 => "0001001111011000000100",
			414 => "0000001000011010011101",
			415 => "0000000000011010011101",
			416 => "0010111011101100001000",
			417 => "0001011000000000000100",
			418 => "0000000000011010011101",
			419 => "1111111000011010011101",
			420 => "0001100101000100000100",
			421 => "1111111000011010011101",
			422 => "0000000000011010011101",
			423 => "0011100110110000000100",
			424 => "1111111000011100000001",
			425 => "0011011010100100011000",
			426 => "0000001010010100001100",
			427 => "0000000011011100000100",
			428 => "1111111000011100000001",
			429 => "0000111100110000000100",
			430 => "0000000000011100000001",
			431 => "0000001000011100000001",
			432 => "0010111011101100000100",
			433 => "0000000000011100000001",
			434 => "0000010110010000000100",
			435 => "0000000000011100000001",
			436 => "1111111000011100000001",
			437 => "0011100100000100001100",
			438 => "0011101100000100001000",
			439 => "0011100001100000000100",
			440 => "1111111000011100000001",
			441 => "0000000000011100000001",
			442 => "1111111000011100000001",
			443 => "0000111001010000000100",
			444 => "1111111000011100000001",
			445 => "0001001100000000000100",
			446 => "0000001000011100000001",
			447 => "0000000000011100000001",
			448 => "0000000111111000101000",
			449 => "0001011111011000010000",
			450 => "0000111100110000001100",
			451 => "0010010101010100001000",
			452 => "0001111000111000000100",
			453 => "0000000000011110000101",
			454 => "0000000000011110000101",
			455 => "0000000000011110000101",
			456 => "0000000000011110000101",
			457 => "0001011001010000010100",
			458 => "0000011000011000001100",
			459 => "0000110011100100000100",
			460 => "0000000000011110000101",
			461 => "0011110000001000000100",
			462 => "0000000000011110000101",
			463 => "0000001000011110000101",
			464 => "0001100010000100000100",
			465 => "0000000000011110000101",
			466 => "0000000000011110000101",
			467 => "0000000000011110000101",
			468 => "0001110001010000010100",
			469 => "0010010101011100001000",
			470 => "0001011000000000000100",
			471 => "0000001000011110000101",
			472 => "0000000000011110000101",
			473 => "0000111100110000000100",
			474 => "0000000000011110000101",
			475 => "0000001110110000000100",
			476 => "0000000000011110000101",
			477 => "0000000000011110000101",
			478 => "0011101000010100000100",
			479 => "1111111000011110000101",
			480 => "0000000000011110000101",
			481 => "0000111100110000101100",
			482 => "0010010101010100001100",
			483 => "0000010001110000000100",
			484 => "0000000000100000001001",
			485 => "0000110011000000000100",
			486 => "0000000000100000001001",
			487 => "0000001000100000001001",
			488 => "0000001001110100001100",
			489 => "0001111011111000000100",
			490 => "1111111000100000001001",
			491 => "0001011111011000000100",
			492 => "0000000000100000001001",
			493 => "0000001000100000001001",
			494 => "0010111011101100001000",
			495 => "0011110010101000000100",
			496 => "0000000000100000001001",
			497 => "0000000000100000001001",
			498 => "0001000110000000000100",
			499 => "1111111000100000001001",
			500 => "0001001010000100000100",
			501 => "0000000000100000001001",
			502 => "0000000000100000001001",
			503 => "0000100011011100000100",
			504 => "1111111000100000001001",
			505 => "0000000111111000001000",
			506 => "0001011001010000000100",
			507 => "0000001000100000001001",
			508 => "0000000000100000001001",
			509 => "0000010011110000001000",
			510 => "0011110100111100000100",
			511 => "0000000000100000001001",
			512 => "0000000000100000001001",
			513 => "1111111000100000001001",
			514 => "0001000101101100101100",
			515 => "0000110011001000001100",
			516 => "0010010111011100001000",
			517 => "0000000110011000000100",
			518 => "0000000000100001110101",
			519 => "0000000000100001110101",
			520 => "1111111000100001110101",
			521 => "0001101101010100011000",
			522 => "0000000100010100010100",
			523 => "0001000101010100001100",
			524 => "0001001010100100001000",
			525 => "0011010111011100000100",
			526 => "0000001000100001110101",
			527 => "0000000000100001110101",
			528 => "1111111000100001110101",
			529 => "0000000001110100000100",
			530 => "0000000000100001110101",
			531 => "0000001000100001110101",
			532 => "0000000000100001110101",
			533 => "0001111011111000000100",
			534 => "0000000000100001110101",
			535 => "0000000000100001110101",
			536 => "0011100101000000000100",
			537 => "1111111000100001110101",
			538 => "0001010100101100000100",
			539 => "0000000000100001110101",
			540 => "0000000000100001110101",
			541 => "0001011000000100010100",
			542 => "0000110011100100001000",
			543 => "0011001011101100000100",
			544 => "0000000000100011111001",
			545 => "0000000000100011111001",
			546 => "0000000010101100001000",
			547 => "0000011000011000000100",
			548 => "0000000000100011111001",
			549 => "0000000000100011111001",
			550 => "0000000000100011111001",
			551 => "0011110011100000101000",
			552 => "0011110000100100010100",
			553 => "0000010110010000001000",
			554 => "0000010111110000000100",
			555 => "0000000000100011111001",
			556 => "0000000000100011111001",
			557 => "0000111001010000000100",
			558 => "0000000000100011111001",
			559 => "0010100100101100000100",
			560 => "0000000000100011111001",
			561 => "0000000000100011111001",
			562 => "0011011010100100001000",
			563 => "0000001110110000000100",
			564 => "0000000000100011111001",
			565 => "0000000000100011111001",
			566 => "0010100100101100000100",
			567 => "0000000000100011111001",
			568 => "0001000011000000000100",
			569 => "0000000000100011111001",
			570 => "0000000000100011111001",
			571 => "0010101011111000000100",
			572 => "0000000000100011111001",
			573 => "0000000000100011111001",
			574 => "0011110000001000000100",
			575 => "1111111000100100111101",
			576 => "0000010111110000000100",
			577 => "1111111000100100111101",
			578 => "0011010110001100000100",
			579 => "0000001000100100111101",
			580 => "0000001010010000010000",
			581 => "0001110011000100001100",
			582 => "0000000011001100000100",
			583 => "0000000000100100111101",
			584 => "0011110101000100000100",
			585 => "1111111000100100111101",
			586 => "0000001000100100111101",
			587 => "1111111000100100111101",
			588 => "0001100010101000000100",
			589 => "1111111000100100111101",
			590 => "0000000000100100111101",
			591 => "0000011000011000101000",
			592 => "0000010111110000001100",
			593 => "0001001101000000000100",
			594 => "0000000000100111000001",
			595 => "0001111011111000000100",
			596 => "0000000000100111000001",
			597 => "0000000000100111000001",
			598 => "0010001001001100000100",
			599 => "0000000000100111000001",
			600 => "0010100100101100001100",
			601 => "0011110000001000000100",
			602 => "0000000000100111000001",
			603 => "0000110011100100000100",
			604 => "0000000000100111000001",
			605 => "0000000000100111000001",
			606 => "0001110100101100000100",
			607 => "0000000000100111000001",
			608 => "0010001111001000000100",
			609 => "0000000000100111000001",
			610 => "0000000000100111000001",
			611 => "0010100100101100010100",
			612 => "0010010101010100000100",
			613 => "0000000000100111000001",
			614 => "0010010101101100000100",
			615 => "0000000000100111000001",
			616 => "0010110011010000001000",
			617 => "0010001111001000000100",
			618 => "0000000000100111000001",
			619 => "0000000000100111000001",
			620 => "0000000000100111000001",
			621 => "0001011000101000000100",
			622 => "0000000000100111000001",
			623 => "0000000000100111000001",
			624 => "0000000111111000110000",
			625 => "0001110001010000010000",
			626 => "0011010110110100001000",
			627 => "0001110110101100000100",
			628 => "0000000000101001001101",
			629 => "0000000000101001001101",
			630 => "0010010101010100000100",
			631 => "0000000000101001001101",
			632 => "0000000000101001001101",
			633 => "0000110011100100000100",
			634 => "0000000000101001001101",
			635 => "0011011010100100001100",
			636 => "0000010111100100000100",
			637 => "0000000000101001001101",
			638 => "0011110000001000000100",
			639 => "0000000000101001001101",
			640 => "0000000000101001001101",
			641 => "0010001001000100000100",
			642 => "0000000000101001001101",
			643 => "0000010110001100001000",
			644 => "0010101011000000000100",
			645 => "0000000000101001001101",
			646 => "0000000000101001001101",
			647 => "0000000000101001001101",
			648 => "0001110001010000010000",
			649 => "0010010101011100001000",
			650 => "0001011000000000000100",
			651 => "0000000000101001001101",
			652 => "0000000000101001001101",
			653 => "0000000101101000000100",
			654 => "0000000000101001001101",
			655 => "0000000000101001001101",
			656 => "0011101000010100000100",
			657 => "0000000000101001001101",
			658 => "0000000000101001001101",
			659 => "0001011000000100011000",
			660 => "0000010001110000000100",
			661 => "0000000000101011101001",
			662 => "0000000010101100001000",
			663 => "0001011111011000000100",
			664 => "0000000000101011101001",
			665 => "0000000000101011101001",
			666 => "0000110011100100001000",
			667 => "0000110011000000000100",
			668 => "0000000000101011101001",
			669 => "0000000000101011101001",
			670 => "0000000000101011101001",
			671 => "0010101111101000011000",
			672 => "0010011001001000001100",
			673 => "0011110110011000001000",
			674 => "0011110111010000000100",
			675 => "0000000000101011101001",
			676 => "0000000000101011101001",
			677 => "0000000000101011101001",
			678 => "0001011100110000001000",
			679 => "0001011000111000000100",
			680 => "0000000000101011101001",
			681 => "0000000000101011101001",
			682 => "0000000000101011101001",
			683 => "0000000111111000010100",
			684 => "0011010011010000001000",
			685 => "0011110000100100000100",
			686 => "0000000000101011101001",
			687 => "0000000000101011101001",
			688 => "0000010110001100000100",
			689 => "0000000000101011101001",
			690 => "0000011011101100000100",
			691 => "0000000000101011101001",
			692 => "0000000000101011101001",
			693 => "0001110001010000001000",
			694 => "0011111101001100000100",
			695 => "0000000000101011101001",
			696 => "0000000000101011101001",
			697 => "0000000000101011101001",
			698 => "0000100011011100000100",
			699 => "1111111000101100111101",
			700 => "0001011001010000100100",
			701 => "0000111100110000011000",
			702 => "0010010101010100001000",
			703 => "0000010001110000000100",
			704 => "1111111000101100111101",
			705 => "0000001000101100111101",
			706 => "0011100001100000001100",
			707 => "0000000010101100000100",
			708 => "1111111000101100111101",
			709 => "0000100100010100000100",
			710 => "0000000000101100111101",
			711 => "1111111000101100111101",
			712 => "0000000000101100111101",
			713 => "0000001010010100001000",
			714 => "0000111001010000000100",
			715 => "0000001000101100111101",
			716 => "0000001000101100111101",
			717 => "0000000000101100111101",
			718 => "1111111000101100111101",
			719 => "0000010111100100010000",
			720 => "0001001110011000001000",
			721 => "0010000101011100000100",
			722 => "0000000000101111001001",
			723 => "0000000000101111001001",
			724 => "0001010101111000000100",
			725 => "0000000000101111001001",
			726 => "0000000000101111001001",
			727 => "0011110011100000110000",
			728 => "0011011010100100011000",
			729 => "0000001010000000001100",
			730 => "0001010011001000001000",
			731 => "0010001001000100000100",
			732 => "0000000000101111001001",
			733 => "0000000000101111001001",
			734 => "0000000000101111001001",
			735 => "0000001110110000001000",
			736 => "0011100110110000000100",
			737 => "0000000000101111001001",
			738 => "0000001000101111001001",
			739 => "0000000000101111001001",
			740 => "0010100100101100001100",
			741 => "0000100110101000000100",
			742 => "0000000000101111001001",
			743 => "0000100110100100000100",
			744 => "0000000000101111001001",
			745 => "0000000000101111001001",
			746 => "0001000011000000001000",
			747 => "0011100111100000000100",
			748 => "0000000000101111001001",
			749 => "0000000000101111001001",
			750 => "0000000000101111001001",
			751 => "0000111001010000000100",
			752 => "0000000000101111001001",
			753 => "0000000000101111001001",
			754 => "0000110011100100001100",
			755 => "0010010101010100001000",
			756 => "0001111100010000000100",
			757 => "0000000000110001001101",
			758 => "0000000000110001001101",
			759 => "1111111000110001001101",
			760 => "0000010111100100001000",
			761 => "0001011000000100000100",
			762 => "0000000000110001001101",
			763 => "0000000000110001001101",
			764 => "0000011000011000010100",
			765 => "0010100100101100001000",
			766 => "0001011100010000000100",
			767 => "0000001000110001001101",
			768 => "0000000000110001001101",
			769 => "0001110100101100000100",
			770 => "0000000000110001001101",
			771 => "0010001010000100000100",
			772 => "0000000000110001001101",
			773 => "0000000000110001001101",
			774 => "0001000111011100001000",
			775 => "0000010011110000000100",
			776 => "0000000000110001001101",
			777 => "0000000000110001001101",
			778 => "0000101010101000001000",
			779 => "0000100111011000000100",
			780 => "0000000000110001001101",
			781 => "0000000000110001001101",
			782 => "0010100100101100000100",
			783 => "0000000000110001001101",
			784 => "0001111111101000000100",
			785 => "0000000000110001001101",
			786 => "0000000000110001001101",
			787 => "0011100110110000000100",
			788 => "1111111000110010100001",
			789 => "0000110011001000000100",
			790 => "0000000000110010100001",
			791 => "0000010111110000000100",
			792 => "1111111000110010100001",
			793 => "0011011010100100001100",
			794 => "0010100100101100001000",
			795 => "0001001100101000000100",
			796 => "0000001000110010100001",
			797 => "0000000000110010100001",
			798 => "0000000000110010100001",
			799 => "0011101110001000001100",
			800 => "0010100100101100000100",
			801 => "1111111000110010100001",
			802 => "0001011011111000000100",
			803 => "0000001000110010100001",
			804 => "0000000000110010100001",
			805 => "0000000010100000000100",
			806 => "0000001000110010100001",
			807 => "0000000000110010100001",
			808 => "0000100011011100000100",
			809 => "0000000000110011111101",
			810 => "0000101101110000100100",
			811 => "0001110011000100100000",
			812 => "0000110011001000001000",
			813 => "0010010101010100000100",
			814 => "0000000000110011111101",
			815 => "0000000000110011111101",
			816 => "0000111000101000001100",
			817 => "0000010111110000000100",
			818 => "0000000000110011111101",
			819 => "0010100100101100000100",
			820 => "0000001000110011111101",
			821 => "0000000000110011111101",
			822 => "0001111100101100000100",
			823 => "0000000000110011111101",
			824 => "0000111011111000000100",
			825 => "0000000000110011111101",
			826 => "0000000000110011111101",
			827 => "0000000000110011111101",
			828 => "0011110101011000000100",
			829 => "0000000000110011111101",
			830 => "0000000000110011111101",
			831 => "0011100110111000000100",
			832 => "1111111000110101110001",
			833 => "0011101010001000001100",
			834 => "0001100100100000000100",
			835 => "0000000000110101110001",
			836 => "0000000101101000000100",
			837 => "0000001000110101110001",
			838 => "0000000000110101110001",
			839 => "0000111001010000011000",
			840 => "0011100101001100010100",
			841 => "0011111000100100001100",
			842 => "0011100001100000001000",
			843 => "0011110100111100000100",
			844 => "0000000000110101110001",
			845 => "0000000000110101110001",
			846 => "0000000000110101110001",
			847 => "0010010101011100000100",
			848 => "0000000000110101110001",
			849 => "0000000000110101110001",
			850 => "0000000000110101110001",
			851 => "0011100100000100001100",
			852 => "0011110100111100001000",
			853 => "0011100101000000000100",
			854 => "0000000000110101110001",
			855 => "0000000000110101110001",
			856 => "0000000000110101110001",
			857 => "0001001111011000000100",
			858 => "0000001000110101110001",
			859 => "0000000000110101110001",
			860 => "0011110000001000000100",
			861 => "1111111000110111001101",
			862 => "0010010101010100000100",
			863 => "0000001000110111001101",
			864 => "0000110011100100001000",
			865 => "0011011011101100000100",
			866 => "0000000000110111001101",
			867 => "1111111000110111001101",
			868 => "0000000111111000010000",
			869 => "0001100000001100000100",
			870 => "0000001000110111001101",
			871 => "0000111100110000000100",
			872 => "0000000000110111001101",
			873 => "0000111000101000000100",
			874 => "0000001000110111001101",
			875 => "0000000000110111001101",
			876 => "0000010011110000001100",
			877 => "0000001010010000001000",
			878 => "0000100000000000000100",
			879 => "0000000000110111001101",
			880 => "0000000000110111001101",
			881 => "1111111000110111001101",
			882 => "1111111000110111001101",
			883 => "0001111011111000111000",
			884 => "0010010111011100001000",
			885 => "0010100011000000000100",
			886 => "0000000000111001011001",
			887 => "0000001000111001011001",
			888 => "0001011111011000010100",
			889 => "0000111100110000010000",
			890 => "0010010101010100000100",
			891 => "0000000000111001011001",
			892 => "0000010110010000001000",
			893 => "0000010111110000000100",
			894 => "0000000000111001011001",
			895 => "0000000000111001011001",
			896 => "1111111000111001011001",
			897 => "0000000000111001011001",
			898 => "0010001111111100000100",
			899 => "1111111000111001011001",
			900 => "0011011011101100001000",
			901 => "0001011000111000000100",
			902 => "0000001000111001011001",
			903 => "0000000000111001011001",
			904 => "0010101000101000001000",
			905 => "0010000101101100000100",
			906 => "0000000000111001011001",
			907 => "1111111000111001011001",
			908 => "0011011110011000000100",
			909 => "0000000000111001011001",
			910 => "0000000000111001011001",
			911 => "0011000011010000000100",
			912 => "0000001000111001011001",
			913 => "0011010011010000001000",
			914 => "0000010111100100000100",
			915 => "0000000000111001011001",
			916 => "0000000000111001011001",
			917 => "1111111000111001011001",
			918 => "0000010111110000000100",
			919 => "1111111000111011100111",
			920 => "0011010110001100010000",
			921 => "0001011000111000001100",
			922 => "0010001001001100000100",
			923 => "0000000000111011100111",
			924 => "0011100101110100000100",
			925 => "0000000000111011100111",
			926 => "0000001000111011100111",
			927 => "0000000000111011100111",
			928 => "0001111011111000100000",
			929 => "0000010110010000001000",
			930 => "0001000101101100000100",
			931 => "0000001000111011100111",
			932 => "0000000000111011100111",
			933 => "0010011001001000001100",
			934 => "0000000100010100000100",
			935 => "1111111000111011100111",
			936 => "0000001110110000000100",
			937 => "0000000000111011100111",
			938 => "0000000000111011100111",
			939 => "0010111010100100001000",
			940 => "0000111100110000000100",
			941 => "0000000000111011100111",
			942 => "0000000000111011100111",
			943 => "0000000000111011100111",
			944 => "0001110011000100010000",
			945 => "0000010111100100000100",
			946 => "0000000000111011100111",
			947 => "0010101001010100000100",
			948 => "0000000000111011100111",
			949 => "0000000111111000000100",
			950 => "0000001000111011100111",
			951 => "0000000000111011100111",
			952 => "1111111000111011100111",
			953 => "0011100111100000001100",
			954 => "0011001011101100001000",
			955 => "0011000110001100000100",
			956 => "0000000000111100100001",
			957 => "0000000000111100100001",
			958 => "0000000000111100100001",
			959 => "0011100101100000001100",
			960 => "0000111000101000001000",
			961 => "0001110110011100000100",
			962 => "0000000000111100100001",
			963 => "0000000000111100100001",
			964 => "0000000000111100100001",
			965 => "0000111001010000000100",
			966 => "0000000000111100100001",
			967 => "0000000000111100100001",
			968 => "0011100101000000010000",
			969 => "0011001011101100001000",
			970 => "0001001001001000000100",
			971 => "0000000000111101100101",
			972 => "0000000000111101100101",
			973 => "0001001110011000000100",
			974 => "0000000000111101100101",
			975 => "0000000000111101100101",
			976 => "0010001001000100001000",
			977 => "0001100000100100000100",
			978 => "0000000000111101100101",
			979 => "0000000000111101100101",
			980 => "0010100100101100000100",
			981 => "0000000000111101100101",
			982 => "0001001111011000000100",
			983 => "0000000000111101100101",
			984 => "0000000000111101100101",
			985 => "0011100111100000001100",
			986 => "0011001011101100001000",
			987 => "0011000110001100000100",
			988 => "0000000000111110100001",
			989 => "0000000000111110100001",
			990 => "0000000000111110100001",
			991 => "0010111011101100000100",
			992 => "0000000000111110100001",
			993 => "0000101010101000000100",
			994 => "0000000000111110100001",
			995 => "0000111001010000000100",
			996 => "0000000000111110100001",
			997 => "0011101000110100000100",
			998 => "0000000000111110100001",
			999 => "0000000000111110100001",
			1000 => "0011100111100000000100",
			1001 => "0000000000111111011101",
			1002 => "0001011000111000001100",
			1003 => "0000000110010100000100",
			1004 => "0000000000111111011101",
			1005 => "0010111011101100000100",
			1006 => "0000000000111111011101",
			1007 => "0000000000111111011101",
			1008 => "0000111001010000001000",
			1009 => "0010101011111000000100",
			1010 => "0000000000111111011101",
			1011 => "0000000000111111011101",
			1012 => "0011010101010100000100",
			1013 => "0000000000111111011101",
			1014 => "0000000000111111011101",
			1015 => "0000100011011100000100",
			1016 => "0000000001000000011001",
			1017 => "0000111100110000010100",
			1018 => "0010010101010100001000",
			1019 => "0000010001110000000100",
			1020 => "0000000001000000011001",
			1021 => "0000000001000000011001",
			1022 => "0000001000010000001000",
			1023 => "0001111011111000000100",
			1024 => "0000000001000000011001",
			1025 => "0000000001000000011001",
			1026 => "0000000001000000011001",
			1027 => "0001011001010100000100",
			1028 => "0000000001000000011001",
			1029 => "0000000001000000011001",
			1030 => "0000001010010000100000",
			1031 => "0011100110111000001100",
			1032 => "0011001011101100001000",
			1033 => "0011011111011100000100",
			1034 => "0000000001000001100101",
			1035 => "0000000001000001100101",
			1036 => "0000000001000001100101",
			1037 => "0000000011001100001000",
			1038 => "0011101010001000000100",
			1039 => "0000000001000001100101",
			1040 => "0000000001000001100101",
			1041 => "0011110011100000001000",
			1042 => "0010010101101100000100",
			1043 => "0000000001000001100101",
			1044 => "0000000001000001100101",
			1045 => "0000000001000001100101",
			1046 => "0011110101011000000100",
			1047 => "0000000001000001100101",
			1048 => "0000000001000001100101",
			1049 => "0011000011010000100100",
			1050 => "0000111100110000010100",
			1051 => "0010010101010100001000",
			1052 => "0001101010111100000100",
			1053 => "0000000001000010111001",
			1054 => "0000000001000010111001",
			1055 => "0001111011111000001000",
			1056 => "0011010110110100000100",
			1057 => "0000000001000010111001",
			1058 => "0000000001000010111001",
			1059 => "0000000001000010111001",
			1060 => "0000001010010100001000",
			1061 => "0001011001010000000100",
			1062 => "0000001001000010111001",
			1063 => "0000000001000010111001",
			1064 => "0010011100101000000100",
			1065 => "0000000001000010111001",
			1066 => "0000000001000010111001",
			1067 => "0011110111111100000100",
			1068 => "0000000001000010111001",
			1069 => "0000000001000010111001",
			1070 => "0011100111100000001100",
			1071 => "0011001011101100001000",
			1072 => "0011000110001100000100",
			1073 => "0000000001000100001101",
			1074 => "0000000001000100001101",
			1075 => "0000000001000100001101",
			1076 => "0011110011100000011000",
			1077 => "0011011110011000001000",
			1078 => "0001110100101100000100",
			1079 => "0000000001000100001101",
			1080 => "0000000001000100001101",
			1081 => "0010100100101100001000",
			1082 => "0011100110000100000100",
			1083 => "0000000001000100001101",
			1084 => "0000000001000100001101",
			1085 => "0001000011000000000100",
			1086 => "0000000001000100001101",
			1087 => "0000000001000100001101",
			1088 => "0011110101011000000100",
			1089 => "0000000001000100001101",
			1090 => "0000000001000100001101",
			1091 => "0011100111100000000100",
			1092 => "1111111001000101000001",
			1093 => "0001110011000100010100",
			1094 => "0011100101100000010000",
			1095 => "0001011001010000001100",
			1096 => "0001111011111000001000",
			1097 => "0010010101011100000100",
			1098 => "0000001001000101000001",
			1099 => "0000000001000101000001",
			1100 => "0000010001000101000001",
			1101 => "1111111001000101000001",
			1102 => "0000000001000101000001",
			1103 => "1111111001000101000001",
			1104 => "0011110000100100010000",
			1105 => "0001001110011000001100",
			1106 => "0000010110010000001000",
			1107 => "0000010111110000000100",
			1108 => "0000000001000110001101",
			1109 => "0000000001000110001101",
			1110 => "0000000001000110001101",
			1111 => "1111111001000110001101",
			1112 => "0010010101010100000100",
			1113 => "0000000001000110001101",
			1114 => "0000001010010000010000",
			1115 => "0001110011000100001100",
			1116 => "0001111100101100001000",
			1117 => "0001011000000000000100",
			1118 => "0000000001000110001101",
			1119 => "0000000001000110001101",
			1120 => "0000000001000110001101",
			1121 => "0000000001000110001101",
			1122 => "1111111001000110001101",
			1123 => "0010111011101100010000",
			1124 => "0000000010100100000100",
			1125 => "0000000001000111101001",
			1126 => "0000010001110000000100",
			1127 => "0000000001000111101001",
			1128 => "0011100110111000000100",
			1129 => "0000000001000111101001",
			1130 => "0000000001000111101001",
			1131 => "0000101010101000001100",
			1132 => "0010000101101100000100",
			1133 => "0000000001000111101001",
			1134 => "0011110101111100000100",
			1135 => "0000000001000111101001",
			1136 => "0000000001000111101001",
			1137 => "0001000111011100000100",
			1138 => "0000000001000111101001",
			1139 => "0000010110001100001000",
			1140 => "0010101011000000000100",
			1141 => "0000000001000111101001",
			1142 => "0000000001000111101001",
			1143 => "0010001111011000000100",
			1144 => "0000000001000111101001",
			1145 => "0000000001000111101001",
			1146 => "0011100110111000000100",
			1147 => "1111111001001000100101",
			1148 => "0001011001010000011000",
			1149 => "0011011010100100010000",
			1150 => "0011101000110100001100",
			1151 => "0000001010000000000100",
			1152 => "0000000001001000100101",
			1153 => "0000100000000000000100",
			1154 => "0000011001001000100101",
			1155 => "0000010001001000100101",
			1156 => "0000001001001000100101",
			1157 => "0010101000101000000100",
			1158 => "1111111001001000100101",
			1159 => "0000001001001000100101",
			1160 => "1111111001001000100101",
			1161 => "0000111100110000100000",
			1162 => "0010111011101100001100",
			1163 => "0000000110010100000100",
			1164 => "0000000001001010000001",
			1165 => "0011100110111000000100",
			1166 => "0000000001001010000001",
			1167 => "0000000001001010000001",
			1168 => "0000001001110100010000",
			1169 => "0001111011111000000100",
			1170 => "0000000001001010000001",
			1171 => "0001000101010100000100",
			1172 => "0000000001001010000001",
			1173 => "0001111011000000000100",
			1174 => "0000000001001010000001",
			1175 => "0000000001001010000001",
			1176 => "1111111001001010000001",
			1177 => "0001011001010000001100",
			1178 => "0000001010010100001000",
			1179 => "0011111100111100000100",
			1180 => "0000000001001010000001",
			1181 => "0000000001001010000001",
			1182 => "0000000001001010000001",
			1183 => "0000000001001010000001",
			1184 => "0011100110110000000100",
			1185 => "1111111001001011010101",
			1186 => "0011011010100100010100",
			1187 => "0000111100110000001100",
			1188 => "0010011100101000001000",
			1189 => "0001010011001000000100",
			1190 => "0000000001001011010101",
			1191 => "0000000001001011010101",
			1192 => "1111111001001011010101",
			1193 => "0000001010010100000100",
			1194 => "0000001001001011010101",
			1195 => "1111111001001011010101",
			1196 => "0011100100000100001000",
			1197 => "0000101010101000000100",
			1198 => "0000000001001011010101",
			1199 => "1111111001001011010101",
			1200 => "0000111001010000000100",
			1201 => "1111111001001011010101",
			1202 => "0000001010111000000100",
			1203 => "0000001001001011010101",
			1204 => "0000000001001011010101",
			1205 => "0001000101101100101000",
			1206 => "0001111011111000011100",
			1207 => "0001111000101000010000",
			1208 => "0000111111011000000100",
			1209 => "1111111001001100111001",
			1210 => "0010010101011100001000",
			1211 => "0011100110110000000100",
			1212 => "0000000001001100111001",
			1213 => "0000001001001100111001",
			1214 => "0000000001001100111001",
			1215 => "0001011000000000001000",
			1216 => "0000001100001000000100",
			1217 => "1111111001001100111001",
			1218 => "0000000001001100111001",
			1219 => "0000000001001100111001",
			1220 => "0001110011000100001000",
			1221 => "0010101001010100000100",
			1222 => "0000000001001100111001",
			1223 => "0000001001001100111001",
			1224 => "1111111001001100111001",
			1225 => "0011100101000000000100",
			1226 => "1111111001001100111001",
			1227 => "0001010100101100000100",
			1228 => "0000000001001100111001",
			1229 => "0000000001001100111001",
			1230 => "0011110000001000000100",
			1231 => "1111111001001110000101",
			1232 => "0000000111111000011000",
			1233 => "0001011111011000000100",
			1234 => "0000000001001110000101",
			1235 => "0011011010100100001000",
			1236 => "0000111100110000000100",
			1237 => "0000001001001110000101",
			1238 => "0000001001001110000101",
			1239 => "0000100110101000001000",
			1240 => "0010100100101100000100",
			1241 => "1111111001001110000101",
			1242 => "0000001001001110000101",
			1243 => "0000001001001110000101",
			1244 => "0001010101111000000100",
			1245 => "0000001001001110000101",
			1246 => "0001011000000000000100",
			1247 => "0000000001001110000101",
			1248 => "1111111001001110000101",
			1249 => "0000111100110000101000",
			1250 => "0010011100101000011100",
			1251 => "0011011011101100010100",
			1252 => "0011001011101100001000",
			1253 => "0000000110010100000100",
			1254 => "0000000001001111110001",
			1255 => "0000000001001111110001",
			1256 => "0000000011001100001000",
			1257 => "0001011000000100000100",
			1258 => "0000000001001111110001",
			1259 => "0000000001001111110001",
			1260 => "0000000001001111110001",
			1261 => "0000110011001000000100",
			1262 => "0000000001001111110001",
			1263 => "0000000001001111110001",
			1264 => "0011011011101100001000",
			1265 => "0001000110000000000100",
			1266 => "0000000001001111110001",
			1267 => "0000000001001111110001",
			1268 => "0000000001001111110001",
			1269 => "0000100011011100000100",
			1270 => "0000000001001111110001",
			1271 => "0001011001010000001000",
			1272 => "0000001010010100000100",
			1273 => "0000001001001111110001",
			1274 => "0000000001001111110001",
			1275 => "0000000001001111110001",
			1276 => "0001100000010000000100",
			1277 => "1111111001010000110101",
			1278 => "0001011001010000011100",
			1279 => "0000111100110000010100",
			1280 => "0010111011101100001000",
			1281 => "0001100000001000000100",
			1282 => "0000000001010000110101",
			1283 => "0000001001010000110101",
			1284 => "0011111000100100001000",
			1285 => "0010000101101100000100",
			1286 => "1111111001010000110101",
			1287 => "0000001001010000110101",
			1288 => "1111111001010000110101",
			1289 => "0011110100110100000100",
			1290 => "0000001001010000110101",
			1291 => "0000001001010000110101",
			1292 => "1111111001010000110101",
			1293 => "0010111011101100010100",
			1294 => "0000000010100100000100",
			1295 => "0000000001010010110001",
			1296 => "0001011000000000001000",
			1297 => "0000010111110000000100",
			1298 => "0000000001010010110001",
			1299 => "0000001001010010110001",
			1300 => "0011001110011000000100",
			1301 => "0000000001010010110001",
			1302 => "0000000001010010110001",
			1303 => "0000101010101000010000",
			1304 => "0010000101101100001000",
			1305 => "0000001010000000000100",
			1306 => "0000000001010010110001",
			1307 => "0000000001010010110001",
			1308 => "0011110000001000000100",
			1309 => "0000000001010010110001",
			1310 => "0000001001010010110001",
			1311 => "0000111001010000010000",
			1312 => "0001000110000000001000",
			1313 => "0000010110010000000100",
			1314 => "0000000001010010110001",
			1315 => "1111111001010010110001",
			1316 => "0001100000001000000100",
			1317 => "0000000001010010110001",
			1318 => "0000000001010010110001",
			1319 => "0011101000110100000100",
			1320 => "0000000001010010110001",
			1321 => "0000001101011000000100",
			1322 => "0000000001010010110001",
			1323 => "0000000001010010110001",
			1324 => "0001011000000100011000",
			1325 => "0001110100101100010000",
			1326 => "0001111000101000001100",
			1327 => "0010111011101100001000",
			1328 => "0001100000010000000100",
			1329 => "0000000001010100101101",
			1330 => "0000000001010100101101",
			1331 => "0000000001010100101101",
			1332 => "0000000001010100101101",
			1333 => "0000110011100100000100",
			1334 => "0000000001010100101101",
			1335 => "0000000001010100101101",
			1336 => "0011110000100100001100",
			1337 => "0000010110010000001000",
			1338 => "0000010111110000000100",
			1339 => "0000000001010100101101",
			1340 => "0000000001010100101101",
			1341 => "0000000001010100101101",
			1342 => "0011110011100000010100",
			1343 => "0011011010100100001000",
			1344 => "0000001110110000000100",
			1345 => "0000000001010100101101",
			1346 => "0000000001010100101101",
			1347 => "0010100100101100000100",
			1348 => "0000000001010100101101",
			1349 => "0010101011111000000100",
			1350 => "0000000001010100101101",
			1351 => "0000000001010100101101",
			1352 => "0010101011111000000100",
			1353 => "0000000001010100101101",
			1354 => "0000000001010100101101",
			1355 => "0011110000100100010000",
			1356 => "0001001110011000001100",
			1357 => "0000010110010000001000",
			1358 => "0000010111110000000100",
			1359 => "0000000001010110001001",
			1360 => "0000000001010110001001",
			1361 => "0000000001010110001001",
			1362 => "1111111001010110001001",
			1363 => "0010010101010100000100",
			1364 => "0000000001010110001001",
			1365 => "0000001010010000011000",
			1366 => "0000111100110000001100",
			1367 => "0001011000000100000100",
			1368 => "1111111001010110001001",
			1369 => "0011011110011000000100",
			1370 => "0000000001010110001001",
			1371 => "0000000001010110001001",
			1372 => "0001111100101100000100",
			1373 => "0000000001010110001001",
			1374 => "0001000101111000000100",
			1375 => "0000001001010110001001",
			1376 => "0000000001010110001001",
			1377 => "1111111001010110001001",
			1378 => "0011100110110000000100",
			1379 => "1111111001010111101101",
			1380 => "0011011010100100011000",
			1381 => "0000001010010100001100",
			1382 => "0000000010100100001000",
			1383 => "0010011001001000000100",
			1384 => "0000000001010111101101",
			1385 => "0000001001010111101101",
			1386 => "0000001001010111101101",
			1387 => "0010111011101100000100",
			1388 => "0000000001010111101101",
			1389 => "0000010110010000000100",
			1390 => "0000000001010111101101",
			1391 => "1111111001010111101101",
			1392 => "0011100100000100001100",
			1393 => "0000101010101000000100",
			1394 => "0000000001010111101101",
			1395 => "0010101000101000000100",
			1396 => "1111111001010111101101",
			1397 => "1111111001010111101101",
			1398 => "0000111001010000000100",
			1399 => "1111111001010111101101",
			1400 => "0001001100000000000100",
			1401 => "0000001001010111101101",
			1402 => "0000000001010111101101",
			1403 => "0011100001100000101000",
			1404 => "0010010101010100001100",
			1405 => "0001001110011000001000",
			1406 => "0001111000000000000100",
			1407 => "0000000001011001110001",
			1408 => "0000000001011001110001",
			1409 => "0000000001011001110001",
			1410 => "0011010110110100001100",
			1411 => "0000111101001000001000",
			1412 => "0000111000000000000100",
			1413 => "0000000001011001110001",
			1414 => "0000000001011001110001",
			1415 => "0000000001011001110001",
			1416 => "0000111001010000001000",
			1417 => "0011111000100100000100",
			1418 => "0000000001011001110001",
			1419 => "0000000001011001110001",
			1420 => "0000111000101000000100",
			1421 => "0000000001011001110001",
			1422 => "0000000001011001110001",
			1423 => "0011110011100000010100",
			1424 => "0011011010100100000100",
			1425 => "0000000001011001110001",
			1426 => "0011110100110100000100",
			1427 => "0000000001011001110001",
			1428 => "0011110000011100001000",
			1429 => "0010101001011000000100",
			1430 => "0000000001011001110001",
			1431 => "0000000001011001110001",
			1432 => "0000000001011001110001",
			1433 => "0000111001010000000100",
			1434 => "0000000001011001110001",
			1435 => "0000000001011001110001",
			1436 => "0001100000010000000100",
			1437 => "1111111001011010111101",
			1438 => "0001011001010000100000",
			1439 => "0000001010010100001100",
			1440 => "0000100111011000000100",
			1441 => "0000000001011010111101",
			1442 => "0011101100000100000100",
			1443 => "0000010001011010111101",
			1444 => "0000001001011010111101",
			1445 => "0001001010100100000100",
			1446 => "0000001001011010111101",
			1447 => "0001110001010000001000",
			1448 => "0010111110011000000100",
			1449 => "0000001001011010111101",
			1450 => "1111111001011010111101",
			1451 => "0001011100110000000100",
			1452 => "1111111001011010111101",
			1453 => "1111111001011010111101",
			1454 => "1111111001011010111101",
			1455 => "0001111011111000100000",
			1456 => "0011010110001100001100",
			1457 => "0000010111110000000100",
			1458 => "0000000001011100111001",
			1459 => "0001111100010000000100",
			1460 => "0000000001011100111001",
			1461 => "0000000001011100111001",
			1462 => "0010010101010100000100",
			1463 => "0000000001011100111001",
			1464 => "0001001100101000000100",
			1465 => "0000000001011100111001",
			1466 => "0001000101101100000100",
			1467 => "0000000001011100111001",
			1468 => "0001011000000100000100",
			1469 => "0000000001011100111001",
			1470 => "0000000001011100111001",
			1471 => "0000000111111000011100",
			1472 => "0001111011000000001100",
			1473 => "0001011001010000001000",
			1474 => "0010101001010100000100",
			1475 => "0000000001011100111001",
			1476 => "0000000001011100111001",
			1477 => "0000000001011100111001",
			1478 => "0000111001010000000100",
			1479 => "0000000001011100111001",
			1480 => "0010001001000100000100",
			1481 => "0000000001011100111001",
			1482 => "0001001000000100000100",
			1483 => "0000000001011100111001",
			1484 => "0000000001011100111001",
			1485 => "0000000001011100111001",
			1486 => "0000100011011100000100",
			1487 => "1111111001011110011101",
			1488 => "0000000111111000011100",
			1489 => "0011011010100100010000",
			1490 => "0000110011001000000100",
			1491 => "1111111001011110011101",
			1492 => "0001011001010000001000",
			1493 => "0001100000010000000100",
			1494 => "0000000001011110011101",
			1495 => "0000001001011110011101",
			1496 => "0000000001011110011101",
			1497 => "0010100100101100000100",
			1498 => "1111111001011110011101",
			1499 => "0001001111011000000100",
			1500 => "0000001001011110011101",
			1501 => "0000000001011110011101",
			1502 => "0001011111011000000100",
			1503 => "0000000001011110011101",
			1504 => "0011011110011000001000",
			1505 => "0000110011100100000100",
			1506 => "0000000001011110011101",
			1507 => "1111111001011110011101",
			1508 => "0001011100110000000100",
			1509 => "0000000001011110011101",
			1510 => "1111111001011110011101",
			1511 => "0011110000001000000100",
			1512 => "1111111001011111111001",
			1513 => "0000000111111000010100",
			1514 => "0001011111011000000100",
			1515 => "1111111001011111111001",
			1516 => "0000111000101000001100",
			1517 => "0001100100100000000100",
			1518 => "0000011001011111111001",
			1519 => "0001111001011000000100",
			1520 => "0000001001011111111001",
			1521 => "1111111001011111111001",
			1522 => "0000000001011111111001",
			1523 => "0001010101111000000100",
			1524 => "0000001001011111111001",
			1525 => "0001110001010000001100",
			1526 => "0010001111111100000100",
			1527 => "1111111001011111111001",
			1528 => "0010111110011000000100",
			1529 => "0000001001011111111001",
			1530 => "1111111001011111111001",
			1531 => "0011101000010100000100",
			1532 => "1111111001011111111001",
			1533 => "0000000001011111111001",
			1534 => "0000111100110000110000",
			1535 => "0010010101010100001100",
			1536 => "0000010001110000000100",
			1537 => "0000000001100010010101",
			1538 => "0001100001111000000100",
			1539 => "0000000001100010010101",
			1540 => "0000001001100010010101",
			1541 => "0000101011100000010000",
			1542 => "0010011100101000001100",
			1543 => "0001000101011100001000",
			1544 => "0001110110101100000100",
			1545 => "0000000001100010010101",
			1546 => "0000000001100010010101",
			1547 => "0000000001100010010101",
			1548 => "0000000001100010010101",
			1549 => "0010111011101100001000",
			1550 => "0011010110001100000100",
			1551 => "0000000001100010010101",
			1552 => "0000000001100010010101",
			1553 => "0010001111001000000100",
			1554 => "1111111001100010010101",
			1555 => "0000000100010100000100",
			1556 => "0000000001100010010101",
			1557 => "0000000001100010010101",
			1558 => "0000111000101000010100",
			1559 => "0000001010010100001000",
			1560 => "0011111100111100000100",
			1561 => "0000000001100010010101",
			1562 => "0000001001100010010101",
			1563 => "0000010011110000001000",
			1564 => "0011110100111100000100",
			1565 => "0000000001100010010101",
			1566 => "0000000001100010010101",
			1567 => "0000000001100010010101",
			1568 => "0011100100000100000100",
			1569 => "1111111001100010010101",
			1570 => "0000001101011000000100",
			1571 => "0000000001100010010101",
			1572 => "0000000001100010010101",
			1573 => "0000111100110000110000",
			1574 => "0010010101010100001100",
			1575 => "0000010001110000000100",
			1576 => "0000000001100100110001",
			1577 => "0001100001111000000100",
			1578 => "0000000001100100110001",
			1579 => "0000001001100100110001",
			1580 => "0001011111011000001100",
			1581 => "0000010110010000001000",
			1582 => "0000010111110000000100",
			1583 => "0000000001100100110001",
			1584 => "0000000001100100110001",
			1585 => "1111111001100100110001",
			1586 => "0000001111101100010000",
			1587 => "0011011110011000001100",
			1588 => "0000110011100100000100",
			1589 => "0000000001100100110001",
			1590 => "0001001001000100000100",
			1591 => "0000001001100100110001",
			1592 => "0000000001100100110001",
			1593 => "0000000001100100110001",
			1594 => "0011001110011000000100",
			1595 => "0000000001100100110001",
			1596 => "1111111001100100110001",
			1597 => "0000111000101000010100",
			1598 => "0000001010010100001000",
			1599 => "0011111100111100000100",
			1600 => "0000000001100100110001",
			1601 => "0000001001100100110001",
			1602 => "0000010011110000001000",
			1603 => "0011110100111100000100",
			1604 => "0000000001100100110001",
			1605 => "0000000001100100110001",
			1606 => "0000000001100100110001",
			1607 => "0011100100000100000100",
			1608 => "1111111001100100110001",
			1609 => "0000001101011000000100",
			1610 => "0000000001100100110001",
			1611 => "0000000001100100110001",
			1612 => "0000010111100100001100",
			1613 => "0001010101111000001000",
			1614 => "0000111111011000000100",
			1615 => "0000000001100110111101",
			1616 => "0000000001100110111101",
			1617 => "0000000001100110111101",
			1618 => "0000011000011000011000",
			1619 => "0001001010100100001000",
			1620 => "0001001101000000000100",
			1621 => "0000000001100110111101",
			1622 => "0000000001100110111101",
			1623 => "0001001001001000000100",
			1624 => "0000001001100110111101",
			1625 => "0001110100101100000100",
			1626 => "0000000001100110111101",
			1627 => "0010001111001000000100",
			1628 => "0000000001100110111101",
			1629 => "0000000001100110111101",
			1630 => "0001000011010000001100",
			1631 => "0011011011101100000100",
			1632 => "0000000001100110111101",
			1633 => "0010111010100100000100",
			1634 => "0000000001100110111101",
			1635 => "0000000001100110111101",
			1636 => "0001011100010000001100",
			1637 => "0001011000000100001000",
			1638 => "0001011111011000000100",
			1639 => "0000000001100110111101",
			1640 => "0000000001100110111101",
			1641 => "0000000001100110111101",
			1642 => "0000000110010100001000",
			1643 => "0011100100010000000100",
			1644 => "0000000001100110111101",
			1645 => "0000000001100110111101",
			1646 => "0000000001100110111101",
			1647 => "0011100110110000000100",
			1648 => "1111111001101000000001",
			1649 => "0001110011000100011100",
			1650 => "0000110011001000000100",
			1651 => "0000000001101000000001",
			1652 => "0000010111110000000100",
			1653 => "1111111001101000000001",
			1654 => "0001111000101000000100",
			1655 => "0000001001101000000001",
			1656 => "0000000111111000001000",
			1657 => "0000000110101000000100",
			1658 => "0000000001101000000001",
			1659 => "0000001001101000000001",
			1660 => "0000010011110000000100",
			1661 => "0000000001101000000001",
			1662 => "1111111001101000000001",
			1663 => "1111111001101000000001",
			1664 => "0011110000001000000100",
			1665 => "1111111001101001010101",
			1666 => "0010010101010100000100",
			1667 => "0000001001101001010101",
			1668 => "0000110011100100001000",
			1669 => "0011011011101100000100",
			1670 => "0000000001101001010101",
			1671 => "1111111001101001010101",
			1672 => "0000000111111000010000",
			1673 => "0001100000001100000100",
			1674 => "0000001001101001010101",
			1675 => "0011001010100100000100",
			1676 => "0000000001101001010101",
			1677 => "0000000110010100000100",
			1678 => "0000001001101001010101",
			1679 => "0000000001101001010101",
			1680 => "0000010011110000001000",
			1681 => "0010111110011000000100",
			1682 => "0000000001101001010101",
			1683 => "1111111001101001010101",
			1684 => "1111111001101001010101",
			1685 => "0000010111100100010100",
			1686 => "0001001110011000001000",
			1687 => "0000101001110100000100",
			1688 => "0000000001101011101001",
			1689 => "0000000001101011101001",
			1690 => "0001010101111000001000",
			1691 => "0001011101101000000100",
			1692 => "0000000001101011101001",
			1693 => "0000000001101011101001",
			1694 => "0000000001101011101001",
			1695 => "0011010110001100001000",
			1696 => "0001111100110000000100",
			1697 => "0000000001101011101001",
			1698 => "0000000001101011101001",
			1699 => "0001111011111000011000",
			1700 => "0010011001001000001100",
			1701 => "0001111000101000001000",
			1702 => "0011001011101100000100",
			1703 => "0000000001101011101001",
			1704 => "0000000001101011101001",
			1705 => "0000000001101011101001",
			1706 => "0001000101101100001000",
			1707 => "0001110001010000000100",
			1708 => "0000000001101011101001",
			1709 => "0000000001101011101001",
			1710 => "0000000001101011101001",
			1711 => "0001110011000100010100",
			1712 => "0011010011010000001000",
			1713 => "0000000110111100000100",
			1714 => "0000001001101011101001",
			1715 => "0000000001101011101001",
			1716 => "0000010110001100000100",
			1717 => "0000000001101011101001",
			1718 => "0001011000101000000100",
			1719 => "0000000001101011101001",
			1720 => "0000000001101011101001",
			1721 => "0000000001101011101001",
			1722 => "0011100110110000000100",
			1723 => "1111111001101101000101",
			1724 => "0011010110001100000100",
			1725 => "0000001001101101000101",
			1726 => "0000001010010000100000",
			1727 => "0011010011010000010100",
			1728 => "0001110100101100001000",
			1729 => "0000001101111000000100",
			1730 => "0000000001101101000101",
			1731 => "0000001001101101000101",
			1732 => "0000010111100100000100",
			1733 => "0000000001101101000101",
			1734 => "0000001000010000000100",
			1735 => "0000001001101101000101",
			1736 => "0000000001101101000101",
			1737 => "0010101111101000001000",
			1738 => "0011110100111100000100",
			1739 => "1111111001101101000101",
			1740 => "0000000001101101000101",
			1741 => "1111111001101101000101",
			1742 => "0001100010101000000100",
			1743 => "1111111001101101000101",
			1744 => "0000000001101101000101",
			1745 => "0011110000001000000100",
			1746 => "1111111001101110101001",
			1747 => "0000010111110000001000",
			1748 => "0000110011001000000100",
			1749 => "0000000001101110101001",
			1750 => "1111111001101110101001",
			1751 => "0000110011001000001000",
			1752 => "0001111001010000000100",
			1753 => "0000000001101110101001",
			1754 => "1111111001101110101001",
			1755 => "0011011010100100010000",
			1756 => "0010100100101100001100",
			1757 => "0001001001000100001000",
			1758 => "0011110111001100000100",
			1759 => "0000001001101110101001",
			1760 => "0000000001101110101001",
			1761 => "1111111001101110101001",
			1762 => "0000000001101110101001",
			1763 => "0011110111101100001100",
			1764 => "0010100100101100000100",
			1765 => "1111111001101110101001",
			1766 => "0001000011000000000100",
			1767 => "0000001001101110101001",
			1768 => "0000000001101110101001",
			1769 => "0000001001101110101001",
			1770 => "0000010111110000001000",
			1771 => "0001111011111000000100",
			1772 => "0000000001110000101101",
			1773 => "0000000001110000101101",
			1774 => "0000100111110100010000",
			1775 => "0001010011001000001000",
			1776 => "0001010101111000000100",
			1777 => "0000000001110000101101",
			1778 => "0000000001110000101101",
			1779 => "0000010110010000000100",
			1780 => "0000000001110000101101",
			1781 => "0000000001110000101101",
			1782 => "0011110011100000100100",
			1783 => "0011011010100100010000",
			1784 => "0000001110110000001100",
			1785 => "0001011001010000001000",
			1786 => "0000110011001000000100",
			1787 => "0000000001110000101101",
			1788 => "0000001001110000101101",
			1789 => "0000000001110000101101",
			1790 => "0000000001110000101101",
			1791 => "0000101010101000001000",
			1792 => "0000000011111000000100",
			1793 => "0000000001110000101101",
			1794 => "0000000001110000101101",
			1795 => "0011110111001100001000",
			1796 => "0000010110001100000100",
			1797 => "0000000001110000101101",
			1798 => "0000000001110000101101",
			1799 => "0000000001110000101101",
			1800 => "0000111001010000000100",
			1801 => "0000000001110000101101",
			1802 => "0000000001110000101101",
			1803 => "0000010111100100011000",
			1804 => "0001001110011000001100",
			1805 => "0010001001000100001000",
			1806 => "0001111100010000000100",
			1807 => "0000000001110011101001",
			1808 => "0000000001110011101001",
			1809 => "0000000001110011101001",
			1810 => "0001010101111000001000",
			1811 => "0001010011000000000100",
			1812 => "0000000001110011101001",
			1813 => "0000000001110011101001",
			1814 => "0000000001110011101001",
			1815 => "0000011000011000011000",
			1816 => "0001001010100100001000",
			1817 => "0001001101000000000100",
			1818 => "0000000001110011101001",
			1819 => "0000000001110011101001",
			1820 => "0001001001001000000100",
			1821 => "0000000001110011101001",
			1822 => "0001110100101100000100",
			1823 => "0000000001110011101001",
			1824 => "0010001010000100000100",
			1825 => "0000000001110011101001",
			1826 => "0000000001110011101001",
			1827 => "0001111100101100011100",
			1828 => "0001011100010000010100",
			1829 => "0001001110011000001000",
			1830 => "0001110110101100000100",
			1831 => "0000000001110011101001",
			1832 => "0000000001110011101001",
			1833 => "0001011000000100001000",
			1834 => "0001011111011000000100",
			1835 => "0000000001110011101001",
			1836 => "0000000001110011101001",
			1837 => "0000000001110011101001",
			1838 => "0001000110000000000100",
			1839 => "0000000001110011101001",
			1840 => "0000000001110011101001",
			1841 => "0001110110011100010000",
			1842 => "0011010101010100000100",
			1843 => "0000000001110011101001",
			1844 => "0000111001010000000100",
			1845 => "0000000001110011101001",
			1846 => "0000111011111000000100",
			1847 => "0000000001110011101001",
			1848 => "0000000001110011101001",
			1849 => "0000000001110011101001",
			1850 => "0010010101010100001100",
			1851 => "0000010001110000000100",
			1852 => "0000000001110101100111",
			1853 => "0011111000001000000100",
			1854 => "0000000001110101100111",
			1855 => "0000001001110101100111",
			1856 => "0000101101110000110000",
			1857 => "0011010110001100001000",
			1858 => "0000010111100100000100",
			1859 => "0000000001110101100111",
			1860 => "0000001001110101100111",
			1861 => "0001110100101100010100",
			1862 => "0000001101111000001100",
			1863 => "0000111001010000000100",
			1864 => "1111111001110101100111",
			1865 => "0010111010100100000100",
			1866 => "0000000001110101100111",
			1867 => "0000000001110101100111",
			1868 => "0011101111010100000100",
			1869 => "0000000001110101100111",
			1870 => "0000000001110101100111",
			1871 => "0011011110011000000100",
			1872 => "0000000001110101100111",
			1873 => "0010100100101100001000",
			1874 => "0000100110101000000100",
			1875 => "1111111001110101100111",
			1876 => "0000001001110101100111",
			1877 => "0001000101111000000100",
			1878 => "0000001001110101100111",
			1879 => "0000000001110101100111",
			1880 => "1111111001110101100111",
			1881 => "0001100101111100010000",
			1882 => "0011100110111000000100",
			1883 => "1100000001110110100001",
			1884 => "0010011001001000000100",
			1885 => "1110001001110110100001",
			1886 => "0010011001000100000100",
			1887 => "1100100001110110100001",
			1888 => "1100000001110110100001",
			1889 => "0010010101101100001000",
			1890 => "0000111100110000000100",
			1891 => "1110100001110110100001",
			1892 => "1111111001110110100001",
			1893 => "0000101101111000000100",
			1894 => "1100010001110110100001",
			1895 => "1100000001110110100001",
			1896 => "0011100111100000000100",
			1897 => "1111111001110111001101",
			1898 => "0011000111011100010000",
			1899 => "0011100101100000001100",
			1900 => "0001111011111000001000",
			1901 => "0011111110011100000100",
			1902 => "0000000001110111001101",
			1903 => "0000001001110111001101",
			1904 => "0000001001110111001101",
			1905 => "0000000001110111001101",
			1906 => "1111111001110111001101",
			1907 => "0011100111100000001100",
			1908 => "0011011101000000001000",
			1909 => "0011011111011100000100",
			1910 => "0000000001111000010001",
			1911 => "0000000001111000010001",
			1912 => "0000000001111000010001",
			1913 => "0011101100000100001000",
			1914 => "0001011100110000000100",
			1915 => "0000000001111000010001",
			1916 => "0000000001111000010001",
			1917 => "0001111100101100000100",
			1918 => "0000000001111000010001",
			1919 => "0000111100110000000100",
			1920 => "0000000001111000010001",
			1921 => "0001011000101000000100",
			1922 => "0000000001111000010001",
			1923 => "0000000001111000010001",
			1924 => "0011100111100000001100",
			1925 => "0011011101000000001000",
			1926 => "0000111100010000000100",
			1927 => "0000000001111001011101",
			1928 => "0000000001111001011101",
			1929 => "0000000001111001011101",
			1930 => "0001111011111000001100",
			1931 => "0001111000101000000100",
			1932 => "0000000001111001011101",
			1933 => "0001011000000000000100",
			1934 => "0000000001111001011101",
			1935 => "0000000001111001011101",
			1936 => "0011000011010000000100",
			1937 => "0000000001111001011101",
			1938 => "0001000110000000000100",
			1939 => "0000000001111001011101",
			1940 => "0001000101111000000100",
			1941 => "0000000001111001011101",
			1942 => "0000000001111001011101",
			1943 => "0000010111100100010100",
			1944 => "0001001110011000001100",
			1945 => "0010001001000100001000",
			1946 => "0001111100010000000100",
			1947 => "0000000001111010110001",
			1948 => "0000000001111010110001",
			1949 => "0000000001111010110001",
			1950 => "0001011101101000000100",
			1951 => "0000000001111010110001",
			1952 => "0000000001111010110001",
			1953 => "0000110011100100001000",
			1954 => "0011001011101100000100",
			1955 => "0000000001111010110001",
			1956 => "0000000001111010110001",
			1957 => "0001011001010000001100",
			1958 => "0011100101100000001000",
			1959 => "0011110000001000000100",
			1960 => "0000000001111010110001",
			1961 => "0000000001111010110001",
			1962 => "0000000001111010110001",
			1963 => "0000000001111010110001",
			1964 => "0001000111011100010000",
			1965 => "0000100010101100001000",
			1966 => "0000111100110000000100",
			1967 => "0000000001111100001101",
			1968 => "0000000001111100001101",
			1969 => "0000111111011000000100",
			1970 => "0000000001111100001101",
			1971 => "0000000001111100001101",
			1972 => "0000101010101000010000",
			1973 => "0001111111101000000100",
			1974 => "0000000001111100001101",
			1975 => "0010101001010100000100",
			1976 => "0000000001111100001101",
			1977 => "0001000011000000000100",
			1978 => "0000000001111100001101",
			1979 => "0000000001111100001101",
			1980 => "0010111011101100001000",
			1981 => "0010101000101000000100",
			1982 => "0000000001111100001101",
			1983 => "0000000001111100001101",
			1984 => "0001011000000100000100",
			1985 => "0000000001111100001101",
			1986 => "0000000001111100001101",
			1987 => "0000000111111000011000",
			1988 => "0011110000001000000100",
			1989 => "0000000001111101100001",
			1990 => "0001011111011000000100",
			1991 => "0000000001111101100001",
			1992 => "0011011010100100001000",
			1993 => "0011110000100100000100",
			1994 => "0000000001111101100001",
			1995 => "0000000001111101100001",
			1996 => "0010100100101100000100",
			1997 => "0000000001111101100001",
			1998 => "0000000001111101100001",
			1999 => "0001110001010000001100",
			2000 => "0010111110011000001000",
			2001 => "0001100111010000000100",
			2002 => "0000000001111101100001",
			2003 => "0000000001111101100001",
			2004 => "0000000001111101100001",
			2005 => "0011101000010100000100",
			2006 => "0000000001111101100001",
			2007 => "0000000001111101100001",
			2008 => "0011110000100100010100",
			2009 => "0001011000000100001000",
			2010 => "0000111000000000000100",
			2011 => "0000000001111110111101",
			2012 => "0000000001111110111101",
			2013 => "0000111001010000000100",
			2014 => "0000000001111110111101",
			2015 => "0000111111101000000100",
			2016 => "0000000001111110111101",
			2017 => "0000000001111110111101",
			2018 => "0011110011100000010100",
			2019 => "0000101101110000010000",
			2020 => "0011011010100100001000",
			2021 => "0001011000000100000100",
			2022 => "0000000001111110111101",
			2023 => "0000000001111110111101",
			2024 => "0000111001010000000100",
			2025 => "0000000001111110111101",
			2026 => "0000000001111110111101",
			2027 => "0000000001111110111101",
			2028 => "0000111001010000000100",
			2029 => "0000000001111110111101",
			2030 => "0000000001111110111101",
			2031 => "0011100110111000000100",
			2032 => "1111111001111111111001",
			2033 => "0001110011000100011000",
			2034 => "0001111011111000001100",
			2035 => "0010111011101100000100",
			2036 => "0000000001111111111001",
			2037 => "0001011000000000000100",
			2038 => "1111111001111111111001",
			2039 => "0000000001111111111001",
			2040 => "0011011110011000000100",
			2041 => "0000001001111111111001",
			2042 => "0010100100101100000100",
			2043 => "0000000001111111111001",
			2044 => "0000001001111111111001",
			2045 => "1111111001111111111001",
			2046 => "0011100111100000001100",
			2047 => "0011011101000000001000",
			2048 => "0000010110010000000100",
			2049 => "0000000010000001001101",
			2050 => "0000000010000001001101",
			2051 => "1111111010000001001101",
			2052 => "0011110011100000011000",
			2053 => "0010000101101100001000",
			2054 => "0011111000100100000100",
			2055 => "0000000010000001001101",
			2056 => "0000001010000001001101",
			2057 => "0011010011010000000100",
			2058 => "0000001010000001001101",
			2059 => "0000010110001100000100",
			2060 => "1111111010000001001101",
			2061 => "0000011110011000000100",
			2062 => "0000000010000001001101",
			2063 => "0000000010000001001101",
			2064 => "0001011000000100000100",
			2065 => "0000000010000001001101",
			2066 => "1111111010000001001101",
			2067 => "0011110011111100100100",
			2068 => "0001110100101100010100",
			2069 => "0011011110011000001100",
			2070 => "0011010110110100001000",
			2071 => "0011011111011100000100",
			2072 => "0000000010000010110001",
			2073 => "0000000010000010110001",
			2074 => "0000000010000010110001",
			2075 => "0010010101101100000100",
			2076 => "0000000010000010110001",
			2077 => "0000000010000010110001",
			2078 => "0011011110011000000100",
			2079 => "0000000010000010110001",
			2080 => "0010100100101100000100",
			2081 => "0000000010000010110001",
			2082 => "0001001010000100000100",
			2083 => "0000000010000010110001",
			2084 => "0000000010000010110001",
			2085 => "0000101101011000001000",
			2086 => "0001100000100100000100",
			2087 => "0000000010000010110001",
			2088 => "0000000010000010110001",
			2089 => "0001100010101000000100",
			2090 => "0000000010000010110001",
			2091 => "0000000010000010110001",
			2092 => "0011100110111000000100",
			2093 => "1111111010000011101101",
			2094 => "0001011001010000011000",
			2095 => "0011011010100100010000",
			2096 => "0011101000110100001100",
			2097 => "0000001010000000000100",
			2098 => "0000000010000011101101",
			2099 => "0000100000000000000100",
			2100 => "0000011010000011101101",
			2101 => "0000010010000011101101",
			2102 => "0000001010000011101101",
			2103 => "0010101000101000000100",
			2104 => "1111111010000011101101",
			2105 => "0000001010000011101101",
			2106 => "1111111010000011101101",
			2107 => "0011100001100000101000",
			2108 => "0010010101010100001100",
			2109 => "0001001110011000001000",
			2110 => "0001111000000000000100",
			2111 => "0000000010000101011001",
			2112 => "0000000010000101011001",
			2113 => "0000000010000101011001",
			2114 => "0011010110110100001100",
			2115 => "0000111101001000001000",
			2116 => "0000111000000000000100",
			2117 => "0000000010000101011001",
			2118 => "0000000010000101011001",
			2119 => "0000000010000101011001",
			2120 => "0000111001010000001000",
			2121 => "0011111000100100000100",
			2122 => "0000000010000101011001",
			2123 => "0000000010000101011001",
			2124 => "0000111000101000000100",
			2125 => "0000000010000101011001",
			2126 => "0000000010000101011001",
			2127 => "0011110011100000001000",
			2128 => "0011010111011100000100",
			2129 => "0000000010000101011001",
			2130 => "0000000010000101011001",
			2131 => "0001100101100100000100",
			2132 => "0000000010000101011001",
			2133 => "0000000010000101011001",
			2134 => "0011000011010000100100",
			2135 => "0001110100101100011100",
			2136 => "0010010101010100001000",
			2137 => "0011100001000100000100",
			2138 => "0000000010000110101101",
			2139 => "0000000010000110101101",
			2140 => "0011010110110100001000",
			2141 => "0000100010101100000100",
			2142 => "0000000010000110101101",
			2143 => "0000000010000110101101",
			2144 => "0000010110010000001000",
			2145 => "0000111100110000000100",
			2146 => "0000000010000110101101",
			2147 => "0000000010000110101101",
			2148 => "0000000010000110101101",
			2149 => "0000000100010100000100",
			2150 => "0000000010000110101101",
			2151 => "0000000010000110101101",
			2152 => "0011110111111100000100",
			2153 => "0000000010000110101101",
			2154 => "0000000010000110101101",
			2155 => "0011100111100000001100",
			2156 => "0011001011101100001000",
			2157 => "0011000110001100000100",
			2158 => "0000000010001000001001",
			2159 => "0000000010001000001001",
			2160 => "0000000010001000001001",
			2161 => "0011100101100000011100",
			2162 => "0000111000101000010100",
			2163 => "0000100011011100000100",
			2164 => "0000000010001000001001",
			2165 => "0000001010010000001000",
			2166 => "0001110110011100000100",
			2167 => "0000000010001000001001",
			2168 => "0000000010001000001001",
			2169 => "0000000010100000000100",
			2170 => "0000000010001000001001",
			2171 => "0000000010001000001001",
			2172 => "0011100100000100000100",
			2173 => "0000000010001000001001",
			2174 => "0000000010001000001001",
			2175 => "0000111001010000000100",
			2176 => "0000000010001000001001",
			2177 => "0000000010001000001001",
			2178 => "0011100110110000000100",
			2179 => "1111111010001001010101",
			2180 => "0000000111111000011000",
			2181 => "0001011111011000000100",
			2182 => "0000000010001001010101",
			2183 => "0011011010100100001000",
			2184 => "0000111100110000000100",
			2185 => "0000000010001001010101",
			2186 => "0000001010001001010101",
			2187 => "0010100100101100000100",
			2188 => "1111111010001001010101",
			2189 => "0011100110000100000100",
			2190 => "0000000010001001010101",
			2191 => "0000001010001001010101",
			2192 => "0001110001010000001000",
			2193 => "0010010101011100000100",
			2194 => "0000001010001001010101",
			2195 => "1111111010001001010101",
			2196 => "1111111010001001010101",
			2197 => "0000111100110000101000",
			2198 => "0010011100101000011100",
			2199 => "0011011011101100010100",
			2200 => "0001010101111000001000",
			2201 => "0010101000000100000100",
			2202 => "0000000010001011000001",
			2203 => "0000000010001011000001",
			2204 => "0001011000000100000100",
			2205 => "0000000010001011000001",
			2206 => "0000001011001100000100",
			2207 => "0000000010001011000001",
			2208 => "0000000010001011000001",
			2209 => "0000110011001000000100",
			2210 => "0000000010001011000001",
			2211 => "0000000010001011000001",
			2212 => "0011011011101100001000",
			2213 => "0001000110000000000100",
			2214 => "0000000010001011000001",
			2215 => "0000000010001011000001",
			2216 => "0000000010001011000001",
			2217 => "0000100011011100000100",
			2218 => "0000000010001011000001",
			2219 => "0001011001010000001000",
			2220 => "0000001010010100000100",
			2221 => "0000000010001011000001",
			2222 => "0000000010001011000001",
			2223 => "0000000010001011000001",
			2224 => "0001101010110000100000",
			2225 => "0001011000000100001100",
			2226 => "0000111000000000001000",
			2227 => "0011001011101100000100",
			2228 => "0000000010001101000101",
			2229 => "0000000010001101000101",
			2230 => "0000000010001101000101",
			2231 => "0000010110010000001000",
			2232 => "0000010111110000000100",
			2233 => "0000000010001101000101",
			2234 => "0000000010001101000101",
			2235 => "0011110010101000000100",
			2236 => "0000000010001101000101",
			2237 => "0011110101100100000100",
			2238 => "0000000010001101000101",
			2239 => "0000000010001101000101",
			2240 => "0011100101100000011000",
			2241 => "0000001010010000001100",
			2242 => "0000111000101000001000",
			2243 => "0001110110011100000100",
			2244 => "0000000010001101000101",
			2245 => "0000000010001101000101",
			2246 => "0000000010001101000101",
			2247 => "0011100101000000000100",
			2248 => "0000000010001101000101",
			2249 => "0011100100000100000100",
			2250 => "0000000010001101000101",
			2251 => "0000000010001101000101",
			2252 => "0000111101001000000100",
			2253 => "0000000010001101000101",
			2254 => "0011100001111000000100",
			2255 => "0000000010001101000101",
			2256 => "0000000010001101000101",
			2257 => "0011100110110000000100",
			2258 => "1111111010001110011001",
			2259 => "0000000111111000011000",
			2260 => "0011100100010000000100",
			2261 => "0000010010001110011001",
			2262 => "0011110010101000001100",
			2263 => "0011110110011000001000",
			2264 => "0011110000001000000100",
			2265 => "1111111010001110011001",
			2266 => "0000001010001110011001",
			2267 => "1111111010001110011001",
			2268 => "0000111100110000000100",
			2269 => "0000000010001110011001",
			2270 => "0000001010001110011001",
			2271 => "0001110001010000001000",
			2272 => "0011101000101100000100",
			2273 => "1111111010001110011001",
			2274 => "0000001010001110011001",
			2275 => "0011100000010000000100",
			2276 => "1111111010001110011001",
			2277 => "0000000010001110011001",
			2278 => "0001100000010000000100",
			2279 => "1111111010001111011101",
			2280 => "0001011001010000011100",
			2281 => "0010111011101100001000",
			2282 => "0001111000101000000100",
			2283 => "0000010010001111011101",
			2284 => "0000001010001111011101",
			2285 => "0000110011100100000100",
			2286 => "1111111010001111011101",
			2287 => "0000001010010100001000",
			2288 => "0000101010101000000100",
			2289 => "0000010010001111011101",
			2290 => "0000001010001111011101",
			2291 => "0011100011101000000100",
			2292 => "1111111010001111011101",
			2293 => "0000000010001111011101",
			2294 => "1111111010001111011101",
			2295 => "0000111100110000101000",
			2296 => "0010010111011100001000",
			2297 => "0010001001001100000100",
			2298 => "0000000010010001001001",
			2299 => "0000000010010001001001",
			2300 => "0000101011100000001000",
			2301 => "0010111110011000000100",
			2302 => "0000000010010001001001",
			2303 => "0000000010010001001001",
			2304 => "0010111011101100001100",
			2305 => "0001011000000100000100",
			2306 => "0000000010010001001001",
			2307 => "0010101001010100000100",
			2308 => "0000000010010001001001",
			2309 => "0000000010010001001001",
			2310 => "0010001111001000000100",
			2311 => "0000000010010001001001",
			2312 => "0010000000110000000100",
			2313 => "0000000010010001001001",
			2314 => "0000000010010001001001",
			2315 => "0000100011011100000100",
			2316 => "0000000010010001001001",
			2317 => "0001011001010000001000",
			2318 => "0011100110110000000100",
			2319 => "0000000010010001001001",
			2320 => "0000000010010001001001",
			2321 => "0000000010010001001001",
			2322 => "0010111011101100010100",
			2323 => "0000000010100100000100",
			2324 => "0000000010010011001101",
			2325 => "0001011000000000001000",
			2326 => "0000010111110000000100",
			2327 => "0000000010010011001101",
			2328 => "0000001010010011001101",
			2329 => "0010101000101000000100",
			2330 => "0000000010010011001101",
			2331 => "0000000010010011001101",
			2332 => "0000101010101000010100",
			2333 => "0000100011011100001100",
			2334 => "0001010011001000001000",
			2335 => "0000111000000000000100",
			2336 => "0000000010010011001101",
			2337 => "0000000010010011001101",
			2338 => "0000000010010011001101",
			2339 => "0001000011000000000100",
			2340 => "0000001010010011001101",
			2341 => "0000000010010011001101",
			2342 => "0000111001010000010000",
			2343 => "0011100101001100001100",
			2344 => "0011100101000000000100",
			2345 => "0000000010010011001101",
			2346 => "0000010101011100000100",
			2347 => "0000000010010011001101",
			2348 => "0000000010010011001101",
			2349 => "1111111010010011001101",
			2350 => "0011101000110100000100",
			2351 => "0000000010010011001101",
			2352 => "0000001101011000000100",
			2353 => "0000000010010011001101",
			2354 => "0000000010010011001101",
			2355 => "0011000011010000101000",
			2356 => "0001111011111000100000",
			2357 => "0010001001000100011000",
			2358 => "0000101011111100001000",
			2359 => "0000111100110000000100",
			2360 => "0000000010010101000001",
			2361 => "0000000010010101000001",
			2362 => "0000010001110000000100",
			2363 => "0000000010010101000001",
			2364 => "0010001001001100000100",
			2365 => "0000000010010101000001",
			2366 => "0010111011101100000100",
			2367 => "0000000010010101000001",
			2368 => "0000000010010101000001",
			2369 => "0001001010000100000100",
			2370 => "0000000010010101000001",
			2371 => "0000000010010101000001",
			2372 => "0001000011010000000100",
			2373 => "0000000010010101000001",
			2374 => "0000000010010101000001",
			2375 => "0000111001010000000100",
			2376 => "0000000010010101000001",
			2377 => "0000111111101000001000",
			2378 => "0011100010110100000100",
			2379 => "0000000010010101000001",
			2380 => "0000000010010101000001",
			2381 => "0001101001111000000100",
			2382 => "0000000010010101000001",
			2383 => "0000000010010101000001",
			2384 => "0011110000001000000100",
			2385 => "1111111010010110011101",
			2386 => "0000000111111000011000",
			2387 => "0000110011100100000100",
			2388 => "1111111010010110011101",
			2389 => "0011011010100100001000",
			2390 => "0000001101011100000100",
			2391 => "0000010010010110011101",
			2392 => "0000001010010110011101",
			2393 => "0000111001010000000100",
			2394 => "1111111010010110011101",
			2395 => "0000000110111100000100",
			2396 => "0000000010010110011101",
			2397 => "0000001010010110011101",
			2398 => "0001001010100100000100",
			2399 => "0000001010010110011101",
			2400 => "0001110001010000001000",
			2401 => "0011001110011000000100",
			2402 => "0000001010010110011101",
			2403 => "1111111010010110011101",
			2404 => "0001011100110000000100",
			2405 => "1111111010010110011101",
			2406 => "1111111010010110011101",
			2407 => "0001011000000100010100",
			2408 => "0000110011100100001000",
			2409 => "0011001011101100000100",
			2410 => "0000000010011000100001",
			2411 => "0000000010011000100001",
			2412 => "0000000010101100001000",
			2413 => "0000011000011000000100",
			2414 => "0000000010011000100001",
			2415 => "0000000010011000100001",
			2416 => "0000000010011000100001",
			2417 => "0011110011100000101000",
			2418 => "0011110000100100010100",
			2419 => "0000010110010000001000",
			2420 => "0000010111110000000100",
			2421 => "0000000010011000100001",
			2422 => "0000000010011000100001",
			2423 => "0000111001010000000100",
			2424 => "0000000010011000100001",
			2425 => "0010100100101100000100",
			2426 => "0000000010011000100001",
			2427 => "0000000010011000100001",
			2428 => "0011011010100100001000",
			2429 => "0000001110110000000100",
			2430 => "0000000010011000100001",
			2431 => "0000000010011000100001",
			2432 => "0010100100101100000100",
			2433 => "0000000010011000100001",
			2434 => "0001000011000000000100",
			2435 => "0000000010011000100001",
			2436 => "0000000010011000100001",
			2437 => "0010101011111000000100",
			2438 => "0000000010011000100001",
			2439 => "0000000010011000100001",
			2440 => "0011100111100000001100",
			2441 => "0011011101000000001000",
			2442 => "0000111100010000000100",
			2443 => "0000000010011010000101",
			2444 => "0000000010011010000101",
			2445 => "0000000010011010000101",
			2446 => "0000110011100100000100",
			2447 => "0000000010011010000101",
			2448 => "0000111000101000011000",
			2449 => "0011100101100000010000",
			2450 => "0001001001000100000100",
			2451 => "0000000010011010000101",
			2452 => "0010001111001000000100",
			2453 => "0000000010011010000101",
			2454 => "0001110000111100000100",
			2455 => "0000000010011010000101",
			2456 => "0000000010011010000101",
			2457 => "0011010011010000000100",
			2458 => "0000000010011010000101",
			2459 => "0000000010011010000101",
			2460 => "0011100100000100000100",
			2461 => "0000000010011010000101",
			2462 => "0000001010111000000100",
			2463 => "0000000010011010000101",
			2464 => "0000000010011010000101",
			2465 => "0000011000011000101000",
			2466 => "0000010111110000001100",
			2467 => "0001001101000000000100",
			2468 => "0000000010011100001001",
			2469 => "0001111011111000000100",
			2470 => "0000000010011100001001",
			2471 => "0000000010011100001001",
			2472 => "0010001001001100000100",
			2473 => "0000000010011100001001",
			2474 => "0010100100101100001100",
			2475 => "0011110000001000000100",
			2476 => "0000000010011100001001",
			2477 => "0000110011100100000100",
			2478 => "0000000010011100001001",
			2479 => "0000000010011100001001",
			2480 => "0001110100101100000100",
			2481 => "0000000010011100001001",
			2482 => "0010001111001000000100",
			2483 => "0000000010011100001001",
			2484 => "0000000010011100001001",
			2485 => "0010100100101100010100",
			2486 => "0010010101010100000100",
			2487 => "0000000010011100001001",
			2488 => "0010010101101100000100",
			2489 => "0000000010011100001001",
			2490 => "0010110011010000001000",
			2491 => "0010001111001000000100",
			2492 => "0000000010011100001001",
			2493 => "0000000010011100001001",
			2494 => "0000000010011100001001",
			2495 => "0001011000101000000100",
			2496 => "0000000010011100001001",
			2497 => "0000000010011100001001",
			2498 => "0000000111111000110000",
			2499 => "0001110001010000010000",
			2500 => "0011010110110100001000",
			2501 => "0001110110101100000100",
			2502 => "0000000010011110010101",
			2503 => "0000000010011110010101",
			2504 => "0010010101010100000100",
			2505 => "0000000010011110010101",
			2506 => "0000000010011110010101",
			2507 => "0000110011100100000100",
			2508 => "0000000010011110010101",
			2509 => "0011011010100100001100",
			2510 => "0000010111100100000100",
			2511 => "0000000010011110010101",
			2512 => "0011110000001000000100",
			2513 => "0000000010011110010101",
			2514 => "0000000010011110010101",
			2515 => "0010001001000100000100",
			2516 => "0000000010011110010101",
			2517 => "0000010110001100001000",
			2518 => "0010101011000000000100",
			2519 => "0000000010011110010101",
			2520 => "0000000010011110010101",
			2521 => "0000000010011110010101",
			2522 => "0001110001010000010000",
			2523 => "0010010101011100001000",
			2524 => "0001011000000000000100",
			2525 => "0000000010011110010101",
			2526 => "0000000010011110010101",
			2527 => "0000000101101000000100",
			2528 => "0000000010011110010101",
			2529 => "0000000010011110010101",
			2530 => "0011101000010100000100",
			2531 => "0000000010011110010101",
			2532 => "0000000010011110010101",
			2533 => "0001011000000100011000",
			2534 => "0000010001110000000100",
			2535 => "0000000010100000110001",
			2536 => "0000000010101100001000",
			2537 => "0001011111011000000100",
			2538 => "0000000010100000110001",
			2539 => "0000000010100000110001",
			2540 => "0000110011100100001000",
			2541 => "0000110011000000000100",
			2542 => "0000000010100000110001",
			2543 => "0000000010100000110001",
			2544 => "0000000010100000110001",
			2545 => "0010101111101000011000",
			2546 => "0010011001001000001100",
			2547 => "0011110110011000001000",
			2548 => "0011110111010000000100",
			2549 => "0000000010100000110001",
			2550 => "0000000010100000110001",
			2551 => "0000000010100000110001",
			2552 => "0001011100110000001000",
			2553 => "0001011000111000000100",
			2554 => "0000000010100000110001",
			2555 => "0000000010100000110001",
			2556 => "0000000010100000110001",
			2557 => "0000000111111000010100",
			2558 => "0011010011010000001000",
			2559 => "0011110000100100000100",
			2560 => "0000000010100000110001",
			2561 => "0000000010100000110001",
			2562 => "0000010110001100000100",
			2563 => "0000000010100000110001",
			2564 => "0000011011101100000100",
			2565 => "0000000010100000110001",
			2566 => "0000000010100000110001",
			2567 => "0001110001010000001000",
			2568 => "0011111101001100000100",
			2569 => "0000000010100000110001",
			2570 => "0000000010100000110001",
			2571 => "0000000010100000110001",
			2572 => "0000100011011100000100",
			2573 => "1111111010100010000101",
			2574 => "0001011001010000100100",
			2575 => "0000111100110000011000",
			2576 => "0010010101010100001000",
			2577 => "0000010001110000000100",
			2578 => "1111111010100010000101",
			2579 => "0000001010100010000101",
			2580 => "0011100001100000001100",
			2581 => "0010101000101000001000",
			2582 => "0000100100010100000100",
			2583 => "1111111010100010000101",
			2584 => "1111111010100010000101",
			2585 => "1111111010100010000101",
			2586 => "0000000010100010000101",
			2587 => "0000001010010100001000",
			2588 => "0000111001010000000100",
			2589 => "0000001010100010000101",
			2590 => "0000001010100010000101",
			2591 => "0000000010100010000101",
			2592 => "1111111010100010000101",
			2593 => "0011100110110000000100",
			2594 => "1111111010100011001001",
			2595 => "0001110011000100011100",
			2596 => "0000110011001000000100",
			2597 => "0000000010100011001001",
			2598 => "0000010111110000000100",
			2599 => "1111111010100011001001",
			2600 => "0001111000101000000100",
			2601 => "0000001010100011001001",
			2602 => "0001111011111000001000",
			2603 => "0011110100110100000100",
			2604 => "0000000010100011001001",
			2605 => "0000000010100011001001",
			2606 => "0011000011010000000100",
			2607 => "0000001010100011001001",
			2608 => "0000000010100011001001",
			2609 => "1111111010100011001001",
			2610 => "0011110000001000000100",
			2611 => "1111111010100100101101",
			2612 => "0000000111111000011000",
			2613 => "0001011111011000000100",
			2614 => "0000000010100100101101",
			2615 => "0011011010100100001000",
			2616 => "0000000100010100000100",
			2617 => "0000001010100100101101",
			2618 => "0000000010100100101101",
			2619 => "0010100100101100000100",
			2620 => "1111111010100100101101",
			2621 => "0000000000101000000100",
			2622 => "0000000010100100101101",
			2623 => "0000000010100100101101",
			2624 => "0001010101111000000100",
			2625 => "0000000010100100101101",
			2626 => "0011101000010100010000",
			2627 => "0001110001010000001100",
			2628 => "0011010110001100000100",
			2629 => "1111111010100100101101",
			2630 => "0010111110011000000100",
			2631 => "0000001010100100101101",
			2632 => "0000000010100100101101",
			2633 => "1111111010100100101101",
			2634 => "0000000010100100101101",
			2635 => "0011110000001000000100",
			2636 => "1111111010100101111001",
			2637 => "0000010111110000000100",
			2638 => "1111111010100101111001",
			2639 => "0011010110001100000100",
			2640 => "0000001010100101111001",
			2641 => "0000001010010000010100",
			2642 => "0011011011101100000100",
			2643 => "0000000010100101111001",
			2644 => "0011011010100100001000",
			2645 => "0010101111101000000100",
			2646 => "0000000010100101111001",
			2647 => "0000001010100101111001",
			2648 => "0011100100000100000100",
			2649 => "1111111010100101111001",
			2650 => "0000000010100101111001",
			2651 => "0001100010101000000100",
			2652 => "1111111010100101111001",
			2653 => "0000000010100101111001",
			2654 => "0000100011011100000100",
			2655 => "0000000010100111010101",
			2656 => "0000101101110000100100",
			2657 => "0001110011000100100000",
			2658 => "0000110011001000001000",
			2659 => "0010010101010100000100",
			2660 => "0000000010100111010101",
			2661 => "0000000010100111010101",
			2662 => "0000111000101000001100",
			2663 => "0000010111110000000100",
			2664 => "0000000010100111010101",
			2665 => "0011100110110000000100",
			2666 => "0000000010100111010101",
			2667 => "0000000010100111010101",
			2668 => "0001111100101100000100",
			2669 => "0000000010100111010101",
			2670 => "0000111011111000000100",
			2671 => "0000000010100111010101",
			2672 => "0000000010100111010101",
			2673 => "0000000010100111010101",
			2674 => "0011110101011000000100",
			2675 => "0000000010100111010101",
			2676 => "0000000010100111010101",
			2677 => "0010010101010100001100",
			2678 => "0000010001110000000100",
			2679 => "0000000010101001001001",
			2680 => "0011111000001000000100",
			2681 => "0000000010101001001001",
			2682 => "0000001010101001001001",
			2683 => "0000101101110000101100",
			2684 => "0011010110001100001000",
			2685 => "0011001110011000000100",
			2686 => "0000001010101001001001",
			2687 => "0000000010101001001001",
			2688 => "0001111011111000010100",
			2689 => "0000111100010000001000",
			2690 => "0000001101111000000100",
			2691 => "1111111010101001001001",
			2692 => "0000000010101001001001",
			2693 => "0000111000101000001000",
			2694 => "0000010001100100000100",
			2695 => "0000000010101001001001",
			2696 => "0000000010101001001001",
			2697 => "1111111010101001001001",
			2698 => "0001110011000100001100",
			2699 => "0000010111100100000100",
			2700 => "0000000010101001001001",
			2701 => "0011010011010000000100",
			2702 => "0000001010101001001001",
			2703 => "0000000010101001001001",
			2704 => "1111111010101001001001",
			2705 => "1111111010101001001001",
			2706 => "0000110011100100001100",
			2707 => "0010010101010100001000",
			2708 => "0001111100010000000100",
			2709 => "0000000010101011010101",
			2710 => "0000000010101011010101",
			2711 => "1111111010101011010101",
			2712 => "0000010111100100001000",
			2713 => "0001011000000100000100",
			2714 => "0000000010101011010101",
			2715 => "0000000010101011010101",
			2716 => "0000011000011000010100",
			2717 => "0010100100101100001000",
			2718 => "0001011100010000000100",
			2719 => "0000001010101011010101",
			2720 => "0000000010101011010101",
			2721 => "0001110100101100000100",
			2722 => "0000000010101011010101",
			2723 => "0010001010000100000100",
			2724 => "0000000010101011010101",
			2725 => "0000000010101011010101",
			2726 => "0001000111011100001000",
			2727 => "0000010011110000000100",
			2728 => "0000000010101011010101",
			2729 => "0000000010101011010101",
			2730 => "0000101010101000001000",
			2731 => "0000100111011000000100",
			2732 => "0000000010101011010101",
			2733 => "0000000010101011010101",
			2734 => "0001111111101000001000",
			2735 => "0000001011001100000100",
			2736 => "0000000010101011010101",
			2737 => "0000000010101011010101",
			2738 => "0000010110001100000100",
			2739 => "0000000010101011010101",
			2740 => "0000000010101011010101",
			2741 => "0001111011111000111000",
			2742 => "0010010111011100001000",
			2743 => "0011011111011100000100",
			2744 => "0000000010101110000001",
			2745 => "0000000010101110000001",
			2746 => "0011011110011000100000",
			2747 => "0011010110001100010100",
			2748 => "0010101111101000001100",
			2749 => "0000111100010000001000",
			2750 => "0001001101000000000100",
			2751 => "0000000010101110000001",
			2752 => "0000000010101110000001",
			2753 => "0000000010101110000001",
			2754 => "0010100100101100000100",
			2755 => "0000000010101110000001",
			2756 => "0000000010101110000001",
			2757 => "0001010101111000001000",
			2758 => "0001011101101000000100",
			2759 => "0000000010101110000001",
			2760 => "0000000010101110000001",
			2761 => "0000000010101110000001",
			2762 => "0010101000101000001000",
			2763 => "0001001110011000000100",
			2764 => "0000000010101110000001",
			2765 => "0000000010101110000001",
			2766 => "0001001001000100000100",
			2767 => "0000000010101110000001",
			2768 => "0000000010101110000001",
			2769 => "0000000111111000011100",
			2770 => "0001111011000000001100",
			2771 => "0001011001010000001000",
			2772 => "0010101001010100000100",
			2773 => "0000000010101110000001",
			2774 => "0000000010101110000001",
			2775 => "0000000010101110000001",
			2776 => "0000111001010000000100",
			2777 => "0000000010101110000001",
			2778 => "0010001001000100000100",
			2779 => "0000000010101110000001",
			2780 => "0001001000000100000100",
			2781 => "0000000010101110000001",
			2782 => "0000000010101110000001",
			2783 => "0000000010101110000001",
			2784 => "0000010111110000000100",
			2785 => "1111111010110000000111",
			2786 => "0011010110001100001100",
			2787 => "0001011000111000001000",
			2788 => "0011101110100000000100",
			2789 => "0000000010110000000111",
			2790 => "0000001010110000000111",
			2791 => "0000000010110000000111",
			2792 => "0001111011111000100000",
			2793 => "0000010110010000001000",
			2794 => "0001000101101100000100",
			2795 => "0000001010110000000111",
			2796 => "0000000010110000000111",
			2797 => "0010011001001000001100",
			2798 => "0000000100010100000100",
			2799 => "1111111010110000000111",
			2800 => "0000001110110000000100",
			2801 => "0000000010110000000111",
			2802 => "0000000010110000000111",
			2803 => "0010111010100100001000",
			2804 => "0000111100110000000100",
			2805 => "0000000010110000000111",
			2806 => "0000000010110000000111",
			2807 => "0000000010110000000111",
			2808 => "0001110011000100010000",
			2809 => "0000010111100100000100",
			2810 => "0000000010110000000111",
			2811 => "0010101001010100000100",
			2812 => "0000000010110000000111",
			2813 => "0000000111111000000100",
			2814 => "0000001010110000000111",
			2815 => "0000000010110000000111",
			2816 => "1111111010110000000111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(953, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1881, initial_addr_3'length));
	end generate gen_rom_6;

	gen_rom_7: if SELECT_ROM = 7 generate
		bank <= (
			0 => "0000100111000100100100",
			1 => "0000000111110100011100",
			2 => "0000011001100100000100",
			3 => "1111111000000001011101",
			4 => "0011100110100000010000",
			5 => "0001100010000000001100",
			6 => "0000000100111100001000",
			7 => "0001111001010100000100",
			8 => "0000000000000001011101",
			9 => "0000000000000001011101",
			10 => "1111111000000001011101",
			11 => "0000000000000001011101",
			12 => "0010111110011000000100",
			13 => "0000000000000001011101",
			14 => "1111111000000001011101",
			15 => "0011101111110000000100",
			16 => "0000001000000001011101",
			17 => "0000000000000001011101",
			18 => "0000010000011000001000",
			19 => "0011011011101100000100",
			20 => "0000000000000001011101",
			21 => "0000000000000001011101",
			22 => "1111111000000001011101",
			23 => "0001101111010100101000",
			24 => "0000000000011100100000",
			25 => "0011111110100000011100",
			26 => "0001100000110100010100",
			27 => "0001101111000100001100",
			28 => "0001100110100000001000",
			29 => "0000000010111100000100",
			30 => "0000000000000011000001",
			31 => "0000000000000011000001",
			32 => "0000001000000011000001",
			33 => "0001000000111100000100",
			34 => "0000000000000011000001",
			35 => "0000000000000011000001",
			36 => "0000001011011000000100",
			37 => "0000000000000011000001",
			38 => "0000000000000011000001",
			39 => "0000000000000011000001",
			40 => "0001111001010100000100",
			41 => "0000000000000011000001",
			42 => "0000000000000011000001",
			43 => "0000010111110000001000",
			44 => "0010110011010000000100",
			45 => "0000000000000011000001",
			46 => "0000000000000011000001",
			47 => "1111111000000011000001",
			48 => "0011101110111100101000",
			49 => "0001000010111000100000",
			50 => "0001001100001100011100",
			51 => "0011001011101100001000",
			52 => "0010001001001100000100",
			53 => "0000000000000100010101",
			54 => "0000001000000100010101",
			55 => "0001000111011100000100",
			56 => "1111111000000100010101",
			57 => "0000111110111000001000",
			58 => "0010101010011100000100",
			59 => "0000000000000100010101",
			60 => "0000001000000100010101",
			61 => "0001001110111000000100",
			62 => "1111111000000100010101",
			63 => "0000000000000100010101",
			64 => "1111111000000100010101",
			65 => "0001111000101000000100",
			66 => "0000001000000100010101",
			67 => "1111111000000100010101",
			68 => "1111111000000100010101",
			69 => "0000101000010100111000",
			70 => "0011101010100000101000",
			71 => "0000000011101100011000",
			72 => "0011000101011100010000",
			73 => "0010000011010000000100",
			74 => "0000000000000111100001",
			75 => "0001011001100000000100",
			76 => "0000000000000111100001",
			77 => "0000010001110000000100",
			78 => "0000000000000111100001",
			79 => "0000000000000111100001",
			80 => "0000010011010000000100",
			81 => "0000000000000111100001",
			82 => "0000000000000111100001",
			83 => "0000011000011000001000",
			84 => "0011100010001100000100",
			85 => "0000000000000111100001",
			86 => "0000000000000111100001",
			87 => "0011100001101000000100",
			88 => "0000000000000111100001",
			89 => "0000000000000111100001",
			90 => "0011010101011100001100",
			91 => "0010001111111100001000",
			92 => "0001101111111000000100",
			93 => "0000000000000111100001",
			94 => "0000000000000111100001",
			95 => "0000000000000111100001",
			96 => "0000000000000111100001",
			97 => "0011101010011000001100",
			98 => "0000010110001100001000",
			99 => "0000000010111100000100",
			100 => "0000000000000111100001",
			101 => "0000000000000111100001",
			102 => "0000000000000111100001",
			103 => "0001101111010100011000",
			104 => "0010001111001000010000",
			105 => "0010001111111100001000",
			106 => "0010000101011100000100",
			107 => "0000000000000111100001",
			108 => "0000000000000111100001",
			109 => "0000111110111000000100",
			110 => "0000000000000111100001",
			111 => "0000000000000111100001",
			112 => "0011110010001000000100",
			113 => "0000000000000111100001",
			114 => "0000000000000111100001",
			115 => "0000011000111100001000",
			116 => "0001011001010000000100",
			117 => "0000000000000111100001",
			118 => "0000000000000111100001",
			119 => "0000000000000111100001",
			120 => "0001100100010000111000",
			121 => "0001010110001100001100",
			122 => "0001001001100100000100",
			123 => "0000000000001001010101",
			124 => "0000010011110000000100",
			125 => "1111111000001001010101",
			126 => "0000000000001001010101",
			127 => "0010001001001100010100",
			128 => "0001101010011000010000",
			129 => "0001101001111100001100",
			130 => "0001011001001000000100",
			131 => "0000000000001001010101",
			132 => "0000001110010000000100",
			133 => "1111111000001001010101",
			134 => "0000000000001001010101",
			135 => "0000000000001001010101",
			136 => "1111111000001001010101",
			137 => "0011001010100100001000",
			138 => "0010001111111100000100",
			139 => "0000000000001001010101",
			140 => "0000001000001001010101",
			141 => "0001011000000100000100",
			142 => "1111111000001001010101",
			143 => "0001100110110000001000",
			144 => "0001101111010100000100",
			145 => "0000000000001001010101",
			146 => "1111111000001001010101",
			147 => "0000001000001001010101",
			148 => "1111111000001001010101",
			149 => "0001011100001100111000",
			150 => "0010110111011100110000",
			151 => "0010001111111100010000",
			152 => "0011000110110100000100",
			153 => "0000000000001100010001",
			154 => "0011111100000100000100",
			155 => "0000000000001100010001",
			156 => "0000111111101000000100",
			157 => "0000000000001100010001",
			158 => "0000000000001100010001",
			159 => "0011010011010000011000",
			160 => "0011011011101100001100",
			161 => "0000101001111100000100",
			162 => "0000000000001100010001",
			163 => "0011100000010100000100",
			164 => "0000000000001100010001",
			165 => "0000000000001100010001",
			166 => "0000010110010000000100",
			167 => "0000000000001100010001",
			168 => "0001100011101100000100",
			169 => "0000000000001100010001",
			170 => "0000000000001100010001",
			171 => "0000001011101000000100",
			172 => "0000000000001100010001",
			173 => "0000000000001100010001",
			174 => "0010000101011100000100",
			175 => "0000000000001100010001",
			176 => "0000000000001100010001",
			177 => "0010101100110100011100",
			178 => "0010110101010100001100",
			179 => "0000111000100000001000",
			180 => "0010010110000000000100",
			181 => "0000000000001100010001",
			182 => "0000000000001100010001",
			183 => "0000000000001100010001",
			184 => "0000010001110000000100",
			185 => "0000000000001100010001",
			186 => "0001110001010000001000",
			187 => "0000110001001000000100",
			188 => "0000000000001100010001",
			189 => "0000000000001100010001",
			190 => "0000000000001100010001",
			191 => "0001111001010000000100",
			192 => "0000000000001100010001",
			193 => "0010011000000100000100",
			194 => "0000000000001100010001",
			195 => "0000000000001100010001",
			196 => "0000000100011000111100",
			197 => "0011101111100100101100",
			198 => "0010001001000100100000",
			199 => "0010101011000000010100",
			200 => "0011100001101000001100",
			201 => "0001110011010000000100",
			202 => "0000000000001111110101",
			203 => "0000010111100100000100",
			204 => "0000000000001111110101",
			205 => "0000000000001111110101",
			206 => "0001011000111000000100",
			207 => "0000000000001111110101",
			208 => "0000000000001111110101",
			209 => "0000111001000000001000",
			210 => "0011000111011100000100",
			211 => "0000000000001111110101",
			212 => "0000000000001111110101",
			213 => "0000000000001111110101",
			214 => "0001001000000000001000",
			215 => "0010110111011100000100",
			216 => "0000000000001111110101",
			217 => "0000000000001111110101",
			218 => "0000000000001111110101",
			219 => "0010000101011100001000",
			220 => "0000001101010000000100",
			221 => "0000000000001111110101",
			222 => "0000000000001111110101",
			223 => "0010001111001000000100",
			224 => "0000000000001111110101",
			225 => "0000000000001111110101",
			226 => "0011101010011000010000",
			227 => "0000010110001100001100",
			228 => "0001111101001000000100",
			229 => "0000000000001111110101",
			230 => "0001111001010000000100",
			231 => "0000000000001111110101",
			232 => "0000000000001111110101",
			233 => "0000000000001111110101",
			234 => "0011100110100000010100",
			235 => "0010001111111100001000",
			236 => "0010110111011100000100",
			237 => "0000000000001111110101",
			238 => "0000000000001111110101",
			239 => "0011110101110100001000",
			240 => "0001101001011100000100",
			241 => "0000000000001111110101",
			242 => "0000000000001111110101",
			243 => "0000000000001111110101",
			244 => "0000011000111100001000",
			245 => "0010111110011000000100",
			246 => "0000000000001111110101",
			247 => "0000000000001111110101",
			248 => "0001011110010100000100",
			249 => "0000000000001111110101",
			250 => "0001010001011100000100",
			251 => "0000000000001111110101",
			252 => "0000000000001111110101",
			253 => "0001100100010000111000",
			254 => "0011001001001000101000",
			255 => "0000011001100100001000",
			256 => "0011100000010100000100",
			257 => "1111111000010001101001",
			258 => "0000001000010001101001",
			259 => "0010101100110100011100",
			260 => "0000101100111000010000",
			261 => "0011101101111100001000",
			262 => "0000001100000100000100",
			263 => "0000001000010001101001",
			264 => "1111111000010001101001",
			265 => "0011110000010100000100",
			266 => "0000001000010001101001",
			267 => "0000000000010001101001",
			268 => "0011101001111100000100",
			269 => "1111111000010001101001",
			270 => "0010101011000000000100",
			271 => "0000000000010001101001",
			272 => "0000001000010001101001",
			273 => "1111111000010001101001",
			274 => "0001010010111000000100",
			275 => "1111111000010001101001",
			276 => "0000001011000100001000",
			277 => "0011101011110000000100",
			278 => "0000000000010001101001",
			279 => "0000001000010001101001",
			280 => "1111111000010001101001",
			281 => "1111111000010001101001",
			282 => "0000100111010001000100",
			283 => "0001010101111000010100",
			284 => "0011001011101100001000",
			285 => "0000001110010100000100",
			286 => "0000100000010100011101",
			287 => "0000010000010100011101",
			288 => "0011001110011000000100",
			289 => "0000001000010100011101",
			290 => "0011001010100100000100",
			291 => "0000000000010100011101",
			292 => "1111111000010100011101",
			293 => "0010001111111100010000",
			294 => "0011011011101100001000",
			295 => "0001000110011100000100",
			296 => "1111111000010100011101",
			297 => "0000000000010100011101",
			298 => "0001011110001100000100",
			299 => "0000000000010100011101",
			300 => "0000010000010100011101",
			301 => "0010110101101100011100",
			302 => "0000010111100100010000",
			303 => "0011100010001100001000",
			304 => "0010101001010100000100",
			305 => "0000010000010100011101",
			306 => "1111111000010100011101",
			307 => "0000000000001100000100",
			308 => "0000011000010100011101",
			309 => "0000001000010100011101",
			310 => "0000110001001000001000",
			311 => "0000000111101000000100",
			312 => "0000011000010100011101",
			313 => "0000001000010100011101",
			314 => "0000101000010100011101",
			315 => "1111111000010100011101",
			316 => "0011101110111100010100",
			317 => "0011110100101000010000",
			318 => "0010101101001000000100",
			319 => "0000001000010100011101",
			320 => "0010100001101000001000",
			321 => "0001001001000000000100",
			322 => "1111111000010100011101",
			323 => "0000001000010100011101",
			324 => "1111111000010100011101",
			325 => "0000010000010100011101",
			326 => "1111111000010100011101",
			327 => "0000100111010001000100",
			328 => "0001010011000000010000",
			329 => "0011001110011000001100",
			330 => "0010000011010000000100",
			331 => "1111111000010111011001",
			332 => "0011000110110100000100",
			333 => "0000010000010111011001",
			334 => "0000001000010111011001",
			335 => "1111111000010111011001",
			336 => "0000010110010000011000",
			337 => "0011011011101100001100",
			338 => "0000111011000000001000",
			339 => "0010000101011100000100",
			340 => "1111111000010111011001",
			341 => "0000001000010111011001",
			342 => "1111111000010111011001",
			343 => "0001011110001100000100",
			344 => "0000000000010111011001",
			345 => "0000000100100000000100",
			346 => "0000010000010111011001",
			347 => "0000000000010111011001",
			348 => "0011000110000000011000",
			349 => "0011000011010000001000",
			350 => "0000011001100000000100",
			351 => "0000010000010111011001",
			352 => "0000010000010111011001",
			353 => "0001011001011000001000",
			354 => "0010110111011100000100",
			355 => "0000001000010111011001",
			356 => "1111111000010111011001",
			357 => "0011101111100100000100",
			358 => "0000001000010111011001",
			359 => "0000010000010111011001",
			360 => "1111111000010111011001",
			361 => "0011101110111100011000",
			362 => "0011110100001100001000",
			363 => "0000001101001100000100",
			364 => "0000000000010111011001",
			365 => "1111111000010111011001",
			366 => "0001111000101000001100",
			367 => "0010001111111100001000",
			368 => "0011000101010100000100",
			369 => "1111111000010111011001",
			370 => "0000001000010111011001",
			371 => "0000010000010111011001",
			372 => "1111111000010111011001",
			373 => "1111111000010111011001",
			374 => "0000000100011000111100",
			375 => "0011101111100100101100",
			376 => "0010001001000100100000",
			377 => "0010101011000000010100",
			378 => "0001011001010100001100",
			379 => "0011000110110100000100",
			380 => "0000000000011010110101",
			381 => "0000010001100100000100",
			382 => "0000000000011010110101",
			383 => "0000000000011010110101",
			384 => "0010010101101100000100",
			385 => "0000000000011010110101",
			386 => "0000000000011010110101",
			387 => "0000111001000000001000",
			388 => "0011000111011100000100",
			389 => "0000000000011010110101",
			390 => "0000000000011010110101",
			391 => "0000000000011010110101",
			392 => "0001001000000000001000",
			393 => "0010110111011100000100",
			394 => "0000000000011010110101",
			395 => "0000000000011010110101",
			396 => "0000000000011010110101",
			397 => "0010000101011100001000",
			398 => "0000001101010000000100",
			399 => "0000000000011010110101",
			400 => "0000000000011010110101",
			401 => "0010001111001000000100",
			402 => "0000000000011010110101",
			403 => "0000000000011010110101",
			404 => "0000011000111100001100",
			405 => "0011101001110000000100",
			406 => "0000000000011010110101",
			407 => "0000001000010000000100",
			408 => "0000000000011010110101",
			409 => "0000000000011010110101",
			410 => "0001000101010100001000",
			411 => "0000000011100000000100",
			412 => "0000000000011010110101",
			413 => "0000000000011010110101",
			414 => "0000010000011000001000",
			415 => "0001100011010100000100",
			416 => "0000000000011010110101",
			417 => "0000000000011010110101",
			418 => "0001101111000100001100",
			419 => "0001100110100000001000",
			420 => "0011101111111000000100",
			421 => "0000000000011010110101",
			422 => "0000000000011010110101",
			423 => "0000000000011010110101",
			424 => "0001101111110100000100",
			425 => "0000000000011010110101",
			426 => "0001101111010100000100",
			427 => "0000000000011010110101",
			428 => "0000000000011010110101",
			429 => "0000001100000100110100",
			430 => "0001011100001100101100",
			431 => "0010111010100100011000",
			432 => "0010000101011100001100",
			433 => "0000001001000000000100",
			434 => "0000000000011110000001",
			435 => "0011010110110100000100",
			436 => "1111111000011110000001",
			437 => "0000000000011110000001",
			438 => "0001000110001100000100",
			439 => "0000000000011110000001",
			440 => "0000100011010100000100",
			441 => "0000001000011110000001",
			442 => "0000000000011110000001",
			443 => "0011011010100100001000",
			444 => "0000011000011000000100",
			445 => "1111111000011110000001",
			446 => "0000000000011110000001",
			447 => "0011101001000000000100",
			448 => "1111111000011110000001",
			449 => "0001010100101100000100",
			450 => "0000000000011110000001",
			451 => "0000000000011110000001",
			452 => "0011000101010100000100",
			453 => "0000000000011110000001",
			454 => "0000001000011110000001",
			455 => "0001000010111000101100",
			456 => "0011101101111100001000",
			457 => "0010000000110000000100",
			458 => "1111111000011110000001",
			459 => "0000000000011110000001",
			460 => "0000000100100000001100",
			461 => "0001011110111000000100",
			462 => "0000000000011110000001",
			463 => "0011100101110000000100",
			464 => "0000000000011110000001",
			465 => "0000001000011110000001",
			466 => "0011100010011100001000",
			467 => "0010111001001000000100",
			468 => "1111111000011110000001",
			469 => "0000000000011110000001",
			470 => "0001101111000100001000",
			471 => "0000010110010000000100",
			472 => "0000000000011110000001",
			473 => "0000000000011110000001",
			474 => "0001100010000000000100",
			475 => "1111111000011110000001",
			476 => "0000000000011110000001",
			477 => "0000110001101000000100",
			478 => "0000001000011110000001",
			479 => "1111111000011110000001",
			480 => "0010001001000101010000",
			481 => "0011100010011100101100",
			482 => "0000001100000100011000",
			483 => "0011100010001100010100",
			484 => "0010110110001100001000",
			485 => "0000001110010100000100",
			486 => "0000000000100010000101",
			487 => "0000000000100010000101",
			488 => "0000010111100100000100",
			489 => "0000000000100010000101",
			490 => "0010111010100100000100",
			491 => "0000000000100010000101",
			492 => "0000000000100010000101",
			493 => "0000000000100010000101",
			494 => "0010101010011100010000",
			495 => "0001111000111000001100",
			496 => "0000111100101100001000",
			497 => "0001111000000100000100",
			498 => "0000000000100010000101",
			499 => "0000000000100010000101",
			500 => "0000000000100010000101",
			501 => "0000000000100010000101",
			502 => "0000000000100010000101",
			503 => "0001010011000100001100",
			504 => "0000011000011000000100",
			505 => "0000000000100010000101",
			506 => "0001111100110000000100",
			507 => "0000000000100010000101",
			508 => "0000000000100010000101",
			509 => "0000111110111000001100",
			510 => "0010001001001100000100",
			511 => "0000000000100010000101",
			512 => "0000100111000100000100",
			513 => "0000000000100010000101",
			514 => "0000000000100010000101",
			515 => "0000000100111100001000",
			516 => "0000111110001100000100",
			517 => "0000000000100010000101",
			518 => "0000000000100010000101",
			519 => "0000000000100010000101",
			520 => "0001101010011000011100",
			521 => "0011011001001000010100",
			522 => "0001010110000000001100",
			523 => "0000001000100000001000",
			524 => "0001010101011100000100",
			525 => "0000000000100010000101",
			526 => "0000000000100010000101",
			527 => "0000000000100010000101",
			528 => "0010111100101000000100",
			529 => "0000001000100010000101",
			530 => "0000000000100010000101",
			531 => "0001001000111000000100",
			532 => "0000000000100010000101",
			533 => "0000000000100010000101",
			534 => "0010101101001000001000",
			535 => "0010101100010000000100",
			536 => "0000000000100010000101",
			537 => "0000000000100010000101",
			538 => "0011111110111100001000",
			539 => "0010110011000000000100",
			540 => "0000000000100010000101",
			541 => "0000000000100010000101",
			542 => "0001011101101100000100",
			543 => "0000000000100010000101",
			544 => "0000000000100010000101",
			545 => "0011101110111101010000",
			546 => "0011001001001000111100",
			547 => "0000011000011000101000",
			548 => "0011101010100000010000",
			549 => "0010110110001100000100",
			550 => "0000001000100100110001",
			551 => "0001010101101100000100",
			552 => "1111111000100100110001",
			553 => "0001111010000100000100",
			554 => "0000001000100100110001",
			555 => "0000000000100100110001",
			556 => "0011011011101100001100",
			557 => "0010110011010000001000",
			558 => "0001000110101100000100",
			559 => "0000000000100100110001",
			560 => "0000001000100100110001",
			561 => "1111111000100100110001",
			562 => "0010110011010000000100",
			563 => "0000000000100100110001",
			564 => "0010100000111100000100",
			565 => "0000001000100100110001",
			566 => "0000001000100100110001",
			567 => "0011111010011000001100",
			568 => "0001011011101100000100",
			569 => "0000000000100100110001",
			570 => "0001001011101100000100",
			571 => "0000001000100100110001",
			572 => "0000001000100100110001",
			573 => "0010001111001000000100",
			574 => "0000001000100100110001",
			575 => "0000000000100100110001",
			576 => "0001010010111000001000",
			577 => "0001010001001000000100",
			578 => "1111111000100100110001",
			579 => "1111111000100100110001",
			580 => "0000001011000100001000",
			581 => "0011101011110000000100",
			582 => "0000000000100100110001",
			583 => "0000001000100100110001",
			584 => "1111111000100100110001",
			585 => "0000000101111100000100",
			586 => "0000000000100100110001",
			587 => "1111111000100100110001",
			588 => "0001111000101000110100",
			589 => "0011101110111100110000",
			590 => "0000001000000100000100",
			591 => "1111111000100110101101",
			592 => "0010001001001100001100",
			593 => "0000010110010000001000",
			594 => "0011011011101100000100",
			595 => "1111111000100110101101",
			596 => "0000000000100110101101",
			597 => "0000000000100110101101",
			598 => "0011000011010000010000",
			599 => "0000010110010000001000",
			600 => "0000001110100000000100",
			601 => "0000001000100110101101",
			602 => "1111111000100110101101",
			603 => "0001011101001000000100",
			604 => "0000001000100110101101",
			605 => "0000001000100110101101",
			606 => "0001011001011000001000",
			607 => "0010110011010000000100",
			608 => "0000000000100110101101",
			609 => "1111111000100110101101",
			610 => "0011010111011100000100",
			611 => "0000000000100110101101",
			612 => "0000001000100110101101",
			613 => "1111111000100110101101",
			614 => "0011001110011000001000",
			615 => "0000000110111100000100",
			616 => "0000001000100110101101",
			617 => "1111111000100110101101",
			618 => "1111111000100110101101",
			619 => "0000001011011101001000",
			620 => "0010000101011100010100",
			621 => "0000001011111000000100",
			622 => "0000000000101010100001",
			623 => "0000010000011000001100",
			624 => "0010111010100100001000",
			625 => "0010101111111100000100",
			626 => "0000000000101010100001",
			627 => "0000000000101010100001",
			628 => "0000000000101010100001",
			629 => "0000000000101010100001",
			630 => "0001111000000000011100",
			631 => "0011000011010000001000",
			632 => "0001000110001100000100",
			633 => "0000000000101010100001",
			634 => "0000001000101010100001",
			635 => "0000010001100100001100",
			636 => "0001001100101100001000",
			637 => "0010011001000100000100",
			638 => "0000000000101010100001",
			639 => "1111111000101010100001",
			640 => "0000000000101010100001",
			641 => "0011101001011000000100",
			642 => "0000000000101010100001",
			643 => "0000000000101010100001",
			644 => "0011010101011100010000",
			645 => "0000010001110000001000",
			646 => "0011001001001000000100",
			647 => "0000000000101010100001",
			648 => "0000000000101010100001",
			649 => "0011101010100000000100",
			650 => "0000000000101010100001",
			651 => "0000001000101010100001",
			652 => "0000010011010000000100",
			653 => "0000000000101010100001",
			654 => "0000000000101010100001",
			655 => "0001101101000100010000",
			656 => "0011010111011100000100",
			657 => "1111111000101010100001",
			658 => "0001000011110100001000",
			659 => "0011011100101000000100",
			660 => "0000000000101010100001",
			661 => "0000000000101010100001",
			662 => "0000000000101010100001",
			663 => "0001101111000100001000",
			664 => "0000000010101000000100",
			665 => "0000001000101010100001",
			666 => "0000000000101010100001",
			667 => "0000010000011000001100",
			668 => "0010001001001100000100",
			669 => "0000000000101010100001",
			670 => "0011101110111100000100",
			671 => "0000000000101010100001",
			672 => "0000000000101010100001",
			673 => "0001100010000000000100",
			674 => "1111111000101010100001",
			675 => "0010001111001000001000",
			676 => "0010001111111100000100",
			677 => "0000000000101010100001",
			678 => "0000000000101010100001",
			679 => "0000000000101010100001",
			680 => "0000001100000100101100",
			681 => "0010000011010000000100",
			682 => "0000000000101101110101",
			683 => "0001100100000000100100",
			684 => "0000000111001000011000",
			685 => "0011000101011100010000",
			686 => "0001010110001100001000",
			687 => "0010100110010000000100",
			688 => "0000000000101101110101",
			689 => "0000000000101101110101",
			690 => "0000010001110000000100",
			691 => "0000000000101101110101",
			692 => "0000000000101101110101",
			693 => "0000010011010000000100",
			694 => "0000000000101101110101",
			695 => "0000000000101101110101",
			696 => "0000011000011000001000",
			697 => "0000000011101000000100",
			698 => "0000000000101101110101",
			699 => "0000000000101101110101",
			700 => "0000000000101101110101",
			701 => "0000000000101101110101",
			702 => "0001001110111000101100",
			703 => "0011101010011000010000",
			704 => "0011010111011100000100",
			705 => "0000000000101101110101",
			706 => "0011011100101000001000",
			707 => "0000000110011000000100",
			708 => "0000000000101101110101",
			709 => "0000000000101101110101",
			710 => "0000000000101101110101",
			711 => "0000110011001000001100",
			712 => "0000111111011000000100",
			713 => "0000000000101101110101",
			714 => "0000000001110100000100",
			715 => "0000000000101101110101",
			716 => "0000000000101101110101",
			717 => "0011010110001100001000",
			718 => "0001101110010000000100",
			719 => "0000000000101101110101",
			720 => "0000000000101101110101",
			721 => "0001000000111100000100",
			722 => "0000000000101101110101",
			723 => "0000000000101101110101",
			724 => "0010100001101000001000",
			725 => "0000111110111000000100",
			726 => "0000000000101101110101",
			727 => "0000000000101101110101",
			728 => "0001000010001100000100",
			729 => "0000000000101101110101",
			730 => "0001001111100100000100",
			731 => "0000000000101101110101",
			732 => "0000000000101101110101",
			733 => "0000000100011001001000",
			734 => "0011100101110000111000",
			735 => "0000001100000100100100",
			736 => "0011100001101000011000",
			737 => "0010110110001100001000",
			738 => "0000000001101000000100",
			739 => "0000000000110001011001",
			740 => "0000000000110001011001",
			741 => "0000010111100100001000",
			742 => "0010001111001000000100",
			743 => "0000000000110001011001",
			744 => "0000000000110001011001",
			745 => "0001000101011100000100",
			746 => "0000000000110001011001",
			747 => "0000000000110001011001",
			748 => "0011000101010100001000",
			749 => "0010101001010100000100",
			750 => "0000000000110001011001",
			751 => "0000000000110001011001",
			752 => "0000000000110001011001",
			753 => "0010001111111100001000",
			754 => "0011101010100000000100",
			755 => "0000000000110001011001",
			756 => "0000000000110001011001",
			757 => "0010001001000100000100",
			758 => "0000000000110001011001",
			759 => "0010000000110000000100",
			760 => "0000000000110001011001",
			761 => "0000000000110001011001",
			762 => "0000010110010000001000",
			763 => "0010101001000000000100",
			764 => "0000000000110001011001",
			765 => "0000000000110001011001",
			766 => "0011010101010100000100",
			767 => "0000000000110001011001",
			768 => "0000000000110001011001",
			769 => "0011101111111000000100",
			770 => "0000000000110001011001",
			771 => "0001100011010100010100",
			772 => "0001100000110100001100",
			773 => "0011100000010100001000",
			774 => "0011110011010100000100",
			775 => "0000000000110001011001",
			776 => "0000000000110001011001",
			777 => "0000000000110001011001",
			778 => "0000000011100000000100",
			779 => "0000000000110001011001",
			780 => "0000000000110001011001",
			781 => "0001111101001000010000",
			782 => "0000010110010000001000",
			783 => "0000000011111000000100",
			784 => "0000000000110001011001",
			785 => "0000000000110001011001",
			786 => "0001110110101100000100",
			787 => "0000000000110001011001",
			788 => "0000000000110001011001",
			789 => "0000000000110001011001",
			790 => "0000101000010100111000",
			791 => "0011101010100000101000",
			792 => "0000000011101100011000",
			793 => "0011000101011100010000",
			794 => "0010000011010000000100",
			795 => "0000000000110100110101",
			796 => "0001011001100000000100",
			797 => "0000000000110100110101",
			798 => "0000010001110000000100",
			799 => "0000000000110100110101",
			800 => "0000000000110100110101",
			801 => "0000010011010000000100",
			802 => "0000000000110100110101",
			803 => "0000000000110100110101",
			804 => "0000011000011000001000",
			805 => "0011100010001100000100",
			806 => "0000000000110100110101",
			807 => "0000000000110100110101",
			808 => "0011100001101000000100",
			809 => "0000000000110100110101",
			810 => "0000000000110100110101",
			811 => "0011010101011100001100",
			812 => "0010001111111100001000",
			813 => "0001101111111000000100",
			814 => "0000000000110100110101",
			815 => "0000000000110100110101",
			816 => "0000000000110100110101",
			817 => "0000000000110100110101",
			818 => "0001101101000100000100",
			819 => "0000000000110100110101",
			820 => "0001001000000100011000",
			821 => "0000110011001000001100",
			822 => "0000111111011000000100",
			823 => "0000000000110100110101",
			824 => "0001110110101100000100",
			825 => "0000000000110100110101",
			826 => "0000000000110100110101",
			827 => "0011001010100100001000",
			828 => "0011001110011000000100",
			829 => "0000000000110100110101",
			830 => "0000000000110100110101",
			831 => "0000000000110100110101",
			832 => "0000000010101000000100",
			833 => "0000000000110100110101",
			834 => "0001111101001000001100",
			835 => "0000000000011100000100",
			836 => "0000000000110100110101",
			837 => "0000001001110100000100",
			838 => "0000000000110100110101",
			839 => "0000000000110100110101",
			840 => "0001000010111000000100",
			841 => "0000000000110100110101",
			842 => "0011101110000000000100",
			843 => "0000000000110100110101",
			844 => "0000000000110100110101",
			845 => "0000100111010001001000",
			846 => "0001010011000000010000",
			847 => "0011001110011000001100",
			848 => "0010000011010000000100",
			849 => "1111111000110111111001",
			850 => "0000010111100100000100",
			851 => "0000001000110111111001",
			852 => "0000010000110111111001",
			853 => "1111111000110111111001",
			854 => "0000010110010000011000",
			855 => "0011011010100100010100",
			856 => "0000000001111000001100",
			857 => "0011100010001100001000",
			858 => "0000000111001000000100",
			859 => "0000000000110111111001",
			860 => "1111111000110111111001",
			861 => "0000001000110111111001",
			862 => "0011100010011100000100",
			863 => "1111111000110111111001",
			864 => "0000000000110111111001",
			865 => "0000001000110111111001",
			866 => "0011000110000000011100",
			867 => "0011000011010000001100",
			868 => "0010101100010000001000",
			869 => "0000010011110000000100",
			870 => "0000010000110111111001",
			871 => "0000001000110111111001",
			872 => "0000001000110111111001",
			873 => "0001011001011000001000",
			874 => "0010110111011100000100",
			875 => "0000001000110111111001",
			876 => "1111111000110111111001",
			877 => "0011101111100100000100",
			878 => "0000001000110111111001",
			879 => "0000010000110111111001",
			880 => "1111111000110111111001",
			881 => "0011101110111100011000",
			882 => "0011110100001100001000",
			883 => "0000001101001100000100",
			884 => "0000000000110111111001",
			885 => "1111111000110111111001",
			886 => "0001111000101000001100",
			887 => "0010001111111100001000",
			888 => "0011000101010100000100",
			889 => "1111111000110111111001",
			890 => "0000001000110111111001",
			891 => "0000001000110111111001",
			892 => "1111111000110111111001",
			893 => "1111111000110111111001",
			894 => "0001110001010000110000",
			895 => "0001100100010000101100",
			896 => "0000001000000100000100",
			897 => "1111111000111001011101",
			898 => "0010001001001100010000",
			899 => "0010000011010000000100",
			900 => "1111111000111001011101",
			901 => "0000000001111000001000",
			902 => "0011000011010000000100",
			903 => "0000000000111001011101",
			904 => "0000001000111001011101",
			905 => "1111111000111001011101",
			906 => "0011001010100100001100",
			907 => "0010001111111100000100",
			908 => "0000001000111001011101",
			909 => "0011011011101100000100",
			910 => "0000001000111001011101",
			911 => "0000001000111001011101",
			912 => "0001011000000100000100",
			913 => "1111111000111001011101",
			914 => "0011101101000100000100",
			915 => "0000000000111001011101",
			916 => "0000001000111001011101",
			917 => "1111111000111001011101",
			918 => "1111111000111001011101",
			919 => "0001100100010000110100",
			920 => "0010000011010000000100",
			921 => "1111111000111011001001",
			922 => "0001000111100100001000",
			923 => "0000101000000100000100",
			924 => "0000000000111011001001",
			925 => "1111111000111011001001",
			926 => "0011001010100100001000",
			927 => "0010001111111100000100",
			928 => "0000000000111011001001",
			929 => "0000001000111011001001",
			930 => "0001011001011000010000",
			931 => "0010010110000000001000",
			932 => "0000010111100100000100",
			933 => "1111111000111011001001",
			934 => "0000000000111011001001",
			935 => "0001111100010000000100",
			936 => "0000000000111011001001",
			937 => "1111111000111011001001",
			938 => "0000010111110000001000",
			939 => "0001110110101100000100",
			940 => "0000001000111011001001",
			941 => "0000000000111011001001",
			942 => "0011011110011000000100",
			943 => "0000000000111011001001",
			944 => "0000000000111011001001",
			945 => "1111111000111011001001",
			946 => "0000101010111101000100",
			947 => "0011100100000000111000",
			948 => "0010011010000100100000",
			949 => "0011111010110100011100",
			950 => "0000000111001000010000",
			951 => "0001010110001100001000",
			952 => "0001110111011100000100",
			953 => "0000000000111111010101",
			954 => "0000000000111111010101",
			955 => "0010010110000000000100",
			956 => "0000000000111111010101",
			957 => "0000000000111111010101",
			958 => "0011011010100100001000",
			959 => "0000010000011000000100",
			960 => "0000000000111111010101",
			961 => "0000000000111111010101",
			962 => "0000000000111111010101",
			963 => "0000000000111111010101",
			964 => "0010001001000100001000",
			965 => "0010011111011000000100",
			966 => "0000000000111111010101",
			967 => "0000000000111111010101",
			968 => "0001111100010000001000",
			969 => "0000000110100000000100",
			970 => "0000000000111111010101",
			971 => "0000000000111111010101",
			972 => "0010001010000100000100",
			973 => "0000000000111111010101",
			974 => "0000000000111111010101",
			975 => "0011010101010100001000",
			976 => "0010010110000000000100",
			977 => "0000000000111111010101",
			978 => "0000000000111111010101",
			979 => "0000000000111111010101",
			980 => "0011101010011000011000",
			981 => "0011011010100100001000",
			982 => "0010010011000000000100",
			983 => "0000000000111111010101",
			984 => "0000000000111111010101",
			985 => "0001001000000100000100",
			986 => "0000000000111111010101",
			987 => "0011010101010100000100",
			988 => "0000000000111111010101",
			989 => "0011101001111100000100",
			990 => "0000000000111111010101",
			991 => "0000000000111111010101",
			992 => "0001100011010100010000",
			993 => "0011110101110100001000",
			994 => "0011110010001000000100",
			995 => "0000000000111111010101",
			996 => "0000000000111111010101",
			997 => "0011001001001000000100",
			998 => "0000000000111111010101",
			999 => "0000000000111111010101",
			1000 => "0001111101001000010000",
			1001 => "0001011100010000000100",
			1002 => "0000000000111111010101",
			1003 => "0011011011101100001000",
			1004 => "0011010110001100000100",
			1005 => "0000000000111111010101",
			1006 => "0000000000111111010101",
			1007 => "0000000000111111010101",
			1008 => "0011001110011000001000",
			1009 => "0001000101011100000100",
			1010 => "0000000000111111010101",
			1011 => "0000000000111111010101",
			1012 => "0000000000111111010101",
			1013 => "0001100100010001000100",
			1014 => "0011010101011100111000",
			1015 => "0001000010111000110000",
			1016 => "0000011000011000011000",
			1017 => "0001001100010000001100",
			1018 => "0011000110110100000100",
			1019 => "0000001001000001100001",
			1020 => "0010101100010000000100",
			1021 => "0000000001000001100001",
			1022 => "1111111001000001100001",
			1023 => "0001111000000100000100",
			1024 => "1111111001000001100001",
			1025 => "0000110011000100000100",
			1026 => "0000000001000001100001",
			1027 => "0000000001000001100001",
			1028 => "0000000100011000010000",
			1029 => "0011000101011100001000",
			1030 => "0010101110011000000100",
			1031 => "0000000001000001100001",
			1032 => "0000001001000001100001",
			1033 => "0011010111011100000100",
			1034 => "0000000001000001100001",
			1035 => "0000000001000001100001",
			1036 => "0001100010000000000100",
			1037 => "1111111001000001100001",
			1038 => "0000000001000001100001",
			1039 => "0001111000101000000100",
			1040 => "0000001001000001100001",
			1041 => "1111111001000001100001",
			1042 => "0001111000111000001000",
			1043 => "0001101100001100000100",
			1044 => "0000000001000001100001",
			1045 => "0000001001000001100001",
			1046 => "1111111001000001100001",
			1047 => "1111111001000001100001",
			1048 => "0010001001001100010000",
			1049 => "0001111100000000001100",
			1050 => "0010000011010000000100",
			1051 => "0000000001000100010101",
			1052 => "0011000011010000000100",
			1053 => "0000000001000100010101",
			1054 => "0000000001000100010101",
			1055 => "1111111001000100010101",
			1056 => "0001000010111001000100",
			1057 => "0000111110111000110100",
			1058 => "0001001100101100100000",
			1059 => "0010110111011100010000",
			1060 => "0000011000011000001000",
			1061 => "0000000111000100000100",
			1062 => "0000000001000100010101",
			1063 => "0000000001000100010101",
			1064 => "0001000011000000000100",
			1065 => "0000000001000100010101",
			1066 => "0000001001000100010101",
			1067 => "0001001111101000001000",
			1068 => "0010000101011100000100",
			1069 => "0000000001000100010101",
			1070 => "1111111001000100010101",
			1071 => "0000111011000000000100",
			1072 => "0000000001000100010101",
			1073 => "0000000001000100010101",
			1074 => "0010010110000000000100",
			1075 => "0000000001000100010101",
			1076 => "0001010001111100001000",
			1077 => "0000000000001100000100",
			1078 => "0000001001000100010101",
			1079 => "0000000001000100010101",
			1080 => "0000110001001000000100",
			1081 => "0000000001000100010101",
			1082 => "0000000001000100010101",
			1083 => "0001001110111000001000",
			1084 => "0011001001001000000100",
			1085 => "1111111001000100010101",
			1086 => "0000000001000100010101",
			1087 => "0000001100111100000100",
			1088 => "0000000001000100010101",
			1089 => "0000000001000100010101",
			1090 => "0001111000101000000100",
			1091 => "0000001001000100010101",
			1092 => "0000000001000100010101",
			1093 => "0000000111001000011000",
			1094 => "0001010110001100001000",
			1095 => "0001110101010100000100",
			1096 => "0000000001000111100001",
			1097 => "0000000001000111100001",
			1098 => "0011000101011100001000",
			1099 => "0010001001001100000100",
			1100 => "0000000001000111100001",
			1101 => "0000000001000111100001",
			1102 => "0000010011010000000100",
			1103 => "0000000001000111100001",
			1104 => "0000000001000111100001",
			1105 => "0011100010001100001000",
			1106 => "0010001111001000000100",
			1107 => "0000000001000111100001",
			1108 => "0000000001000111100001",
			1109 => "0001010011000100101000",
			1110 => "0000011000011000001100",
			1111 => "0001010101111000001000",
			1112 => "0001010011000000000100",
			1113 => "0000000001000111100001",
			1114 => "0000000001000111100001",
			1115 => "1111111001000111100001",
			1116 => "0011010011010000001100",
			1117 => "0001010101111000000100",
			1118 => "0000000001000111100001",
			1119 => "0010101001010100000100",
			1120 => "0000000001000111100001",
			1121 => "0000000001000111100001",
			1122 => "0000001011101000001000",
			1123 => "0011111010011000000100",
			1124 => "0000000001000111100001",
			1125 => "0000000001000111100001",
			1126 => "0000100111000100000100",
			1127 => "0000000001000111100001",
			1128 => "0000000001000111100001",
			1129 => "0000001100000100000100",
			1130 => "0000000001000111100001",
			1131 => "0001100000110100010000",
			1132 => "0000000010111100001000",
			1133 => "0001101010011000000100",
			1134 => "0000000001000111100001",
			1135 => "0000000001000111100001",
			1136 => "0010001111001000000100",
			1137 => "0000000001000111100001",
			1138 => "0000000001000111100001",
			1139 => "0010001111001000001000",
			1140 => "0011001001001000000100",
			1141 => "0000000001000111100001",
			1142 => "0000000001000111100001",
			1143 => "0000000001000111100001",
			1144 => "0000000000100100111100",
			1145 => "0000001000000100000100",
			1146 => "1111111001001001111101",
			1147 => "0000011001100100000100",
			1148 => "1111111001001001111101",
			1149 => "0010110101011100011100",
			1150 => "0000011000011000010000",
			1151 => "0011101001101100001000",
			1152 => "0011001110011000000100",
			1153 => "0000001001001001111101",
			1154 => "0000000001001001111101",
			1155 => "0011011110011000000100",
			1156 => "0000000001001001111101",
			1157 => "0000001001001001111101",
			1158 => "0000000111101000001000",
			1159 => "0010101110011000000100",
			1160 => "0000001001001001111101",
			1161 => "0000001001001001111101",
			1162 => "0000001001001001111101",
			1163 => "0001001111101000001100",
			1164 => "0000010011010000001000",
			1165 => "0001001010000100000100",
			1166 => "1111111001001001111101",
			1167 => "1111111001001001111101",
			1168 => "0000000001001001111101",
			1169 => "0010100001111100001000",
			1170 => "0000111001000000000100",
			1171 => "0000001001001001111101",
			1172 => "0000001001001001111101",
			1173 => "1111111001001001111101",
			1174 => "0011101110111100010000",
			1175 => "0001100000110100000100",
			1176 => "1111111001001001111101",
			1177 => "0000010110010000000100",
			1178 => "0000001001001001111101",
			1179 => "0011111111010100000100",
			1180 => "0000000001001001111101",
			1181 => "1111111001001001111101",
			1182 => "1111111001001001111101",
			1183 => "0001100100010000111100",
			1184 => "0010000011010000000100",
			1185 => "1111111001001011111001",
			1186 => "0011010101011100101100",
			1187 => "0010001001000100010100",
			1188 => "0010101100110100010000",
			1189 => "0010101010011100001000",
			1190 => "0010011010000100000100",
			1191 => "0000000001001011111001",
			1192 => "0000000001001011111001",
			1193 => "0001011010100000000100",
			1194 => "0000001001001011111001",
			1195 => "0000000001001011111001",
			1196 => "1111111001001011111001",
			1197 => "0000010111100100001100",
			1198 => "0001111000000000000100",
			1199 => "0000000001001011111001",
			1200 => "0010011111011000000100",
			1201 => "0000001001001011111001",
			1202 => "0000000001001011111001",
			1203 => "0001101111000100001000",
			1204 => "0011011010100100000100",
			1205 => "0000000001001011111001",
			1206 => "0000001001001011111001",
			1207 => "0000000001001011111001",
			1208 => "0001111100010000001000",
			1209 => "0011000101101100000100",
			1210 => "0000001001001011111001",
			1211 => "0000000001001011111001",
			1212 => "1111111001001011111001",
			1213 => "1111111001001011111001",
			1214 => "0001101111010101100100",
			1215 => "0011011110011000101100",
			1216 => "0000111011000000011100",
			1217 => "0000110100101100011000",
			1218 => "0010001111111100001100",
			1219 => "0011000110110100000100",
			1220 => "0000000001001111011101",
			1221 => "0010010101101100000100",
			1222 => "1111111001001111011101",
			1223 => "0000000001001111011101",
			1224 => "0011000011010000000100",
			1225 => "0000001001001111011101",
			1226 => "0001111000000000000100",
			1227 => "0000000001001111011101",
			1228 => "0000000001001111011101",
			1229 => "0000001001001111011101",
			1230 => "0010010011000000001100",
			1231 => "0001000001011000000100",
			1232 => "1111111001001111011101",
			1233 => "0001000011110100000100",
			1234 => "0000000001001111011101",
			1235 => "0000000001001111011101",
			1236 => "0000000001001111011101",
			1237 => "0010110101011100011000",
			1238 => "0001000001011000010100",
			1239 => "0000101100111000001100",
			1240 => "0001001101001000001000",
			1241 => "0011000011010000000100",
			1242 => "0000001001001111011101",
			1243 => "0000000001001111011101",
			1244 => "0000001001001111011101",
			1245 => "0000001011000100000100",
			1246 => "0000000001001111011101",
			1247 => "0000000001001111011101",
			1248 => "0000001001001111011101",
			1249 => "0000110000111100010100",
			1250 => "0010001001000100000100",
			1251 => "1111111001001111011101",
			1252 => "0010001111001000001000",
			1253 => "0011010111011100000100",
			1254 => "0000000001001111011101",
			1255 => "0000000001001111011101",
			1256 => "0000010011010000000100",
			1257 => "0000000001001111011101",
			1258 => "0000000001001111011101",
			1259 => "0010100000111000000100",
			1260 => "0000000001001111011101",
			1261 => "0000001100111100000100",
			1262 => "0000000001001111011101",
			1263 => "0000000001001111011101",
			1264 => "0000010111110000001100",
			1265 => "0010101011000000000100",
			1266 => "0000000001001111011101",
			1267 => "0010100000111100000100",
			1268 => "0000000001001111011101",
			1269 => "0000000001001111011101",
			1270 => "1111111001001111011101",
			1271 => "0001100100010001010100",
			1272 => "0011010101011101001000",
			1273 => "0000011000011000101100",
			1274 => "0011101111100100011000",
			1275 => "0000100100011100001100",
			1276 => "0011111010110100001000",
			1277 => "0010110110001100000100",
			1278 => "0000001001010010001001",
			1279 => "0000000001010010001001",
			1280 => "0000001001010010001001",
			1281 => "0000010111100100001000",
			1282 => "0001101111111000000100",
			1283 => "0000000001010010001001",
			1284 => "1111111001010010001001",
			1285 => "1111111001010010001001",
			1286 => "0001010011000100001000",
			1287 => "0000001101010000000100",
			1288 => "0000000001010010001001",
			1289 => "1111111001010010001001",
			1290 => "0000000100011000000100",
			1291 => "0000001001010010001001",
			1292 => "0011101111111000000100",
			1293 => "1111111001010010001001",
			1294 => "0000000001010010001001",
			1295 => "0000101000110100010000",
			1296 => "0011001100101000001000",
			1297 => "0010101110011000000100",
			1298 => "0000000001010010001001",
			1299 => "0000001001010010001001",
			1300 => "0001010101011100000100",
			1301 => "1111111001010010001001",
			1302 => "0000000001010010001001",
			1303 => "0011100010011100000100",
			1304 => "1111111001010010001001",
			1305 => "0011010011010000000100",
			1306 => "0000001001010010001001",
			1307 => "0000000001010010001001",
			1308 => "0001111100010000001000",
			1309 => "0011000101101100000100",
			1310 => "0000001001010010001001",
			1311 => "1111111001010010001001",
			1312 => "1111111001010010001001",
			1313 => "1111111001010010001001",
			1314 => "0010001001001100010000",
			1315 => "0000001001000000000100",
			1316 => "0000000001010101101101",
			1317 => "0000111100101100001000",
			1318 => "0000111111101000000100",
			1319 => "0000000001010101101101",
			1320 => "0000000001010101101101",
			1321 => "0000000001010101101101",
			1322 => "0010110101011101000100",
			1323 => "0011111110100000110000",
			1324 => "0001111000000000011000",
			1325 => "0000001110100000001100",
			1326 => "0001000111100100000100",
			1327 => "0000000001010101101101",
			1328 => "0010010110000000000100",
			1329 => "0000000001010101101101",
			1330 => "0000000001010101101101",
			1331 => "0011011010100100001000",
			1332 => "0000100100011100000100",
			1333 => "0000000001010101101101",
			1334 => "0000000001010101101101",
			1335 => "0000000001010101101101",
			1336 => "0010001111111100001100",
			1337 => "0011101011110000001000",
			1338 => "0000000101100000000100",
			1339 => "0000000001010101101101",
			1340 => "0000000001010101101101",
			1341 => "0000000001010101101101",
			1342 => "0000011001100000001000",
			1343 => "0001101010100000000100",
			1344 => "0000000001010101101101",
			1345 => "0000000001010101101101",
			1346 => "0000000001010101101101",
			1347 => "0001010011000100001100",
			1348 => "0011001110011000001000",
			1349 => "0000000010101100000100",
			1350 => "0000000001010101101101",
			1351 => "0000000001010101101101",
			1352 => "0000000001010101101101",
			1353 => "0011000101010100000100",
			1354 => "0000000001010101101101",
			1355 => "0000000001010101101101",
			1356 => "0011001100101000001000",
			1357 => "0001100010001100000100",
			1358 => "0000000001010101101101",
			1359 => "0000000001010101101101",
			1360 => "0010011101101000000100",
			1361 => "0000000001010101101101",
			1362 => "0001111100010000000100",
			1363 => "0000000001010101101101",
			1364 => "0001110110101100001000",
			1365 => "0011101110010100000100",
			1366 => "0000000001010101101101",
			1367 => "0000000001010101101101",
			1368 => "0001000001111100000100",
			1369 => "0000000001010101101101",
			1370 => "0000000001010101101101",
			1371 => "0000001100000100110000",
			1372 => "0010000011010000000100",
			1373 => "0000000001011001100001",
			1374 => "0001000110011100101000",
			1375 => "0011000011010000001100",
			1376 => "0000010110010000001000",
			1377 => "0000001010011000000100",
			1378 => "0000000001011001100001",
			1379 => "0000000001011001100001",
			1380 => "0000000001011001100001",
			1381 => "0000011000011000001100",
			1382 => "0000000010110100001000",
			1383 => "0001111000000000000100",
			1384 => "0000000001011001100001",
			1385 => "0000000001011001100001",
			1386 => "0000000001011001100001",
			1387 => "0001111100010000001000",
			1388 => "0011101001011000000100",
			1389 => "0000000001011001100001",
			1390 => "0000000001011001100001",
			1391 => "0010001111001000000100",
			1392 => "0000000001011001100001",
			1393 => "0000000001011001100001",
			1394 => "0000000001011001100001",
			1395 => "0011100101110000011000",
			1396 => "0000010111110000001100",
			1397 => "0001001011111000001000",
			1398 => "0001000011000000000100",
			1399 => "0000000001011001100001",
			1400 => "0000000001011001100001",
			1401 => "0000000001011001100001",
			1402 => "0011010111011100000100",
			1403 => "1111111001011001100001",
			1404 => "0011011100101000000100",
			1405 => "0000000001011001100001",
			1406 => "0000000001011001100001",
			1407 => "0000000010010000001100",
			1408 => "0000010110010000000100",
			1409 => "0000000001011001100001",
			1410 => "0000110001001000000100",
			1411 => "0000001001011001100001",
			1412 => "0000000001011001100001",
			1413 => "0001001110001100011100",
			1414 => "0000011000011000001100",
			1415 => "0011010111011100001000",
			1416 => "0001100110110000000100",
			1417 => "0000000001011001100001",
			1418 => "0000000001011001100001",
			1419 => "0000000001011001100001",
			1420 => "0010101101001000001000",
			1421 => "0001011000111000000100",
			1422 => "0000000001011001100001",
			1423 => "0000000001011001100001",
			1424 => "0001101111000100000100",
			1425 => "0000000001011001100001",
			1426 => "0000000001011001100001",
			1427 => "0000110001101000001000",
			1428 => "0010111100101000000100",
			1429 => "0000000001011001100001",
			1430 => "0000000001011001100001",
			1431 => "0000000001011001100001",
			1432 => "0001100100010001000100",
			1433 => "0010010011001001000000",
			1434 => "0011101010011000100100",
			1435 => "0000101110000100010100",
			1436 => "0000011001100100000100",
			1437 => "1111111001011011101101",
			1438 => "0011001110011000001000",
			1439 => "0011010110110100000100",
			1440 => "0000000001011011101101",
			1441 => "0000001001011011101101",
			1442 => "0001011000000100000100",
			1443 => "1111111001011011101101",
			1444 => "0000000001011011101101",
			1445 => "0010001111001000001100",
			1446 => "0001111101001000001000",
			1447 => "0010101000101000000100",
			1448 => "1111111001011011101101",
			1449 => "1111111001011011101101",
			1450 => "0000000001011011101101",
			1451 => "0000000001011011101101",
			1452 => "0001100011010100001000",
			1453 => "0010101100001100000100",
			1454 => "0000001001011011101101",
			1455 => "0000000001011011101101",
			1456 => "0011110100101000001000",
			1457 => "0001001001000100000100",
			1458 => "0000000001011011101101",
			1459 => "1111111001011011101101",
			1460 => "0010011001001000000100",
			1461 => "1111111001011011101101",
			1462 => "0000010110010000000100",
			1463 => "0000001001011011101101",
			1464 => "0000000001011011101101",
			1465 => "1111111001011011101101",
			1466 => "1111111001011011101101",
			1467 => "0010001001001100001000",
			1468 => "0000001001000000000100",
			1469 => "0000000001011111000001",
			1470 => "0000000001011111000001",
			1471 => "0010110101011101000100",
			1472 => "0011111110100000110000",
			1473 => "0001111000000000011000",
			1474 => "0000001110100000001100",
			1475 => "0001000111100100000100",
			1476 => "0000000001011111000001",
			1477 => "0010010110000000000100",
			1478 => "0000000001011111000001",
			1479 => "0000000001011111000001",
			1480 => "0011011010100100001000",
			1481 => "0000100100011100000100",
			1482 => "0000000001011111000001",
			1483 => "0000000001011111000001",
			1484 => "0000000001011111000001",
			1485 => "0010001111111100001100",
			1486 => "0011101011110000001000",
			1487 => "0000001101010000000100",
			1488 => "0000000001011111000001",
			1489 => "0000000001011111000001",
			1490 => "0000000001011111000001",
			1491 => "0000011001100000001000",
			1492 => "0001101010100000000100",
			1493 => "0000000001011111000001",
			1494 => "0000000001011111000001",
			1495 => "0000000001011111000001",
			1496 => "0001010011000100001100",
			1497 => "0011001110011000001000",
			1498 => "0000000010101100000100",
			1499 => "0000000001011111000001",
			1500 => "0000000001011111000001",
			1501 => "0000000001011111000001",
			1502 => "0011000101010100000100",
			1503 => "0000000001011111000001",
			1504 => "0000000001011111000001",
			1505 => "0011001100101000001000",
			1506 => "0001100010001100000100",
			1507 => "0000000001011111000001",
			1508 => "0000000001011111000001",
			1509 => "0010011101101000000100",
			1510 => "0000000001011111000001",
			1511 => "0001111100010000000100",
			1512 => "0000000001011111000001",
			1513 => "0001110110101100001000",
			1514 => "0011101110010100000100",
			1515 => "0000000001011111000001",
			1516 => "0000000001011111000001",
			1517 => "0001000001111100000100",
			1518 => "0000000001011111000001",
			1519 => "0000000001011111000001",
			1520 => "0011101110111101001000",
			1521 => "0011000110000001000100",
			1522 => "0010001001001100010000",
			1523 => "0010010110000000001000",
			1524 => "0001000111100100000100",
			1525 => "0000000001100001010101",
			1526 => "1111111001100001010101",
			1527 => "0010110111011100000100",
			1528 => "0000001001100001010101",
			1529 => "1111111001100001010101",
			1530 => "0011000011010000010100",
			1531 => "0000001110100000001100",
			1532 => "0001011011101100000100",
			1533 => "0000000001100001010101",
			1534 => "0000001001111100000100",
			1535 => "0000001001100001010101",
			1536 => "0000001001100001010101",
			1537 => "0000010110010000000100",
			1538 => "1111111001100001010101",
			1539 => "0000000001100001010101",
			1540 => "0001011001011000010000",
			1541 => "0010110011010000001000",
			1542 => "0000011000011000000100",
			1543 => "1111111001100001010101",
			1544 => "0000001001100001010101",
			1545 => "0010011001000100000100",
			1546 => "0000000001100001010101",
			1547 => "1111111001100001010101",
			1548 => "0011101111100100001000",
			1549 => "0000000100110000000100",
			1550 => "0000001001100001010101",
			1551 => "0000000001100001010101",
			1552 => "0000000111000000000100",
			1553 => "0000001001100001010101",
			1554 => "0000000001100001010101",
			1555 => "1111111001100001010101",
			1556 => "1111111001100001010101",
			1557 => "0001100100010001100000",
			1558 => "0001111000000000100100",
			1559 => "0000110011000100100000",
			1560 => "0011001100101000011100",
			1561 => "0011000101010100010000",
			1562 => "0000111101001000001000",
			1563 => "0001010110101100000100",
			1564 => "0000000001100100011001",
			1565 => "0000001001100100011001",
			1566 => "0000111011111000000100",
			1567 => "1111111001100100011001",
			1568 => "0000000001100100011001",
			1569 => "0011100001101000001000",
			1570 => "0011011010100100000100",
			1571 => "0000000001100100011001",
			1572 => "0000000001100100011001",
			1573 => "0000001001100100011001",
			1574 => "1111111001100100011001",
			1575 => "1111111001100100011001",
			1576 => "0001010001101000100000",
			1577 => "0010010110000000001100",
			1578 => "0001110110101100001000",
			1579 => "0001111100010000000100",
			1580 => "0000000001100100011001",
			1581 => "0000000001100100011001",
			1582 => "0000001001100100011001",
			1583 => "0000000010010000001100",
			1584 => "0001001100000000001000",
			1585 => "0001111001010100000100",
			1586 => "1111111001100100011001",
			1587 => "0000000001100100011001",
			1588 => "0000000001100100011001",
			1589 => "0001111100110000000100",
			1590 => "0000000001100100011001",
			1591 => "1111111001100100011001",
			1592 => "0010011010000100001000",
			1593 => "0000011001100100000100",
			1594 => "1111111001100100011001",
			1595 => "0000001001100100011001",
			1596 => "0010010011000000001000",
			1597 => "0011001100101000000100",
			1598 => "0000000001100100011001",
			1599 => "1111111001100100011001",
			1600 => "0000100101000100001000",
			1601 => "0010100001101000000100",
			1602 => "0000001001100100011001",
			1603 => "0000000001100100011001",
			1604 => "1111111001100100011001",
			1605 => "1111111001100100011001",
			1606 => "0011100010001001010000",
			1607 => "0010010011001001001100",
			1608 => "0011101010011000110000",
			1609 => "0000101110000100100000",
			1610 => "0000011000011000010000",
			1611 => "0011101111100100001000",
			1612 => "0000000000001100000100",
			1613 => "0000000001100110111101",
			1614 => "1111111001100110111101",
			1615 => "0000010110010000000100",
			1616 => "0000000001100110111101",
			1617 => "0000001001100110111101",
			1618 => "0000100100111000001000",
			1619 => "0001011011101100000100",
			1620 => "0000000001100110111101",
			1621 => "0000001001100110111101",
			1622 => "0001001111011000000100",
			1623 => "1111111001100110111101",
			1624 => "0000000001100110111101",
			1625 => "0010001111001000001100",
			1626 => "0001111101001000001000",
			1627 => "0010101000101000000100",
			1628 => "1111111001100110111101",
			1629 => "1111111001100110111101",
			1630 => "0000000001100110111101",
			1631 => "0000000001100110111101",
			1632 => "0001100011010100001000",
			1633 => "0010101100001100000100",
			1634 => "0000001001100110111101",
			1635 => "0000000001100110111101",
			1636 => "0000000111110100001100",
			1637 => "0010011001001000000100",
			1638 => "1111111001100110111101",
			1639 => "0011110100101000000100",
			1640 => "1111111001100110111101",
			1641 => "0000000001100110111101",
			1642 => "0000111100010000000100",
			1643 => "1111111001100110111101",
			1644 => "0000001001100110111101",
			1645 => "1111111001100110111101",
			1646 => "1111111001100110111101",
			1647 => "0001000010111010000000",
			1648 => "0000001100000100110000",
			1649 => "0001100100000000100100",
			1650 => "0000000111001000011100",
			1651 => "0001000111100100001100",
			1652 => "0000101000000100001000",
			1653 => "0010101001100000000100",
			1654 => "0000000001101011001001",
			1655 => "0000000001101011001001",
			1656 => "1111111001101011001001",
			1657 => "0010010110000000001000",
			1658 => "0000010001110000000100",
			1659 => "0000000001101011001001",
			1660 => "0000001001101011001001",
			1661 => "0000011110011000000100",
			1662 => "1111111001101011001001",
			1663 => "0000000001101011001001",
			1664 => "0011000101010100000100",
			1665 => "1111111001101011001001",
			1666 => "0000000001101011001001",
			1667 => "0000110011001000000100",
			1668 => "0000000001101011001001",
			1669 => "0001101111100100000100",
			1670 => "0000000001101011001001",
			1671 => "0000001001101011001001",
			1672 => "0011101111100100100000",
			1673 => "0010001001000100010100",
			1674 => "0010101001011000001100",
			1675 => "0001101010110100001000",
			1676 => "0010010110000000000100",
			1677 => "0000000001101011001001",
			1678 => "0000001001101011001001",
			1679 => "1111111001101011001001",
			1680 => "0011100101110000000100",
			1681 => "1111111001101011001001",
			1682 => "1111111001101011001001",
			1683 => "0001111000111000000100",
			1684 => "0000000001101011001001",
			1685 => "0010001010000100000100",
			1686 => "0000001001101011001001",
			1687 => "0000000001101011001001",
			1688 => "0001011001011000011000",
			1689 => "0000110011001000001100",
			1690 => "0010010101101100001000",
			1691 => "0000000010000100000100",
			1692 => "0000000001101011001001",
			1693 => "1111111001101011001001",
			1694 => "0000001001101011001001",
			1695 => "0001001001001000001000",
			1696 => "0011110100100000000100",
			1697 => "0000000001101011001001",
			1698 => "0000000001101011001001",
			1699 => "1111111001101011001001",
			1700 => "0000100111010000001100",
			1701 => "0010001111111100000100",
			1702 => "0000000001101011001001",
			1703 => "0000101101010000000100",
			1704 => "0000001001101011001001",
			1705 => "0000000001101011001001",
			1706 => "0011111110100100000100",
			1707 => "1111111001101011001001",
			1708 => "0000010110010000000100",
			1709 => "0000001001101011001001",
			1710 => "0000000001101011001001",
			1711 => "0001111000101000000100",
			1712 => "0000001001101011001001",
			1713 => "1111111001101011001001",
			1714 => "0001100100010001010100",
			1715 => "0011000110000001010000",
			1716 => "0010111110011000010100",
			1717 => "0010000011010000000100",
			1718 => "1111111001101101110111",
			1719 => "0001011000111000001100",
			1720 => "0011001110011000001000",
			1721 => "0010001111111100000100",
			1722 => "0000001001101101110111",
			1723 => "0000001001101101110111",
			1724 => "0000000001101101110111",
			1725 => "0000001001101101110111",
			1726 => "0001000011000000011100",
			1727 => "0010110011010000010000",
			1728 => "0010010101101100001000",
			1729 => "0000100011010100000100",
			1730 => "0000000001101101110111",
			1731 => "1111111001101101110111",
			1732 => "0011011011101100000100",
			1733 => "1111111001101101110111",
			1734 => "0000001001101101110111",
			1735 => "0011000111011100000100",
			1736 => "0000000001101101110111",
			1737 => "0011010101011100000100",
			1738 => "1111111001101101110111",
			1739 => "1111111001101101110111",
			1740 => "0011011010100100010000",
			1741 => "0000111110111000001000",
			1742 => "0001001100101100000100",
			1743 => "0000000001101101110111",
			1744 => "0000000001101101110111",
			1745 => "0011000101011100000100",
			1746 => "1111111001101101110111",
			1747 => "0000000001101101110111",
			1748 => "0010110101011100001000",
			1749 => "0001000110101100000100",
			1750 => "0000000001101101110111",
			1751 => "0000001001101101110111",
			1752 => "0000010111100100000100",
			1753 => "1111111001101101110111",
			1754 => "0000000001101101110111",
			1755 => "1111111001101101110111",
			1756 => "1111111001101101110111",
			1757 => "0001101111010100100100",
			1758 => "0000000000011100011100",
			1759 => "0011111110100000011000",
			1760 => "0001100000110100010000",
			1761 => "0000000000100100001100",
			1762 => "0000011001100100000100",
			1763 => "0000000001101111010001",
			1764 => "0010101100110100000100",
			1765 => "0000000001101111010001",
			1766 => "0000000001101111010001",
			1767 => "1111111001101111010001",
			1768 => "0000001011011000000100",
			1769 => "0000001001101111010001",
			1770 => "0000000001101111010001",
			1771 => "1111111001101111010001",
			1772 => "0001111001010100000100",
			1773 => "0000001001101111010001",
			1774 => "0000000001101111010001",
			1775 => "0000010111110000001000",
			1776 => "0010110011010000000100",
			1777 => "0000000001101111010001",
			1778 => "0000000001101111010001",
			1779 => "1111111001101111010001",
			1780 => "0001000010111000101100",
			1781 => "0000100111000100100000",
			1782 => "0000000111110100011000",
			1783 => "0000011001100100000100",
			1784 => "1111111001110000110101",
			1785 => "0001001100001100010000",
			1786 => "0000000000001100001000",
			1787 => "0011111010110100000100",
			1788 => "0000000001110000110101",
			1789 => "0000000001110000110101",
			1790 => "0001101010011000000100",
			1791 => "1111111001110000110101",
			1792 => "0000000001110000110101",
			1793 => "1111111001110000110101",
			1794 => "0001100100111000000100",
			1795 => "0000001001110000110101",
			1796 => "0000000001110000110101",
			1797 => "0000010000011000001000",
			1798 => "0010111010100100000100",
			1799 => "0000000001110000110101",
			1800 => "0000000001110000110101",
			1801 => "1111111001110000110101",
			1802 => "0000110001101000000100",
			1803 => "0000001001110000110101",
			1804 => "0000000001110000110101",
			1805 => "0000000100011000111000",
			1806 => "0010110101011100100100",
			1807 => "0010001001001100001100",
			1808 => "0000001101010000001000",
			1809 => "0000001001000000000100",
			1810 => "0000000001110011100001",
			1811 => "0000000001110011100001",
			1812 => "0000000001110011100001",
			1813 => "0001000111100100000100",
			1814 => "0000000001110011100001",
			1815 => "0000011001100100000100",
			1816 => "0000000001110011100001",
			1817 => "0000101100111000001000",
			1818 => "0001101101101100000100",
			1819 => "0000000001110011100001",
			1820 => "0000000001110011100001",
			1821 => "0011101001111100000100",
			1822 => "0000000001110011100001",
			1823 => "0000000001110011100001",
			1824 => "0011101111100100010000",
			1825 => "0010011101101000000100",
			1826 => "0000000001110011100001",
			1827 => "0010001001000100000100",
			1828 => "0000000001110011100001",
			1829 => "0010001111001000000100",
			1830 => "0000000001110011100001",
			1831 => "0000000001110011100001",
			1832 => "0000000001110011100001",
			1833 => "0001001110001100011000",
			1834 => "0001111000111000001100",
			1835 => "0001001000000100001000",
			1836 => "0001000101011100000100",
			1837 => "0000000001110011100001",
			1838 => "0000000001110011100001",
			1839 => "0000000001110011100001",
			1840 => "0001100010000000000100",
			1841 => "0000000001110011100001",
			1842 => "0001101111010100000100",
			1843 => "0000000001110011100001",
			1844 => "0000000001110011100001",
			1845 => "0001011010110100000100",
			1846 => "0000000001110011100001",
			1847 => "0000000001110011100001",
			1848 => "0010110101011100110100",
			1849 => "0010001001001100001000",
			1850 => "0000001100001100000100",
			1851 => "0000000001110110000101",
			1852 => "0000000001110110000101",
			1853 => "0000100111000100100100",
			1854 => "0001010110001100001100",
			1855 => "0001000001100100001000",
			1856 => "0001101001000100000100",
			1857 => "0000000001110110000101",
			1858 => "0000000001110110000101",
			1859 => "0000000001110110000101",
			1860 => "0010101100110100010000",
			1861 => "0000011001100100001000",
			1862 => "0001111100010000000100",
			1863 => "0000000001110110000101",
			1864 => "0000000001110110000101",
			1865 => "0001100100010000000100",
			1866 => "0000000001110110000101",
			1867 => "0000000001110110000101",
			1868 => "0000010001110000000100",
			1869 => "0000000001110110000101",
			1870 => "0000000001110110000101",
			1871 => "0000010000011000000100",
			1872 => "0000000001110110000101",
			1873 => "0000000001110110000101",
			1874 => "0011001100101000001000",
			1875 => "0000111001010000000100",
			1876 => "0000000001110110000101",
			1877 => "0000000001110110000101",
			1878 => "0001000001111100010000",
			1879 => "0010011101101000000100",
			1880 => "0000000001110110000101",
			1881 => "0000101000011100000100",
			1882 => "0000000001110110000101",
			1883 => "0011101111110100000100",
			1884 => "0000000001110110000101",
			1885 => "0000000001110110000101",
			1886 => "0000101011010100000100",
			1887 => "0000000001110110000101",
			1888 => "0000000001110110000101",
			1889 => "0000000100110000011100",
			1890 => "0001011001010100001100",
			1891 => "0011001110011000001000",
			1892 => "0010000011010000000100",
			1893 => "0000000001111001001001",
			1894 => "0000000001111001001001",
			1895 => "0000000001111001001001",
			1896 => "0011011011101100000100",
			1897 => "0000000001111001001001",
			1898 => "0011101110010100001000",
			1899 => "0001101110001100000100",
			1900 => "0000000001111001001001",
			1901 => "0000000001111001001001",
			1902 => "0000000001111001001001",
			1903 => "0011101111100100010100",
			1904 => "0000111001000000001100",
			1905 => "0011101010100000001000",
			1906 => "0001101101101100000100",
			1907 => "0000000001111001001001",
			1908 => "0000000001111001001001",
			1909 => "0000000001111001001001",
			1910 => "0010001111111100000100",
			1911 => "0000000001111001001001",
			1912 => "0000000001111001001001",
			1913 => "0000100111010000010000",
			1914 => "0010000101011100001000",
			1915 => "0010110011010000000100",
			1916 => "0000000001111001001001",
			1917 => "0000000001111001001001",
			1918 => "0000111000101000000100",
			1919 => "0000000001111001001001",
			1920 => "0000000001111001001001",
			1921 => "0001111101001000011000",
			1922 => "0001001101101000001000",
			1923 => "0001000101010100000100",
			1924 => "0000000001111001001001",
			1925 => "0000000001111001001001",
			1926 => "0001011100011100001000",
			1927 => "0011001110011000000100",
			1928 => "0000000001111001001001",
			1929 => "0000000001111001001001",
			1930 => "0011000101011100000100",
			1931 => "0000000001111001001001",
			1932 => "0000000001111001001001",
			1933 => "0001000010111000000100",
			1934 => "0000000001111001001001",
			1935 => "0000110001101000000100",
			1936 => "0000000001111001001001",
			1937 => "0000000001111001001001",
			1938 => "0001101111010100111100",
			1939 => "0011101101000100110000",
			1940 => "0000000100110100100100",
			1941 => "0011000110110100000100",
			1942 => "0000000001111011010101",
			1943 => "0011100010001100010000",
			1944 => "0010001001000100001000",
			1945 => "0000011000011000000100",
			1946 => "1111111001111011010101",
			1947 => "0000000001111011010101",
			1948 => "0011001100101000000100",
			1949 => "0000001001111011010101",
			1950 => "0000000001111011010101",
			1951 => "0000000010010000001000",
			1952 => "0001001100000000000100",
			1953 => "0000000001111011010101",
			1954 => "0000000001111011010101",
			1955 => "0001100100100100000100",
			1956 => "1111111001111011010101",
			1957 => "0000000001111011010101",
			1958 => "0011101110000000000100",
			1959 => "1111111001111011010101",
			1960 => "0000101000100100000100",
			1961 => "0000000001111011010101",
			1962 => "0000000001111011010101",
			1963 => "0001010101111000000100",
			1964 => "0000000001111011010101",
			1965 => "0001111111101000000100",
			1966 => "0000001001111011010101",
			1967 => "0000000001111011010101",
			1968 => "0000010111110000001000",
			1969 => "0010110011010000000100",
			1970 => "0000000001111011010101",
			1971 => "0000000001111011010101",
			1972 => "1111111001111011010101",
			1973 => "0001000010111000111000",
			1974 => "0000100111000100101100",
			1975 => "0000000111110100100100",
			1976 => "0000011001100100000100",
			1977 => "1111111001111101010001",
			1978 => "0011001010100100010000",
			1979 => "0010001111111100001000",
			1980 => "0011000110110100000100",
			1981 => "0000000001111101010001",
			1982 => "1111111001111101010001",
			1983 => "0011011011101100000100",
			1984 => "0000000001111101010001",
			1985 => "0000001001111101010001",
			1986 => "0001011100010000001000",
			1987 => "0000000011101000000100",
			1988 => "0000000001111101010001",
			1989 => "1111111001111101010001",
			1990 => "0000111011000000000100",
			1991 => "0000000001111101010001",
			1992 => "0000000001111101010001",
			1993 => "0001100100111000000100",
			1994 => "0000001001111101010001",
			1995 => "0000000001111101010001",
			1996 => "0000010000011000001000",
			1997 => "0010111010100100000100",
			1998 => "0000000001111101010001",
			1999 => "0000000001111101010001",
			2000 => "1111111001111101010001",
			2001 => "0000110001101000000100",
			2002 => "0000001001111101010001",
			2003 => "0000000001111101010001",
			2004 => "0001100100010000111000",
			2005 => "0011001001001000101000",
			2006 => "0000011001100100001000",
			2007 => "0011100000010100000100",
			2008 => "1111111001111111000101",
			2009 => "0000001001111111000101",
			2010 => "0010101100110100011100",
			2011 => "0011001010100100001100",
			2012 => "0010001001001100000100",
			2013 => "0000000001111111000101",
			2014 => "0010001111111100000100",
			2015 => "0000001001111111000101",
			2016 => "0000001001111111000101",
			2017 => "0001001101101000001000",
			2018 => "0000011001100000000100",
			2019 => "1111111001111111000101",
			2020 => "0000000001111111000101",
			2021 => "0000010111110000000100",
			2022 => "0000001001111111000101",
			2023 => "0000000001111111000101",
			2024 => "1111111001111111000101",
			2025 => "0001010010111000000100",
			2026 => "1111111001111111000101",
			2027 => "0000001011000100001000",
			2028 => "0011101011110000000100",
			2029 => "0000000001111111000101",
			2030 => "0000001001111111000101",
			2031 => "1111111001111111000101",
			2032 => "1111111001111111000101",
			2033 => "0001110001010000101100",
			2034 => "0001100100010000101000",
			2035 => "0000001000000100000100",
			2036 => "1111111010000000100001",
			2037 => "0010001001001100001100",
			2038 => "0001101100000000000100",
			2039 => "0000000010000000100001",
			2040 => "0011011011101100000100",
			2041 => "1111111010000000100001",
			2042 => "0000000010000000100001",
			2043 => "0011001010100100001100",
			2044 => "0000010110010000000100",
			2045 => "0000001010000000100001",
			2046 => "0000111101101000000100",
			2047 => "0000001010000000100001",
			2048 => "0000001010000000100001",
			2049 => "0001011000000100000100",
			2050 => "1111111010000000100001",
			2051 => "0011101110000000000100",
			2052 => "0000000010000000100001",
			2053 => "0000001010000000100001",
			2054 => "1111111010000000100001",
			2055 => "1111111010000000100001",
			2056 => "0000101010111101000000",
			2057 => "0001101111100100110000",
			2058 => "0011011010100100011000",
			2059 => "0010110110001100001000",
			2060 => "0000001010100000000100",
			2061 => "0000000010000100000101",
			2062 => "0000000010000100000101",
			2063 => "0010110101010100001000",
			2064 => "0000010001100100000100",
			2065 => "0000000010000100000101",
			2066 => "0000000010000100000101",
			2067 => "0010110101011100000100",
			2068 => "0000000010000100000101",
			2069 => "0000000010000100000101",
			2070 => "0010001111111100001000",
			2071 => "0001111100000000000100",
			2072 => "0000000010000100000101",
			2073 => "0000000010000100000101",
			2074 => "0010111100101000001100",
			2075 => "0001001100101000001000",
			2076 => "0000001011000000000100",
			2077 => "0000000010000100000101",
			2078 => "0000000010000100000101",
			2079 => "0000000010000100000101",
			2080 => "0000000010000100000101",
			2081 => "0011111001110000001100",
			2082 => "0011001001001000001000",
			2083 => "0001001100000000000100",
			2084 => "0000000010000100000101",
			2085 => "0000000010000100000101",
			2086 => "0000000010000100000101",
			2087 => "0000000010000100000101",
			2088 => "0001001000000100001100",
			2089 => "0001000101010100001000",
			2090 => "0011110110110000000100",
			2091 => "0000000010000100000101",
			2092 => "0000000010000100000101",
			2093 => "0000000010000100000101",
			2094 => "0001101101000100010000",
			2095 => "0011101011110000001000",
			2096 => "0011010111011100000100",
			2097 => "0000000010000100000101",
			2098 => "0000000010000100000101",
			2099 => "0011100000100000000100",
			2100 => "0000000010000100000101",
			2101 => "0000000010000100000101",
			2102 => "0000000100111100000100",
			2103 => "0000000010000100000101",
			2104 => "0001111101001000001000",
			2105 => "0000100111000100000100",
			2106 => "0000000010000100000101",
			2107 => "0000000010000100000101",
			2108 => "0001011001111100000100",
			2109 => "0000000010000100000101",
			2110 => "0000110001101000000100",
			2111 => "0000000010000100000101",
			2112 => "0000000010000100000101",
			2113 => "0000000100011001001100",
			2114 => "0011101001101100110000",
			2115 => "0000000111001000100000",
			2116 => "0010010110000000010100",
			2117 => "0001010110001100001100",
			2118 => "0001000000011000000100",
			2119 => "0000000010000111111001",
			2120 => "0001001000011000000100",
			2121 => "0000000010000111111001",
			2122 => "0000000010000111111001",
			2123 => "0010001001001100000100",
			2124 => "0000000010000111111001",
			2125 => "0000000010000111111001",
			2126 => "0000011110011000001000",
			2127 => "0011011011101100000100",
			2128 => "0000000010000111111001",
			2129 => "0000000010000111111001",
			2130 => "0000000010000111111001",
			2131 => "0000011000011000001000",
			2132 => "0010000101011100000100",
			2133 => "0000000010000111111001",
			2134 => "0000000010000111111001",
			2135 => "0010001010000100000100",
			2136 => "0000000010000111111001",
			2137 => "0000000010000111111001",
			2138 => "0010001111011000011000",
			2139 => "0000010001110000001000",
			2140 => "0000000001111000000100",
			2141 => "0000000010000111111001",
			2142 => "0000000010000111111001",
			2143 => "0010000101011100000100",
			2144 => "0000000010000111111001",
			2145 => "0010101100010000000100",
			2146 => "0000000010000111111001",
			2147 => "0010110101011100000100",
			2148 => "0000000010000111111001",
			2149 => "0000000010000111111001",
			2150 => "0000000010000111111001",
			2151 => "0001100000110100010100",
			2152 => "0010001111001000001000",
			2153 => "0001001110010100000100",
			2154 => "0000000010000111111001",
			2155 => "0000000010000111111001",
			2156 => "0001101111000100001000",
			2157 => "0001100110100000000100",
			2158 => "0000000010000111111001",
			2159 => "0000000010000111111001",
			2160 => "0000000010000111111001",
			2161 => "0001101111010100010000",
			2162 => "0001111101001000000100",
			2163 => "0000000010000111111001",
			2164 => "0001000010111000000100",
			2165 => "0000000010000111111001",
			2166 => "0011110011101100000100",
			2167 => "0000000010000111111001",
			2168 => "0000000010000111111001",
			2169 => "0000010111110000001000",
			2170 => "0000011001100100000100",
			2171 => "0000000010000111111001",
			2172 => "0000000010000111111001",
			2173 => "0000000010000111111001",
			2174 => "0000101010111100110100",
			2175 => "0011101010100000100100",
			2176 => "0000001100000100100000",
			2177 => "0001010110001100010000",
			2178 => "0001001001100100000100",
			2179 => "0000000010001011011101",
			2180 => "0001000001100100000100",
			2181 => "0000000010001011011101",
			2182 => "0000010110010000000100",
			2183 => "0000000010001011011101",
			2184 => "0000000010001011011101",
			2185 => "0011001001001000001100",
			2186 => "0010000011010000000100",
			2187 => "0000000010001011011101",
			2188 => "0010110111011100000100",
			2189 => "0000000010001011011101",
			2190 => "0000000010001011011101",
			2191 => "0000000010001011011101",
			2192 => "0000000010001011011101",
			2193 => "0011111001110000001100",
			2194 => "0001110110101100001000",
			2195 => "0010010110000000000100",
			2196 => "0000000010001011011101",
			2197 => "0000000010001011011101",
			2198 => "0000000010001011011101",
			2199 => "0000000010001011011101",
			2200 => "0011101010011000011000",
			2201 => "0011011010100100001000",
			2202 => "0011100000100000000100",
			2203 => "0000000010001011011101",
			2204 => "0000000010001011011101",
			2205 => "0001001000000100000100",
			2206 => "0000000010001011011101",
			2207 => "0011010101010100000100",
			2208 => "0000000010001011011101",
			2209 => "0011101001111100000100",
			2210 => "0000000010001011011101",
			2211 => "0000000010001011011101",
			2212 => "0011111110100000010000",
			2213 => "0010101100001100000100",
			2214 => "0000000010001011011101",
			2215 => "0001000010111000000100",
			2216 => "0000000010001011011101",
			2217 => "0011110010000000000100",
			2218 => "0000000010001011011101",
			2219 => "0000000010001011011101",
			2220 => "0000010111110000001100",
			2221 => "0000111011000000001000",
			2222 => "0001010110011100000100",
			2223 => "0000000010001011011101",
			2224 => "0000000010001011011101",
			2225 => "0000000010001011011101",
			2226 => "0001011110010100000100",
			2227 => "0000000010001011011101",
			2228 => "0001000011000100000100",
			2229 => "0000000010001011011101",
			2230 => "0000000010001011011101",
			2231 => "0011011011101100100000",
			2232 => "0000001110100100010100",
			2233 => "0001010110001100001000",
			2234 => "0000101100010000000100",
			2235 => "0000000010001111000001",
			2236 => "0000000010001111000001",
			2237 => "0000011001100000001000",
			2238 => "0010111110011000000100",
			2239 => "0000000010001111000001",
			2240 => "0000000010001111000001",
			2241 => "0000000010001111000001",
			2242 => "0001100100010000000100",
			2243 => "0000000010001111000001",
			2244 => "0000000011111000000100",
			2245 => "0000000010001111000001",
			2246 => "0000000010001111000001",
			2247 => "0001001110111001000000",
			2248 => "0000000000001100100000",
			2249 => "0011101101111100011000",
			2250 => "0010110011010000001000",
			2251 => "0000010110010000000100",
			2252 => "0000000010001111000001",
			2253 => "0000000010001111000001",
			2254 => "0000011101000000001000",
			2255 => "0001111010000100000100",
			2256 => "0000000010001111000001",
			2257 => "0000000010001111000001",
			2258 => "0011011001001000000100",
			2259 => "0000000010001111000001",
			2260 => "0000000010001111000001",
			2261 => "0001011011000000000100",
			2262 => "0000000010001111000001",
			2263 => "0000000010001111000001",
			2264 => "0010101101001000001100",
			2265 => "0001011000111000001000",
			2266 => "0011011010100100000100",
			2267 => "0000000010001111000001",
			2268 => "0000000010001111000001",
			2269 => "0000000010001111000001",
			2270 => "0011100000010100000100",
			2271 => "0000000010001111000001",
			2272 => "0000010110010000001000",
			2273 => "0001010011000100000100",
			2274 => "0000000010001111000001",
			2275 => "0000000010001111000001",
			2276 => "0001011110010100000100",
			2277 => "0000000010001111000001",
			2278 => "0000000010001111000001",
			2279 => "0010100001101000001000",
			2280 => "0011011010100100000100",
			2281 => "0000000010001111000001",
			2282 => "0000000010001111000001",
			2283 => "0001000010001100000100",
			2284 => "0000000010001111000001",
			2285 => "0010001111001000000100",
			2286 => "0000000010001111000001",
			2287 => "0000000010001111000001",
			2288 => "0000101100111001000000",
			2289 => "0011101010100000101100",
			2290 => "0010110111011100011100",
			2291 => "0000010110010000010000",
			2292 => "0010010110000000001100",
			2293 => "0000001010011000001000",
			2294 => "0011001110011000000100",
			2295 => "0000000010010010101101",
			2296 => "0000000010010010101101",
			2297 => "0000000010010010101101",
			2298 => "0000000010010010101101",
			2299 => "0000001111010100001000",
			2300 => "0001000110001100000100",
			2301 => "0000000010010010101101",
			2302 => "0000001010010010101101",
			2303 => "0000000010010010101101",
			2304 => "0000011101000000000100",
			2305 => "1111111010010010101101",
			2306 => "0010000011001000001000",
			2307 => "0010001010000100000100",
			2308 => "0000000010010010101101",
			2309 => "0000000010010010101101",
			2310 => "0000000010010010101101",
			2311 => "0001010010111000001100",
			2312 => "0011110100100100000100",
			2313 => "0000000010010010101101",
			2314 => "0000010110010000000100",
			2315 => "0000000010010010101101",
			2316 => "0000000010010010101101",
			2317 => "0010101100001100000100",
			2318 => "0000001010010010101101",
			2319 => "0000000010010010101101",
			2320 => "0001100100100100001100",
			2321 => "0010011111011000000100",
			2322 => "1111111010010010101101",
			2323 => "0011000011000000000100",
			2324 => "0000000010010010101101",
			2325 => "0000000010010010101101",
			2326 => "0001001000000100010000",
			2327 => "0010010101101100000100",
			2328 => "1111111010010010101101",
			2329 => "0000110011001000000100",
			2330 => "0000000010010010101101",
			2331 => "0001001001001000000100",
			2332 => "0000000010010010101101",
			2333 => "0000000010010010101101",
			2334 => "0000001100111100000100",
			2335 => "0000000010010010101101",
			2336 => "0010011001000100001000",
			2337 => "0010101001011000000100",
			2338 => "0000000010010010101101",
			2339 => "0000000010010010101101",
			2340 => "0010000101011100001000",
			2341 => "0011101111111000000100",
			2342 => "0000000010010010101101",
			2343 => "0000000010010010101101",
			2344 => "0011100000010100000100",
			2345 => "0000000010010010101101",
			2346 => "0000000010010010101101",
			2347 => "0001100100010000111100",
			2348 => "0011010101011100101100",
			2349 => "0000000111110100101000",
			2350 => "0000011001100100001000",
			2351 => "0010101100110100000100",
			2352 => "1111111010010100101001",
			2353 => "0000000010010100101001",
			2354 => "0000001101001100010000",
			2355 => "0011101111100100001000",
			2356 => "0000000000001100000100",
			2357 => "0000000010010100101001",
			2358 => "1111111010010100101001",
			2359 => "0001010101111000000100",
			2360 => "0000000010010100101001",
			2361 => "0000001010010100101001",
			2362 => "0010011101101000001000",
			2363 => "0010010101101100000100",
			2364 => "1111111010010100101001",
			2365 => "0000001010010100101001",
			2366 => "0001000001111100000100",
			2367 => "1111111010010100101001",
			2368 => "0000001010010100101001",
			2369 => "0000001010010100101001",
			2370 => "0001111100010000001000",
			2371 => "0001101100110100000100",
			2372 => "1111111010010100101001",
			2373 => "0000001010010100101001",
			2374 => "0001110110101100000100",
			2375 => "1111111010010100101001",
			2376 => "1111111010010100101001",
			2377 => "1111111010010100101001",
			2378 => "0011011010100100111100",
			2379 => "0000111011000000101100",
			2380 => "0001001100101100101000",
			2381 => "0010111110011000010000",
			2382 => "0001001001100000000100",
			2383 => "0000000010011000011101",
			2384 => "0010000011010000000100",
			2385 => "0000000010011000011101",
			2386 => "0011101100100000000100",
			2387 => "0000000010011000011101",
			2388 => "0000000010011000011101",
			2389 => "0011001010100100001000",
			2390 => "0000000100110100000100",
			2391 => "0000000010011000011101",
			2392 => "0000000010011000011101",
			2393 => "0001010011000100001000",
			2394 => "0000010011110000000100",
			2395 => "0000000010011000011101",
			2396 => "0000000010011000011101",
			2397 => "0001001001010100000100",
			2398 => "0000000010011000011101",
			2399 => "0000000010011000011101",
			2400 => "0000000010011000011101",
			2401 => "0010010011000000001000",
			2402 => "0010110101010100000100",
			2403 => "0000000010011000011101",
			2404 => "0000000010011000011101",
			2405 => "0011001001001000000100",
			2406 => "0000000010011000011101",
			2407 => "0000000010011000011101",
			2408 => "0001111100010000011100",
			2409 => "0011001100101000001100",
			2410 => "0001011000111000001000",
			2411 => "0001110101111000000100",
			2412 => "0000000010011000011101",
			2413 => "0000000010011000011101",
			2414 => "0000000010011000011101",
			2415 => "0000001010101100001100",
			2416 => "0010010011000000000100",
			2417 => "0000000010011000011101",
			2418 => "0010010101111000000100",
			2419 => "0000000010011000011101",
			2420 => "0000000010011000011101",
			2421 => "0000000010011000011101",
			2422 => "0001001110111000010100",
			2423 => "0011110100101000001100",
			2424 => "0011111001110000001000",
			2425 => "0011100101110000000100",
			2426 => "0000000010011000011101",
			2427 => "0000000010011000011101",
			2428 => "0000000010011000011101",
			2429 => "0001111001010000000100",
			2430 => "0000000010011000011101",
			2431 => "0000000010011000011101",
			2432 => "0010100001101000000100",
			2433 => "0000000010011000011101",
			2434 => "0001000010001100000100",
			2435 => "0000000010011000011101",
			2436 => "0001001111100100000100",
			2437 => "0000000010011000011101",
			2438 => "0000000010011000011101",
			2439 => "0001100100010001010100",
			2440 => "0011101010011000101100",
			2441 => "0000101110000100100000",
			2442 => "0011101111100100010100",
			2443 => "0000000000001100001100",
			2444 => "0010101110111000001000",
			2445 => "0001010110001100000100",
			2446 => "1111111010011011001001",
			2447 => "0000000010011011001001",
			2448 => "0000000010011011001001",
			2449 => "0010101110111000000100",
			2450 => "1111111010011011001001",
			2451 => "0000000010011011001001",
			2452 => "0001000110011100000100",
			2453 => "0000000010011011001001",
			2454 => "0000010110010000000100",
			2455 => "0000000010011011001001",
			2456 => "0000001010011011001001",
			2457 => "0001111101001000000100",
			2458 => "1111111010011011001001",
			2459 => "0010101100110100000100",
			2460 => "0000000010011011001001",
			2461 => "1111111010011011001001",
			2462 => "0010001111001000011000",
			2463 => "0010000101101100010000",
			2464 => "0001000011000000001000",
			2465 => "0000101010101100000100",
			2466 => "0000000010011011001001",
			2467 => "1111111010011011001001",
			2468 => "0010011010000100000100",
			2469 => "0000001010011011001001",
			2470 => "0000000010011011001001",
			2471 => "0001111100101100000100",
			2472 => "0000001010011011001001",
			2473 => "0000000010011011001001",
			2474 => "0011111110100000001100",
			2475 => "0010000000110000001000",
			2476 => "0000101011011000000100",
			2477 => "0000001010011011001001",
			2478 => "0000000010011011001001",
			2479 => "1111111010011011001001",
			2480 => "1111111010011011001001",
			2481 => "1111111010011011001001",
			2482 => "0000000000001100111100",
			2483 => "0011101010100000101100",
			2484 => "0010110110001100001000",
			2485 => "0000001110010100000100",
			2486 => "0000000010011110101101",
			2487 => "0000000010011110101101",
			2488 => "0000011000011000010000",
			2489 => "0001001100101100001100",
			2490 => "0010001001000100000100",
			2491 => "0000000010011110101101",
			2492 => "0010001111001000000100",
			2493 => "0000000010011110101101",
			2494 => "0000000010011110101101",
			2495 => "0000000010011110101101",
			2496 => "0001000111011100001100",
			2497 => "0001010101010100000100",
			2498 => "0000000010011110101101",
			2499 => "0001011001001000000100",
			2500 => "0000000010011110101101",
			2501 => "0000000010011110101101",
			2502 => "0011001001001000000100",
			2503 => "0000000010011110101101",
			2504 => "0000000010011110101101",
			2505 => "0011111001110000001100",
			2506 => "0010100011110100001000",
			2507 => "0001111000000000000100",
			2508 => "0000000010011110101101",
			2509 => "0000000010011110101101",
			2510 => "0000000010011110101101",
			2511 => "0000000010011110101101",
			2512 => "0011101010011000011100",
			2513 => "0001001110001100010100",
			2514 => "0000010110001100010000",
			2515 => "0010000011010000000100",
			2516 => "0000000010011110101101",
			2517 => "0001111001010100001000",
			2518 => "0011001001001000000100",
			2519 => "0000000010011110101101",
			2520 => "0000000010011110101101",
			2521 => "0000000010011110101101",
			2522 => "0000000010011110101101",
			2523 => "0001111000101000000100",
			2524 => "0000000010011110101101",
			2525 => "0000000010011110101101",
			2526 => "0000100111000100011000",
			2527 => "0001111101001000001000",
			2528 => "0001011000111000000100",
			2529 => "0000000010011110101101",
			2530 => "0000000010011110101101",
			2531 => "0000100101000100001100",
			2532 => "0001011111100000001000",
			2533 => "0011110111100000000100",
			2534 => "0000000010011110101101",
			2535 => "0000000010011110101101",
			2536 => "0000000010011110101101",
			2537 => "0000000010011110101101",
			2538 => "0000000010011110101101",
			2539 => "0000100100011100110000",
			2540 => "0011100001101000100000",
			2541 => "0001110111011100000100",
			2542 => "0000000010100010011001",
			2543 => "0010001001000100010000",
			2544 => "0000010111100100000100",
			2545 => "0000000010100010011001",
			2546 => "0000011001100000001000",
			2547 => "0000011000011000000100",
			2548 => "0000000010100010011001",
			2549 => "0000000010100010011001",
			2550 => "0000000010100010011001",
			2551 => "0001010110000000000100",
			2552 => "0000000010100010011001",
			2553 => "0011001100101000000100",
			2554 => "0000000010100010011001",
			2555 => "0000000010100010011001",
			2556 => "0000010110001100001100",
			2557 => "0010000101011100000100",
			2558 => "0000000010100010011001",
			2559 => "0001111000000100000100",
			2560 => "0000000010100010011001",
			2561 => "0000000010100010011001",
			2562 => "0000000010100010011001",
			2563 => "0011101111100100010100",
			2564 => "0011011010100100001100",
			2565 => "0000111011000000001000",
			2566 => "0000010001110000000100",
			2567 => "0000000010100010011001",
			2568 => "0000000010100010011001",
			2569 => "0000000010100010011001",
			2570 => "0000110001001000000100",
			2571 => "0000000010100010011001",
			2572 => "0000000010100010011001",
			2573 => "0000101110000100001100",
			2574 => "0010000101011100000100",
			2575 => "0000000010100010011001",
			2576 => "0011110000110100000100",
			2577 => "0000000010100010011001",
			2578 => "0000000010100010011001",
			2579 => "0001111100010000001100",
			2580 => "0010101000111000000100",
			2581 => "0000000010100010011001",
			2582 => "0010101011111000000100",
			2583 => "0000000010100010011001",
			2584 => "0000000010100010011001",
			2585 => "0000010000011000010000",
			2586 => "0000100011111100001000",
			2587 => "0001101100100000000100",
			2588 => "0000000010100010011001",
			2589 => "0000000010100010011001",
			2590 => "0000111011111000000100",
			2591 => "0000000010100010011001",
			2592 => "0000000010100010011001",
			2593 => "0011101110000000000100",
			2594 => "0000000010100010011001",
			2595 => "0001101111010100000100",
			2596 => "0000000010100010011001",
			2597 => "0000000010100010011001",
			2598 => "0000000111001000100000",
			2599 => "0001010110001100001000",
			2600 => "0001110111011100000100",
			2601 => "0000000010100110001101",
			2602 => "0000000010100110001101",
			2603 => "0010010110000000001100",
			2604 => "0011000101011100001000",
			2605 => "0010000101011100000100",
			2606 => "0000000010100110001101",
			2607 => "0000000010100110001101",
			2608 => "0000000010100110001101",
			2609 => "0000011110011000000100",
			2610 => "0000000010100110001101",
			2611 => "0010000011100100000100",
			2612 => "0000000010100110001101",
			2613 => "0000000010100110001101",
			2614 => "0001001000000100011100",
			2615 => "0011101010011000001100",
			2616 => "0000000110000100001000",
			2617 => "0001100001011100000100",
			2618 => "0000000010100110001101",
			2619 => "0000000010100110001101",
			2620 => "1111111010100110001101",
			2621 => "0011111101100100000100",
			2622 => "0000000010100110001101",
			2623 => "0011000111011100000100",
			2624 => "0000000010100110001101",
			2625 => "0000110011001000000100",
			2626 => "0000000010100110001101",
			2627 => "0000000010100110001101",
			2628 => "0011011010100100100100",
			2629 => "0000111011000000010000",
			2630 => "0000010111100100001100",
			2631 => "0001111000000100000100",
			2632 => "0000000010100110001101",
			2633 => "0011101110111100000100",
			2634 => "0000000010100110001101",
			2635 => "0000000010100110001101",
			2636 => "0000000010100110001101",
			2637 => "0010110101010100001000",
			2638 => "0001110110101100000100",
			2639 => "1111111010100110001101",
			2640 => "0000000010100110001101",
			2641 => "0000010001110000000100",
			2642 => "0000000010100110001101",
			2643 => "0001000011110100000100",
			2644 => "0000000010100110001101",
			2645 => "0000000010100110001101",
			2646 => "0011001100101000001000",
			2647 => "0001101100100000000100",
			2648 => "0000001010100110001101",
			2649 => "0000000010100110001101",
			2650 => "0010110101011100000100",
			2651 => "0000000010100110001101",
			2652 => "0010100000111100001000",
			2653 => "0010101001011000000100",
			2654 => "0000000010100110001101",
			2655 => "0000000010100110001101",
			2656 => "0010001001000100000100",
			2657 => "1111111010100110001101",
			2658 => "0000000010100110001101",
			2659 => "0001111101001001011000",
			2660 => "0001000111011100010100",
			2661 => "0011001011101100001100",
			2662 => "0000000010110100001000",
			2663 => "0010000101011100000100",
			2664 => "0000010010101001101001",
			2665 => "0000011010101001101001",
			2666 => "1111111010101001101001",
			2667 => "0011001110011000000100",
			2668 => "0000000010101001101001",
			2669 => "1111111010101001101001",
			2670 => "0010001111111100011000",
			2671 => "0001010011000100001000",
			2672 => "0001111101101000000100",
			2673 => "0000000010101001101001",
			2674 => "1111111010101001101001",
			2675 => "0000111011000000001000",
			2676 => "0001111000000100000100",
			2677 => "0000000010101001101001",
			2678 => "0000011010101001101001",
			2679 => "0011011110011000000100",
			2680 => "1111111010101001101001",
			2681 => "0000000010101001101001",
			2682 => "0000001011011100011100",
			2683 => "0010110011010000001100",
			2684 => "0001000110101100001000",
			2685 => "0011101010011100000100",
			2686 => "0000011010101001101001",
			2687 => "0000100010101001101001",
			2688 => "0000001010101001101001",
			2689 => "0001010011000100001000",
			2690 => "0010011010000100000100",
			2691 => "0000000010101001101001",
			2692 => "1111111010101001101001",
			2693 => "0011101111100100000100",
			2694 => "0000010010101001101001",
			2695 => "0000011010101001101001",
			2696 => "0011100010011100000100",
			2697 => "1111111010101001101001",
			2698 => "0011011011101100000100",
			2699 => "0000000010101001101001",
			2700 => "0010101011000000000100",
			2701 => "0000001010101001101001",
			2702 => "0000011010101001101001",
			2703 => "0001111000101000010100",
			2704 => "0001011001101100001100",
			2705 => "0001000101111000000100",
			2706 => "1111111010101001101001",
			2707 => "0010110011010000000100",
			2708 => "0000000010101001101001",
			2709 => "1111111010101001101001",
			2710 => "0000111100110100000100",
			2711 => "0000011010101001101001",
			2712 => "0000000010101001101001",
			2713 => "1111111010101001101001",
			2714 => "0011001110011000001100",
			2715 => "0010000011010000000100",
			2716 => "0000000010101100110101",
			2717 => "0000001011110100000100",
			2718 => "0000000010101100110101",
			2719 => "0000000010101100110101",
			2720 => "0001001100101100110100",
			2721 => "0000011000011000010100",
			2722 => "0010000101101100000100",
			2723 => "0000000010101100110101",
			2724 => "0000000110100000000100",
			2725 => "0000000010101100110101",
			2726 => "0000001010101000001000",
			2727 => "0011100100100100000100",
			2728 => "0000000010101100110101",
			2729 => "0000000010101100110101",
			2730 => "0000000010101100110101",
			2731 => "0010110011010000010100",
			2732 => "0001011000111000001000",
			2733 => "0000110011100100000100",
			2734 => "0000000010101100110101",
			2735 => "0000000010101100110101",
			2736 => "0010101101001000000100",
			2737 => "0000000010101100110101",
			2738 => "0000111100110000000100",
			2739 => "0000000010101100110101",
			2740 => "0000000010101100110101",
			2741 => "0001011011000000000100",
			2742 => "0000000010101100110101",
			2743 => "0011100010011100000100",
			2744 => "0000000010101100110101",
			2745 => "0000000010101100110101",
			2746 => "0010101100110100011100",
			2747 => "0000010001110000001000",
			2748 => "0001010001010100000100",
			2749 => "0000000010101100110101",
			2750 => "0000000010101100110101",
			2751 => "0000010111110000000100",
			2752 => "0000000010101100110101",
			2753 => "0010010011000000001000",
			2754 => "0001000000111100000100",
			2755 => "0000000010101100110101",
			2756 => "0000000010101100110101",
			2757 => "0000000100111100000100",
			2758 => "0000000010101100110101",
			2759 => "0000000010101100110101",
			2760 => "0001111001010000000100",
			2761 => "0000000010101100110101",
			2762 => "0010011000000100000100",
			2763 => "0000000010101100110101",
			2764 => "0000000010101100110101",
			2765 => "0001001100101101010100",
			2766 => "0010110111011100111100",
			2767 => "0000000010110100011100",
			2768 => "0000010110010000010000",
			2769 => "0001010110001100000100",
			2770 => "1111111010110000011001",
			2771 => "0000110101010100000100",
			2772 => "0000001010110000011001",
			2773 => "0010001001001100000100",
			2774 => "1111111010110000011001",
			2775 => "0000000010110000011001",
			2776 => "0001010101010100000100",
			2777 => "0000000010110000011001",
			2778 => "0000111100010000000100",
			2779 => "0000001010110000011001",
			2780 => "0000000010110000011001",
			2781 => "0011010011010000011000",
			2782 => "0000011001100000010000",
			2783 => "0001010011000100001000",
			2784 => "0011001010100100000100",
			2785 => "0000000010110000011001",
			2786 => "1111111010110000011001",
			2787 => "0001011100011100000100",
			2788 => "0000001010110000011001",
			2789 => "0000000010110000011001",
			2790 => "0010101101001000000100",
			2791 => "0000001010110000011001",
			2792 => "1111111010110000011001",
			2793 => "0000111101001000000100",
			2794 => "1111111010110000011001",
			2795 => "0000000010110000011001",
			2796 => "0000010111110000001100",
			2797 => "0010011010000100001000",
			2798 => "0001100100000000000100",
			2799 => "1111111010110000011001",
			2800 => "0000001010110000011001",
			2801 => "1111111010110000011001",
			2802 => "0000011110011000000100",
			2803 => "1111111010110000011001",
			2804 => "0010000011001000000100",
			2805 => "0000000010110000011001",
			2806 => "1111111010110000011001",
			2807 => "0000111011000000000100",
			2808 => "0000000010110000011001",
			2809 => "0011011011101100000100",
			2810 => "1111111010110000011001",
			2811 => "0011100101110000000100",
			2812 => "0000000010110000011001",
			2813 => "0010001111111100001000",
			2814 => "0000010001110000000100",
			2815 => "1111111010110000011001",
			2816 => "0000000010110000011001",
			2817 => "0001111000101000001000",
			2818 => "0000001011011100000100",
			2819 => "0000001010110000011001",
			2820 => "0000000010110000011001",
			2821 => "1111111010110000011001",
			2822 => "0010001001001100001000",
			2823 => "0000001011000000000100",
			2824 => "0000000010110011011101",
			2825 => "0000000010110011011101",
			2826 => "0000001100000100101000",
			2827 => "0011100001101000011100",
			2828 => "0011000011010000001000",
			2829 => "0001010110001100000100",
			2830 => "0000000010110011011101",
			2831 => "0000000010110011011101",
			2832 => "0010001001000100001000",
			2833 => "0000011000011000000100",
			2834 => "0000000010110011011101",
			2835 => "0000000010110011011101",
			2836 => "0001110011001000001000",
			2837 => "0001111101101000000100",
			2838 => "0000000010110011011101",
			2839 => "0000000010110011011101",
			2840 => "0000000010110011011101",
			2841 => "0011000101010100001000",
			2842 => "0001001010000100000100",
			2843 => "0000000010110011011101",
			2844 => "0000000010110011011101",
			2845 => "0000000010110011011101",
			2846 => "0011100101110000010000",
			2847 => "0010001111111100000100",
			2848 => "0000000010110011011101",
			2849 => "0010001001000100000100",
			2850 => "0000000010110011011101",
			2851 => "0010001111001000000100",
			2852 => "0000000010110011011101",
			2853 => "0000000010110011011101",
			2854 => "0000000010010000001000",
			2855 => "0011111001110000000100",
			2856 => "0000000010110011011101",
			2857 => "0000000010110011011101",
			2858 => "0011100000100000001100",
			2859 => "0011011010100100000100",
			2860 => "0000000010110011011101",
			2861 => "0001001100011100000100",
			2862 => "0000000010110011011101",
			2863 => "0000000010110011011101",
			2864 => "0001000001011000001000",
			2865 => "0010011101101000000100",
			2866 => "0000000010110011011101",
			2867 => "0000000010110011011101",
			2868 => "0000000100111100000100",
			2869 => "0000000010110011011101",
			2870 => "0000000010110011011101",
			2871 => "0011001110011000001100",
			2872 => "0010000011010000000100",
			2873 => "0000000010110110111001",
			2874 => "0000001011110100000100",
			2875 => "0000000010110110111001",
			2876 => "0000000010110110111001",
			2877 => "0001001100101100111000",
			2878 => "0000011000011000011000",
			2879 => "0010001010000100010100",
			2880 => "0011101111000100001000",
			2881 => "0011010111011100000100",
			2882 => "0000000010110110111001",
			2883 => "0000000010110110111001",
			2884 => "0011011011101100000100",
			2885 => "0000000010110110111001",
			2886 => "0011111110001000000100",
			2887 => "0000000010110110111001",
			2888 => "0000000010110110111001",
			2889 => "0000000010110110111001",
			2890 => "0010110011010000010100",
			2891 => "0001011000111000001000",
			2892 => "0000110011100100000100",
			2893 => "0000000010110110111001",
			2894 => "0000000010110110111001",
			2895 => "0010101101001000000100",
			2896 => "0000000010110110111001",
			2897 => "0000111100110000000100",
			2898 => "0000000010110110111001",
			2899 => "0000000010110110111001",
			2900 => "0001011011000000000100",
			2901 => "0000000010110110111001",
			2902 => "0011100010011100000100",
			2903 => "0000000010110110111001",
			2904 => "0000000010110110111001",
			2905 => "0010101100110100100000",
			2906 => "0011011110011000001100",
			2907 => "0001011110010100000100",
			2908 => "0000000010110110111001",
			2909 => "0010001111111100000100",
			2910 => "0000000010110110111001",
			2911 => "0000000010110110111001",
			2912 => "0000000100111100001100",
			2913 => "0000110000111100001000",
			2914 => "0010100000111100000100",
			2915 => "0000000010110110111001",
			2916 => "0000000010110110111001",
			2917 => "0000000010110110111001",
			2918 => "0000110001001000000100",
			2919 => "0000000010110110111001",
			2920 => "0000000010110110111001",
			2921 => "0001111001010000000100",
			2922 => "0000000010110110111001",
			2923 => "0010011000000100000100",
			2924 => "0000000010110110111001",
			2925 => "0000000010110110111001",
			2926 => "0000000100011001001100",
			2927 => "0010001001001100010100",
			2928 => "0000111100101100010000",
			2929 => "0010000011010000001000",
			2930 => "0000000100111000000100",
			2931 => "0000000010111010011101",
			2932 => "0000000010111010011101",
			2933 => "0000011001100100000100",
			2934 => "0000000010111010011101",
			2935 => "0000000010111010011101",
			2936 => "0000000010111010011101",
			2937 => "0011101111100100110000",
			2938 => "0000001100000100100000",
			2939 => "0011100001101000010000",
			2940 => "0011000011010000001000",
			2941 => "0001000011110000000100",
			2942 => "0000000010111010011101",
			2943 => "0000000010111010011101",
			2944 => "0010001001000100000100",
			2945 => "0000000010111010011101",
			2946 => "0000000010111010011101",
			2947 => "0001001100000000001000",
			2948 => "0011000011010000000100",
			2949 => "0000000010111010011101",
			2950 => "0000000010111010011101",
			2951 => "0011000101010100000100",
			2952 => "0000000010111010011101",
			2953 => "0000000010111010011101",
			2954 => "0000110000111100001100",
			2955 => "0001111000111000001000",
			2956 => "0010010110000000000100",
			2957 => "0000000010111010011101",
			2958 => "0000000010111010011101",
			2959 => "0000000010111010011101",
			2960 => "0000000010111010011101",
			2961 => "0001000011000000000100",
			2962 => "0000000010111010011101",
			2963 => "0000000010111010011101",
			2964 => "0011101111111000001000",
			2965 => "0000010110001100000100",
			2966 => "0000000010111010011101",
			2967 => "0000000010111010011101",
			2968 => "0001000001011000011000",
			2969 => "0001111101001000010100",
			2970 => "0000010111110000001100",
			2971 => "0000111111101000001000",
			2972 => "0001110110101100000100",
			2973 => "0000000010111010011101",
			2974 => "0000000010111010011101",
			2975 => "0000000010111010011101",
			2976 => "0001110110101100000100",
			2977 => "0000000010111010011101",
			2978 => "0000000010111010011101",
			2979 => "0000000010111010011101",
			2980 => "0010100001101000000100",
			2981 => "0000000010111010011101",
			2982 => "0000000010111010011101",
			2983 => "0001001100101101100000",
			2984 => "0010110111011100111100",
			2985 => "0000000010110100011100",
			2986 => "0000010110010000010000",
			2987 => "0001010110001100000100",
			2988 => "1111111010111110100001",
			2989 => "0000110101010100000100",
			2990 => "0000001010111110100001",
			2991 => "0010001001001100000100",
			2992 => "1111111010111110100001",
			2993 => "0000000010111110100001",
			2994 => "0001010101010100000100",
			2995 => "0000000010111110100001",
			2996 => "0000111100010000000100",
			2997 => "0000001010111110100001",
			2998 => "0000000010111110100001",
			2999 => "0011010011010000011000",
			3000 => "0000011001100000010000",
			3001 => "0001010011000100001000",
			3002 => "0011001010100100000100",
			3003 => "0000000010111110100001",
			3004 => "1111111010111110100001",
			3005 => "0000001011100000000100",
			3006 => "0000000010111110100001",
			3007 => "0000001010111110100001",
			3008 => "0010101101001000000100",
			3009 => "0000001010111110100001",
			3010 => "0000000010111110100001",
			3011 => "0000111101001000000100",
			3012 => "1111111010111110100001",
			3013 => "0000000010111110100001",
			3014 => "0000010111110000001100",
			3015 => "0010011010000100001000",
			3016 => "0001100100000000000100",
			3017 => "0000000010111110100001",
			3018 => "0000001010111110100001",
			3019 => "1111111010111110100001",
			3020 => "0000011110011000001100",
			3021 => "0001111100000000001000",
			3022 => "0001110011001000000100",
			3023 => "1111111010111110100001",
			3024 => "0000000010111110100001",
			3025 => "1111111010111110100001",
			3026 => "0011100111010100001000",
			3027 => "0011011010000100000100",
			3028 => "0000000010111110100001",
			3029 => "0000000010111110100001",
			3030 => "1111111010111110100001",
			3031 => "0001001011000000000100",
			3032 => "0000001010111110100001",
			3033 => "0010001001000100011000",
			3034 => "0000010001110000001000",
			3035 => "0000100111010000000100",
			3036 => "0000000010111110100001",
			3037 => "1111111010111110100001",
			3038 => "0011100101110000000100",
			3039 => "0000000010111110100001",
			3040 => "0010101100110100001000",
			3041 => "0001001110111000000100",
			3042 => "0000000010111110100001",
			3043 => "0000001010111110100001",
			3044 => "1111111010111110100001",
			3045 => "0001111000101000000100",
			3046 => "0000001010111110100001",
			3047 => "1111111010111110100001",
			3048 => "0010010011000001010100",
			3049 => "0001010001010101000100",
			3050 => "0000111011111000110000",
			3051 => "0000010111100100010000",
			3052 => "0011000110110100000100",
			3053 => "0000000011000010100101",
			3054 => "0010001001000100001000",
			3055 => "0001100011101100000100",
			3056 => "1111111011000010100101",
			3057 => "0000000011000010100101",
			3058 => "0000000011000010100101",
			3059 => "0011110010110000010000",
			3060 => "0010110011010000001000",
			3061 => "0011010110001100000100",
			3062 => "0000000011000010100101",
			3063 => "0000000011000010100101",
			3064 => "0000001100000100000100",
			3065 => "0000000011000010100101",
			3066 => "0000000011000010100101",
			3067 => "0001011100010000001000",
			3068 => "0001111000101000000100",
			3069 => "1111111011000010100101",
			3070 => "0000000011000010100101",
			3071 => "0010010110000000000100",
			3072 => "0000000011000010100101",
			3073 => "0000000011000010100101",
			3074 => "0011100010001100000100",
			3075 => "0000000011000010100101",
			3076 => "0000111000100000001100",
			3077 => "0000100111000100001000",
			3078 => "0001011100110100000100",
			3079 => "0000000011000010100101",
			3080 => "0000001011000010100101",
			3081 => "0000000011000010100101",
			3082 => "0000000011000010100101",
			3083 => "0000110011110100001000",
			3084 => "0011101001111100000100",
			3085 => "1111111011000010100101",
			3086 => "0000000011000010100101",
			3087 => "0000111100110100000100",
			3088 => "0000000011000010100101",
			3089 => "0000000011000010100101",
			3090 => "0001010001010100010100",
			3091 => "0010110101010100000100",
			3092 => "0000000011000010100101",
			3093 => "0001111000111000001000",
			3094 => "0000000011101100000100",
			3095 => "0000000011000010100101",
			3096 => "0000000011000010100101",
			3097 => "0001010010111000000100",
			3098 => "1111111011000010100101",
			3099 => "0000000011000010100101",
			3100 => "0000100010111100000100",
			3101 => "0000001011000010100101",
			3102 => "0011100000010100001100",
			3103 => "0010001111001000000100",
			3104 => "0000000011000010100101",
			3105 => "0000010011110000000100",
			3106 => "0000000011000010100101",
			3107 => "0000000011000010100101",
			3108 => "0011110011101100001000",
			3109 => "0010001010000100000100",
			3110 => "0000001011000010100101",
			3111 => "0000000011000010100101",
			3112 => "0000000011000010100101",
			3113 => "0011101110111101000000",
			3114 => "0011000110000000111100",
			3115 => "0001011011101100001000",
			3116 => "0001110111011100000100",
			3117 => "0000000011000100110001",
			3118 => "1111111011000100110001",
			3119 => "0000011000011000011100",
			3120 => "0011101010100000010000",
			3121 => "0010111110011000001000",
			3122 => "0000000111001000000100",
			3123 => "0000001011000100110001",
			3124 => "1111111011000100110001",
			3125 => "0000010111110000000100",
			3126 => "0000000011000100110001",
			3127 => "1111111011000100110001",
			3128 => "0011010111011100001000",
			3129 => "0000001011011100000100",
			3130 => "0000001011000100110001",
			3131 => "0000000011000100110001",
			3132 => "0000001011000100110001",
			3133 => "0000100100111000001100",
			3134 => "0010110101011100001000",
			3135 => "0000110101010100000100",
			3136 => "0000001011000100110001",
			3137 => "0000001011000100110001",
			3138 => "0000000011000100110001",
			3139 => "0001001001010100001000",
			3140 => "0010110011010000000100",
			3141 => "0000000011000100110001",
			3142 => "1111111011000100110001",
			3143 => "0000001011000100110001",
			3144 => "1111111011000100110001",
			3145 => "0000000101111100000100",
			3146 => "0000000011000100110001",
			3147 => "1111111011000100110001",
			3148 => "0001110011010000000100",
			3149 => "1110100011000111011101",
			3150 => "0000100111010000111100",
			3151 => "0001011000000000010100",
			3152 => "0011001110011000001000",
			3153 => "0010001001001100000100",
			3154 => "1101011011000111011101",
			3155 => "1110101011000111011101",
			3156 => "0011001010100100000100",
			3157 => "1101100011000111011101",
			3158 => "0001001001000100000100",
			3159 => "1101011011000111011101",
			3160 => "1101100011000111011101",
			3161 => "0010000101101100011000",
			3162 => "0011011110011000001100",
			3163 => "0000010110010000001000",
			3164 => "0000000001111000000100",
			3165 => "1101101011000111011101",
			3166 => "1101011011000111011101",
			3167 => "1101110011000111011101",
			3168 => "0011101101111100000100",
			3169 => "1101101011000111011101",
			3170 => "0000001110101100000100",
			3171 => "1110100011000111011101",
			3172 => "1101111011000111011101",
			3173 => "0011000110000000001100",
			3174 => "0000101000010100001000",
			3175 => "0011000111011100000100",
			3176 => "1110101011000111011101",
			3177 => "1110011011000111011101",
			3178 => "1101111011000111011101",
			3179 => "1101011011000111011101",
			3180 => "0011101110111100010100",
			3181 => "0011110100101000010000",
			3182 => "0010101101001000000100",
			3183 => "1101101011000111011101",
			3184 => "0010100001101000001000",
			3185 => "0001001001000000000100",
			3186 => "1101011011000111011101",
			3187 => "1101101011000111011101",
			3188 => "1101011011000111011101",
			3189 => "1101110011000111011101",
			3190 => "1101011011000111011101",
			3191 => "0000000100011001000100",
			3192 => "0000011001100100000100",
			3193 => "0000000011001010110001",
			3194 => "0011101010100000100100",
			3195 => "0000000111001000010100",
			3196 => "0011000101011100001100",
			3197 => "0001000111100100000100",
			3198 => "0000000011001010110001",
			3199 => "0000010001110000000100",
			3200 => "0000000011001010110001",
			3201 => "0000000011001010110001",
			3202 => "0000010011010000000100",
			3203 => "0000000011001010110001",
			3204 => "0000000011001010110001",
			3205 => "0000011000011000001000",
			3206 => "0010000101011100000100",
			3207 => "0000000011001010110001",
			3208 => "0000000011001010110001",
			3209 => "0011100001101000000100",
			3210 => "0000000011001010110001",
			3211 => "0000000011001010110001",
			3212 => "0011010101011100011000",
			3213 => "0000101010111100001100",
			3214 => "0011001100101000001000",
			3215 => "0011011011101100000100",
			3216 => "0000000011001010110001",
			3217 => "0000000011001010110001",
			3218 => "0000000011001010110001",
			3219 => "0001101010011000000100",
			3220 => "0000000011001010110001",
			3221 => "0010110011010000000100",
			3222 => "0000000011001010110001",
			3223 => "0000000011001010110001",
			3224 => "0000000011001010110001",
			3225 => "0011101111111000000100",
			3226 => "0000000011001010110001",
			3227 => "0001100011010100010000",
			3228 => "0010101100001100000100",
			3229 => "0000000011001010110001",
			3230 => "0001010010011100000100",
			3231 => "0000000011001010110001",
			3232 => "0011110010000000000100",
			3233 => "0000000011001010110001",
			3234 => "0000000011001010110001",
			3235 => "0001111101001000010000",
			3236 => "0001001101101000000100",
			3237 => "0000000011001010110001",
			3238 => "0000100111000100000100",
			3239 => "0000000011001010110001",
			3240 => "0001110110101100000100",
			3241 => "0000000011001010110001",
			3242 => "0000000011001010110001",
			3243 => "0000000011001010110001",
			3244 => "0000001100000100110000",
			3245 => "0010000011010000000100",
			3246 => "0000000011001110100101",
			3247 => "0001000110011100101000",
			3248 => "0011000011010000001100",
			3249 => "0000010110010000001000",
			3250 => "0000001010011000000100",
			3251 => "0000000011001110100101",
			3252 => "0000000011001110100101",
			3253 => "0000000011001110100101",
			3254 => "0000011000011000001100",
			3255 => "0000000010110100001000",
			3256 => "0001111000000000000100",
			3257 => "0000000011001110100101",
			3258 => "0000000011001110100101",
			3259 => "0000000011001110100101",
			3260 => "0001111100010000001000",
			3261 => "0011001001001000000100",
			3262 => "0000000011001110100101",
			3263 => "0000000011001110100101",
			3264 => "0010001111001000000100",
			3265 => "0000000011001110100101",
			3266 => "0000000011001110100101",
			3267 => "0000000011001110100101",
			3268 => "0011100101110000011000",
			3269 => "0000010110010000001100",
			3270 => "0001001011111000001000",
			3271 => "0001000011000000000100",
			3272 => "0000000011001110100101",
			3273 => "0000000011001110100101",
			3274 => "0000000011001110100101",
			3275 => "0011010111011100000100",
			3276 => "1111111011001110100101",
			3277 => "0011011100101000000100",
			3278 => "0000000011001110100101",
			3279 => "0000000011001110100101",
			3280 => "0000000010010000001100",
			3281 => "0000010110010000000100",
			3282 => "0000000011001110100101",
			3283 => "0000110001001000000100",
			3284 => "0000000011001110100101",
			3285 => "0000000011001110100101",
			3286 => "0011011011101100001100",
			3287 => "0001100100010000000100",
			3288 => "0000000011001110100101",
			3289 => "0000000011111000000100",
			3290 => "0000000011001110100101",
			3291 => "0000000011001110100101",
			3292 => "0001101101000100001100",
			3293 => "0011010111011100000100",
			3294 => "0000000011001110100101",
			3295 => "0001011101101100000100",
			3296 => "0000000011001110100101",
			3297 => "0000000011001110100101",
			3298 => "0001101111000100001000",
			3299 => "0000101001111000000100",
			3300 => "0000001011001110100101",
			3301 => "0000000011001110100101",
			3302 => "0001100000110100000100",
			3303 => "0000000011001110100101",
			3304 => "0000000011001110100101",
			3305 => "0001010001101001011100",
			3306 => "0010110111011100111000",
			3307 => "0000100100101000011000",
			3308 => "0011011011101100010000",
			3309 => "0011000110110100000100",
			3310 => "0000001011010010101001",
			3311 => "0010000101011100000100",
			3312 => "1111111011010010101001",
			3313 => "0011001110011000000100",
			3314 => "0000000011010010101001",
			3315 => "0000000011010010101001",
			3316 => "0001100011000100000100",
			3317 => "0000000011010010101001",
			3318 => "0000001011010010101001",
			3319 => "0011101010011000001000",
			3320 => "0001001001010100000100",
			3321 => "1111111011010010101001",
			3322 => "0000000011010010101001",
			3323 => "0010001111111100001000",
			3324 => "0000111111101000000100",
			3325 => "1111111011010010101001",
			3326 => "0000000011010010101001",
			3327 => "0010001111001000001000",
			3328 => "0001100100101000000100",
			3329 => "0000001011010010101001",
			3330 => "0000000011010010101001",
			3331 => "0010001010000100000100",
			3332 => "1111111011010010101001",
			3333 => "0000000011010010101001",
			3334 => "0000001100000100011000",
			3335 => "0011101001101100010100",
			3336 => "0010010110000000001000",
			3337 => "0010110101010100000100",
			3338 => "0000000011010010101001",
			3339 => "0000000011010010101001",
			3340 => "0000011101000000000100",
			3341 => "1111111011010010101001",
			3342 => "0011010101101100000100",
			3343 => "0000000011010010101001",
			3344 => "0000000011010010101001",
			3345 => "0000000011010010101001",
			3346 => "0001111100000000000100",
			3347 => "0000000011010010101001",
			3348 => "0001010000111000000100",
			3349 => "1111111011010010101001",
			3350 => "0000000011010010101001",
			3351 => "0011101010100000000100",
			3352 => "0000000011010010101001",
			3353 => "0001011110010100000100",
			3354 => "0000001011010010101001",
			3355 => "0010001111111100001100",
			3356 => "0011011010100100001000",
			3357 => "0010110101010100000100",
			3358 => "1111111011010010101001",
			3359 => "0000000011010010101001",
			3360 => "0000000011010010101001",
			3361 => "0001001000100000001000",
			3362 => "0000110001001000000100",
			3363 => "0000000011010010101001",
			3364 => "1111111011010010101001",
			3365 => "0000110000111100000100",
			3366 => "0000000011010010101001",
			3367 => "0001011010110100000100",
			3368 => "0000001011010010101001",
			3369 => "0000000011010010101001",
			3370 => "0001100100010001011100",
			3371 => "0001111000000000100000",
			3372 => "0000110011000100011100",
			3373 => "0011001100101000011000",
			3374 => "0011000101010100010000",
			3375 => "0001101110001100001000",
			3376 => "0000011001100100000100",
			3377 => "1111111011010101100101",
			3378 => "0000001011010101100101",
			3379 => "0000011001100000000100",
			3380 => "1111111011010101100101",
			3381 => "0000000011010101100101",
			3382 => "0001001010000100000100",
			3383 => "0000000011010101100101",
			3384 => "0000001011010101100101",
			3385 => "1111111011010101100101",
			3386 => "1111111011010101100101",
			3387 => "0001010001101000100000",
			3388 => "0010010110000000001100",
			3389 => "0001110110101100001000",
			3390 => "0001111100010000000100",
			3391 => "0000000011010101100101",
			3392 => "0000000011010101100101",
			3393 => "0000001011010101100101",
			3394 => "0000000010010000001100",
			3395 => "0001001100000000001000",
			3396 => "0001111001010100000100",
			3397 => "1111111011010101100101",
			3398 => "0000000011010101100101",
			3399 => "0000001011010101100101",
			3400 => "0001111100110000000100",
			3401 => "0000000011010101100101",
			3402 => "1111111011010101100101",
			3403 => "0010011010000100001000",
			3404 => "0000011001100100000100",
			3405 => "1111111011010101100101",
			3406 => "0000001011010101100101",
			3407 => "0010010011000000001000",
			3408 => "0000010111110000000100",
			3409 => "0000000011010101100101",
			3410 => "1111111011010101100101",
			3411 => "0000100101000100001000",
			3412 => "0010100001101000000100",
			3413 => "0000001011010101100101",
			3414 => "0000000011010101100101",
			3415 => "1111111011010101100101",
			3416 => "1111111011010101100101",
			3417 => "0001010001101001011000",
			3418 => "0010110111011100111000",
			3419 => "0000100100101000011000",
			3420 => "0001010110001100001000",
			3421 => "0001110111011100000100",
			3422 => "0000000011011001110001",
			3423 => "1111111011011001110001",
			3424 => "0010000011010000000100",
			3425 => "0000000011011001110001",
			3426 => "0001010001011000001000",
			3427 => "0011000111011100000100",
			3428 => "0000001011011001110001",
			3429 => "0000000011011001110001",
			3430 => "0000000011011001110001",
			3431 => "0011101010011000001000",
			3432 => "0001001001010100000100",
			3433 => "1111111011011001110001",
			3434 => "0000000011011001110001",
			3435 => "0010001111111100001000",
			3436 => "0000111111101000000100",
			3437 => "1111111011011001110001",
			3438 => "0000000011011001110001",
			3439 => "0010001111001000001000",
			3440 => "0001100100101000000100",
			3441 => "0000001011011001110001",
			3442 => "0000000011011001110001",
			3443 => "0010001010000100000100",
			3444 => "1111111011011001110001",
			3445 => "0000000011011001110001",
			3446 => "0000001100000100011000",
			3447 => "0011101001101100010100",
			3448 => "0010010110000000001000",
			3449 => "0010110101010100000100",
			3450 => "0000000011011001110001",
			3451 => "0000000011011001110001",
			3452 => "0000011101000000000100",
			3453 => "1111111011011001110001",
			3454 => "0011010101101100000100",
			3455 => "0000000011011001110001",
			3456 => "0000000011011001110001",
			3457 => "0000001011011001110001",
			3458 => "0010100011110100000100",
			3459 => "1111111011011001110001",
			3460 => "0000000011011001110001",
			3461 => "0001111000000000000100",
			3462 => "0000000011011001110001",
			3463 => "0001011110010100000100",
			3464 => "0000001011011001110001",
			3465 => "0010001111111100001100",
			3466 => "0011101011110000000100",
			3467 => "1111111011011001110001",
			3468 => "0000000100111100000100",
			3469 => "0000000011011001110001",
			3470 => "1111111011011001110001",
			3471 => "0000010111100100001100",
			3472 => "0011011110011000000100",
			3473 => "0000000011011001110001",
			3474 => "0010100001101000000100",
			3475 => "0000001011011001110001",
			3476 => "0000000011011001110001",
			3477 => "0000001100111100001000",
			3478 => "0010101010011100000100",
			3479 => "0000000011011001110001",
			3480 => "0000001011011001110001",
			3481 => "0011110110000100000100",
			3482 => "1111111011011001110001",
			3483 => "0000000011011001110001",
			3484 => "0011011011101100100000",
			3485 => "0000111011000000011100",
			3486 => "0010101001011000011000",
			3487 => "0011000110110100001000",
			3488 => "0000000000110100000100",
			3489 => "0000000011011110000101",
			3490 => "0000000011011110000101",
			3491 => "0010000101011100000100",
			3492 => "1111111011011110000101",
			3493 => "0011000011010000001000",
			3494 => "0001100101110100000100",
			3495 => "0000000011011110000101",
			3496 => "0000000011011110000101",
			3497 => "0000000011011110000101",
			3498 => "0000001011011110000101",
			3499 => "1111111011011110000101",
			3500 => "0011000101011100110000",
			3501 => "0011010101011100101100",
			3502 => "0011111110100000011100",
			3503 => "0010101101001000001100",
			3504 => "0011000101010100001000",
			3505 => "0000110101111000000100",
			3506 => "0000000011011110000101",
			3507 => "0000001011011110000101",
			3508 => "0000000011011110000101",
			3509 => "0011000101010100001000",
			3510 => "0001101010100000000100",
			3511 => "0000000011011110000101",
			3512 => "0000000011011110000101",
			3513 => "0010011101101000000100",
			3514 => "0000000011011110000101",
			3515 => "0000000011011110000101",
			3516 => "0000010111110000001000",
			3517 => "0000111001010100000100",
			3518 => "0000000011011110000101",
			3519 => "0000000011011110000101",
			3520 => "0000110011001000000100",
			3521 => "0000000011011110000101",
			3522 => "1111111011011110000101",
			3523 => "0000000011011110000101",
			3524 => "0010101010011100100100",
			3525 => "0000000000001100010100",
			3526 => "0011100101110000010000",
			3527 => "0010001001000100001000",
			3528 => "0000010111110000000100",
			3529 => "0000000011011110000101",
			3530 => "1111111011011110000101",
			3531 => "0001111000000000000100",
			3532 => "0000000011011110000101",
			3533 => "0000000011011110000101",
			3534 => "0000000011011110000101",
			3535 => "0011010111011100001000",
			3536 => "0000011001100000000100",
			3537 => "1111111011011110000101",
			3538 => "0000000011011110000101",
			3539 => "0001111101001000000100",
			3540 => "0000000011011110000101",
			3541 => "0000000011011110000101",
			3542 => "0010101100001100000100",
			3543 => "0000001011011110000101",
			3544 => "0011101001110000001100",
			3545 => "0000000100011000000100",
			3546 => "0000000011011110000101",
			3547 => "0010001111001000000100",
			3548 => "1111111011011110000101",
			3549 => "0000000011011110000101",
			3550 => "0010100001101000000100",
			3551 => "0000000011011110000101",
			3552 => "0000000011011110000101",
			3553 => "0001110001010001011000",
			3554 => "0001001100110101010000",
			3555 => "0000111011000000110000",
			3556 => "0010011101101000100000",
			3557 => "0001001000000100010000",
			3558 => "0010001111111100001000",
			3559 => "0011000110110100000100",
			3560 => "0000000011100000111001",
			3561 => "1111111011100000111001",
			3562 => "0011001010100100000100",
			3563 => "0000001011100000111001",
			3564 => "0000000011100000111001",
			3565 => "0001111000000100001000",
			3566 => "0001000110101100000100",
			3567 => "0000000011100000111001",
			3568 => "0000000011100000111001",
			3569 => "0000100111000100000100",
			3570 => "0000001011100000111001",
			3571 => "0000000011100000111001",
			3572 => "0010110111011100000100",
			3573 => "0000000011100000111001",
			3574 => "0000001000110100001000",
			3575 => "0000100100101000000100",
			3576 => "0000000011100000111001",
			3577 => "0000000011100000111001",
			3578 => "1111111011100000111001",
			3579 => "0010011101101000001000",
			3580 => "0001111100010000000100",
			3581 => "1111111011100000111001",
			3582 => "0000000011100000111001",
			3583 => "0010001111111100001000",
			3584 => "0010011010000100000100",
			3585 => "0000000011100000111001",
			3586 => "0000000011100000111001",
			3587 => "0000100111010000001000",
			3588 => "0011100100000000000100",
			3589 => "0000000011100000111001",
			3590 => "0000000011100000111001",
			3591 => "0001111101001000000100",
			3592 => "0000000011100000111001",
			3593 => "1111111011100000111001",
			3594 => "0000110010111000000100",
			3595 => "0000000011100000111001",
			3596 => "0000000011100000111001",
			3597 => "0000000011100000111001",
			3598 => "0001100100010001101000",
			3599 => "0011001100101000111100",
			3600 => "0010101100001100111000",
			3601 => "0000000011101100011100",
			3602 => "0000010001110000001100",
			3603 => "0010001001001100000100",
			3604 => "1111111011100100001111",
			3605 => "0010110011010000000100",
			3606 => "0000000011100100001111",
			3607 => "1111111011100100001111",
			3608 => "0011101000100000001000",
			3609 => "0010111010100100000100",
			3610 => "0000001011100100001111",
			3611 => "1111111011100100001111",
			3612 => "0001010110101100000100",
			3613 => "0000001011100100001111",
			3614 => "0000001011100100001111",
			3615 => "0011101001101100001100",
			3616 => "0000011000011000001000",
			3617 => "0000010000011000000100",
			3618 => "0000000011100100001111",
			3619 => "1111111011100100001111",
			3620 => "0000001011100100001111",
			3621 => "0001011001011000001000",
			3622 => "0001011001010100000100",
			3623 => "0000000011100100001111",
			3624 => "1111111011100100001111",
			3625 => "0001111000000000000100",
			3626 => "0000000011100100001111",
			3627 => "0000001011100100001111",
			3628 => "1111111011100100001111",
			3629 => "0000110001001000011000",
			3630 => "0011100101110000010000",
			3631 => "0000000111101000001000",
			3632 => "0000000110000100000100",
			3633 => "1111111011100100001111",
			3634 => "0000000011100100001111",
			3635 => "0000000000010000000100",
			3636 => "1111110011100100001111",
			3637 => "1111111011100100001111",
			3638 => "0001101111111000000100",
			3639 => "0000001011100100001111",
			3640 => "1111111011100100001111",
			3641 => "0000000100111100010000",
			3642 => "0011101111111000001100",
			3643 => "0000000010111100001000",
			3644 => "0010101100110100000100",
			3645 => "0000001011100100001111",
			3646 => "0000000011100100001111",
			3647 => "1111111011100100001111",
			3648 => "0000001011100100001111",
			3649 => "1111111011100100001111",
			3650 => "1111111011100100001111",
			3651 => "0010001001001100001100",
			3652 => "0000001000100000000100",
			3653 => "0000000011100101101001",
			3654 => "0001000110011100000100",
			3655 => "1111111011100101101001",
			3656 => "0000000011100101101001",
			3657 => "0001110001010000100000",
			3658 => "0000000111110100011000",
			3659 => "0011100110100000010000",
			3660 => "0000011001100100000100",
			3661 => "1111111011100101101001",
			3662 => "0011100100100100001000",
			3663 => "0001101111000100000100",
			3664 => "0000000011100101101001",
			3665 => "1111111011100101101001",
			3666 => "0000000011100101101001",
			3667 => "0011101111110000000100",
			3668 => "1111111011100101101001",
			3669 => "0000000011100101101001",
			3670 => "0001010011000100000100",
			3671 => "0000000011100101101001",
			3672 => "0000001011100101101001",
			3673 => "1111111011100101101001",
			3674 => "0010001001001100001100",
			3675 => "0000001000100000000100",
			3676 => "0000000011100111001101",
			3677 => "0001000110011100000100",
			3678 => "1111111011100111001101",
			3679 => "0000000011100111001101",
			3680 => "0001110001010000100100",
			3681 => "0000000111110100011100",
			3682 => "0011100110100000010100",
			3683 => "0000011001100100000100",
			3684 => "1111111011100111001101",
			3685 => "0011101010011000001000",
			3686 => "0001101111000100000100",
			3687 => "0000000011100111001101",
			3688 => "1111111011100111001101",
			3689 => "0010001111111100000100",
			3690 => "0000000011100111001101",
			3691 => "0000001011100111001101",
			3692 => "0011101111110000000100",
			3693 => "1111111011100111001101",
			3694 => "0000000011100111001101",
			3695 => "0001010011000100000100",
			3696 => "0000000011100111001101",
			3697 => "0000001011100111001101",
			3698 => "1111111011100111001101",
			3699 => "0000100111000100110000",
			3700 => "0000000111110100101000",
			3701 => "0000011001100100000100",
			3702 => "1111111011101001000001",
			3703 => "0011100110100000011100",
			3704 => "0010110101011100010000",
			3705 => "0000111110111000001000",
			3706 => "0011101001101100000100",
			3707 => "0000000011101001000001",
			3708 => "0000000011101001000001",
			3709 => "0001001110111000000100",
			3710 => "1111111011101001000001",
			3711 => "0000000011101001000001",
			3712 => "0011001100101000000100",
			3713 => "0000000011101001000001",
			3714 => "0001111100010000000100",
			3715 => "1111111011101001000001",
			3716 => "0000000011101001000001",
			3717 => "0010111110011000000100",
			3718 => "0000000011101001000001",
			3719 => "1111111011101001000001",
			3720 => "0011101111110000000100",
			3721 => "0000001011101001000001",
			3722 => "0000000011101001000001",
			3723 => "0000010000011000001000",
			3724 => "0011011011101100000100",
			3725 => "0000000011101001000001",
			3726 => "0000000011101001000001",
			3727 => "1111111011101001000001",
			3728 => "0010110101011100110100",
			3729 => "0010001001001100001000",
			3730 => "0000001100001100000100",
			3731 => "0000000011101011100101",
			3732 => "0000000011101011100101",
			3733 => "0000100111000100100100",
			3734 => "0001010110001100001100",
			3735 => "0001000001100100001000",
			3736 => "0001101001000100000100",
			3737 => "0000000011101011100101",
			3738 => "0000000011101011100101",
			3739 => "0000000011101011100101",
			3740 => "0010101100110100010000",
			3741 => "0000011001100100001000",
			3742 => "0001111100010000000100",
			3743 => "0000000011101011100101",
			3744 => "0000000011101011100101",
			3745 => "0011101001101100000100",
			3746 => "0000000011101011100101",
			3747 => "0000000011101011100101",
			3748 => "0001001110111000000100",
			3749 => "0000000011101011100101",
			3750 => "0000000011101011100101",
			3751 => "0000010000011000000100",
			3752 => "0000000011101011100101",
			3753 => "0000000011101011100101",
			3754 => "0011001100101000001000",
			3755 => "0000111001010000000100",
			3756 => "0000000011101011100101",
			3757 => "0000000011101011100101",
			3758 => "0001000001111100010000",
			3759 => "0010011101101000000100",
			3760 => "0000000011101011100101",
			3761 => "0000101000011100000100",
			3762 => "0000000011101011100101",
			3763 => "0011101111110100000100",
			3764 => "0000000011101011100101",
			3765 => "0000000011101011100101",
			3766 => "0000101011010100000100",
			3767 => "0000000011101011100101",
			3768 => "0000000011101011100101",
			3769 => "0000001011011101000000",
			3770 => "0011001100101000101000",
			3771 => "0010001001001100001100",
			3772 => "0000001001011000000100",
			3773 => "0000000011101111001001",
			3774 => "0001101001111100000100",
			3775 => "0000000011101111001001",
			3776 => "0000000011101111001001",
			3777 => "0011101001101100010000",
			3778 => "0011110111010100001100",
			3779 => "0001000111100100000100",
			3780 => "0000000011101111001001",
			3781 => "0000010001110000000100",
			3782 => "0000000011101111001001",
			3783 => "0000000011101111001001",
			3784 => "0000000011101111001001",
			3785 => "0000101010111100001000",
			3786 => "0001111100010000000100",
			3787 => "0000000011101111001001",
			3788 => "0000000011101111001001",
			3789 => "0000000011101111001001",
			3790 => "0000110001001000010000",
			3791 => "0010011101101000001000",
			3792 => "0010010110000000000100",
			3793 => "0000000011101111001001",
			3794 => "0000000011101111001001",
			3795 => "0010110101010100000100",
			3796 => "0000000011101111001001",
			3797 => "0000000011101111001001",
			3798 => "0010101100110100000100",
			3799 => "0000000011101111001001",
			3800 => "0000000011101111001001",
			3801 => "0001010001101000011000",
			3802 => "0011110001000000001000",
			3803 => "0000010110110100000100",
			3804 => "1111111011101111001001",
			3805 => "0000000011101111001001",
			3806 => "0001011100011100001100",
			3807 => "0001100100010000001000",
			3808 => "0001000110000000000100",
			3809 => "0000000011101111001001",
			3810 => "0000000011101111001001",
			3811 => "0000000011101111001001",
			3812 => "0000000011101111001001",
			3813 => "0001101101000100001100",
			3814 => "0011010111011100000100",
			3815 => "0000000011101111001001",
			3816 => "0011011001001000000100",
			3817 => "0000000011101111001001",
			3818 => "0000000011101111001001",
			3819 => "0001111000101000001100",
			3820 => "0001000001011000000100",
			3821 => "0000000011101111001001",
			3822 => "0011011110011000000100",
			3823 => "0000000011101111001001",
			3824 => "0000000011101111001001",
			3825 => "0000000011101111001001",
			3826 => "0000000000001100110100",
			3827 => "0011101010100000100100",
			3828 => "0000000111001000011100",
			3829 => "0000111101000000001000",
			3830 => "0001000011110000000100",
			3831 => "0000000011110010110101",
			3832 => "0000000011110010110101",
			3833 => "0010010110000000001100",
			3834 => "0010001001001100000100",
			3835 => "0000000011110010110101",
			3836 => "0000010001110000000100",
			3837 => "0000000011110010110101",
			3838 => "0000000011110010110101",
			3839 => "0000011110011000000100",
			3840 => "0000000011110010110101",
			3841 => "0000000011110010110101",
			3842 => "0000011000011000000100",
			3843 => "0000000011110010110101",
			3844 => "0000000011110010110101",
			3845 => "0001011011000000001000",
			3846 => "0011001010100100000100",
			3847 => "0000000011110010110101",
			3848 => "0000000011110010110101",
			3849 => "0001011001101100000100",
			3850 => "0000000011110010110101",
			3851 => "0000000011110010110101",
			3852 => "0001010001101000100000",
			3853 => "0001001100101000001100",
			3854 => "0010011100101000000100",
			3855 => "0000000011110010110101",
			3856 => "0011000111011100000100",
			3857 => "0000000011110010110101",
			3858 => "0000000011110010110101",
			3859 => "0000010110001100001100",
			3860 => "0000010111110000001000",
			3861 => "0000010001110000000100",
			3862 => "0000000011110010110101",
			3863 => "0000000011110010110101",
			3864 => "0000000011110010110101",
			3865 => "0000011011101100000100",
			3866 => "0000000011110010110101",
			3867 => "0000000011110010110101",
			3868 => "0001101101000100001100",
			3869 => "0000110001001000000100",
			3870 => "0000000011110010110101",
			3871 => "0010001111001000000100",
			3872 => "0000000011110010110101",
			3873 => "0000000011110010110101",
			3874 => "0010101100001100001000",
			3875 => "0010001001000100000100",
			3876 => "0000000011110010110101",
			3877 => "0000000011110010110101",
			3878 => "0001011101101100001000",
			3879 => "0011111000101100000100",
			3880 => "0000000011110010110101",
			3881 => "0000000011110010110101",
			3882 => "0000110001101000000100",
			3883 => "0000000011110010110101",
			3884 => "0000000011110010110101",
			3885 => "0001111000101000110000",
			3886 => "0011101110111100101100",
			3887 => "0000001000000100000100",
			3888 => "1111111011110100101001",
			3889 => "0000010001110000010000",
			3890 => "0001100010011000001100",
			3891 => "0000011001100100000100",
			3892 => "1111111011110100101001",
			3893 => "0000001010101100000100",
			3894 => "0000000011110100101001",
			3895 => "1111111011110100101001",
			3896 => "0000001011110100101001",
			3897 => "0010111100101000010000",
			3898 => "0010101100110100001000",
			3899 => "0001010110001100000100",
			3900 => "0000000011110100101001",
			3901 => "0000001011110100101001",
			3902 => "0001001100001100000100",
			3903 => "0000000011110100101001",
			3904 => "1111111011110100101001",
			3905 => "0001100010011100000100",
			3906 => "1111111011110100101001",
			3907 => "0000001011110100101001",
			3908 => "1111111011110100101001",
			3909 => "0011001110011000001000",
			3910 => "0001000101010100000100",
			3911 => "1111111011110100101001",
			3912 => "0000001011110100101001",
			3913 => "1111111011110100101001",
			3914 => "0001011100001100111000",
			3915 => "0010110111011100110000",
			3916 => "0010001111111100010000",
			3917 => "0011000110110100000100",
			3918 => "0000000011110111101101",
			3919 => "0011111100000100000100",
			3920 => "0000000011110111101101",
			3921 => "0000111111101000000100",
			3922 => "0000000011110111101101",
			3923 => "0000000011110111101101",
			3924 => "0011010011010000011000",
			3925 => "0011011011101100001100",
			3926 => "0000101001111100000100",
			3927 => "0000000011110111101101",
			3928 => "0011100000010100000100",
			3929 => "0000000011110111101101",
			3930 => "0000000011110111101101",
			3931 => "0000010110010000000100",
			3932 => "0000000011110111101101",
			3933 => "0001100011101100000100",
			3934 => "0000000011110111101101",
			3935 => "0000000011110111101101",
			3936 => "0000001011101000000100",
			3937 => "0000000011110111101101",
			3938 => "0000000011110111101101",
			3939 => "0010000101011100000100",
			3940 => "0000000011110111101101",
			3941 => "0000000011110111101101",
			3942 => "0010101100110100100000",
			3943 => "0010110101010100010000",
			3944 => "0000111000100000001100",
			3945 => "0010010110000000000100",
			3946 => "0000000011110111101101",
			3947 => "0001001001011000000100",
			3948 => "0000000011110111101101",
			3949 => "0000000011110111101101",
			3950 => "0000000011110111101101",
			3951 => "0000010001110000000100",
			3952 => "0000000011110111101101",
			3953 => "0001110001010000001000",
			3954 => "0000110001001000000100",
			3955 => "0000000011110111101101",
			3956 => "0000000011110111101101",
			3957 => "0000000011110111101101",
			3958 => "0001111001010000000100",
			3959 => "0000000011110111101101",
			3960 => "0010011000000100000100",
			3961 => "0000000011110111101101",
			3962 => "0000000011110111101101",
			3963 => "0011100010001000111100",
			3964 => "0001010110001100001100",
			3965 => "0001001001100100000100",
			3966 => "0000000011111001101001",
			3967 => "0000010011110000000100",
			3968 => "1111111011111001101001",
			3969 => "0000000011111001101001",
			3970 => "0010001001001100010100",
			3971 => "0001101010011000010000",
			3972 => "0001101001111100001100",
			3973 => "0001011001001000000100",
			3974 => "0000000011111001101001",
			3975 => "0000001110010000000100",
			3976 => "1111111011111001101001",
			3977 => "0000000011111001101001",
			3978 => "0000000011111001101001",
			3979 => "1111111011111001101001",
			3980 => "0011001010100100001000",
			3981 => "0000001110100000000100",
			3982 => "0000001011111001101001",
			3983 => "0000000011111001101001",
			3984 => "0001011000000100000100",
			3985 => "1111111011111001101001",
			3986 => "0011111110100100001000",
			3987 => "0000001011011000000100",
			3988 => "0000000011111001101001",
			3989 => "1111111011111001101001",
			3990 => "0000010110010000000100",
			3991 => "0000001011111001101001",
			3992 => "0000000011111001101001",
			3993 => "1111111011111001101001",
			3994 => "0000100111010000111100",
			3995 => "0011101010001100110000",
			3996 => "0000000000001100100000",
			3997 => "0010000011010000000100",
			3998 => "0000000011111100101101",
			3999 => "0011101101111100010000",
			4000 => "0011000011010000001000",
			4001 => "0011110001010100000100",
			4002 => "0000000011111100101101",
			4003 => "0000000011111100101101",
			4004 => "0000011000011000000100",
			4005 => "0000000011111100101101",
			4006 => "0000000011111100101101",
			4007 => "0001001111011000000100",
			4008 => "0000000011111100101101",
			4009 => "0001011001101100000100",
			4010 => "0000000011111100101101",
			4011 => "0000000011111100101101",
			4012 => "0010101110111000001000",
			4013 => "0011010111011100000100",
			4014 => "0000000011111100101101",
			4015 => "0000000011111100101101",
			4016 => "0000110011110100000100",
			4017 => "0000000011111100101101",
			4018 => "0000000011111100101101",
			4019 => "0001000110011100001000",
			4020 => "0000010110010000000100",
			4021 => "0000000011111100101101",
			4022 => "0000000011111100101101",
			4023 => "0000000011111100101101",
			4024 => "0001111100010000001100",
			4025 => "0010101000111000000100",
			4026 => "0000000011111100101101",
			4027 => "0010111010100100000100",
			4028 => "0000000011111100101101",
			4029 => "0000000011111100101101",
			4030 => "0010101000000000000100",
			4031 => "0000000011111100101101",
			4032 => "0000000111110100001000",
			4033 => "0000011000111100000100",
			4034 => "0000000011111100101101",
			4035 => "0000000011111100101101",
			4036 => "0000001110110100000100",
			4037 => "0000000011111100101101",
			4038 => "0000010000011000001000",
			4039 => "0000011001100100000100",
			4040 => "0000000011111100101101",
			4041 => "0000000011111100101101",
			4042 => "0000000011111100101101",
			4043 => "0001111101001001010000",
			4044 => "0001000111011100010100",
			4045 => "0011001011101100001100",
			4046 => "0000000010110100001000",
			4047 => "0010000101011100000100",
			4048 => "0000001011111111111001",
			4049 => "0000010011111111111001",
			4050 => "1111111011111111111001",
			4051 => "0011001110011000000100",
			4052 => "0000000011111111111001",
			4053 => "1111111011111111111001",
			4054 => "0010000101011100010000",
			4055 => "0010010110000000001000",
			4056 => "0001011110111000000100",
			4057 => "1111111011111111111001",
			4058 => "0000000011111111111001",
			4059 => "0001010001010100000100",
			4060 => "0000010011111111111001",
			4061 => "1111111011111111111001",
			4062 => "0000001011011100011000",
			4063 => "0011001001001000010000",
			4064 => "0000011000011000001000",
			4065 => "0011101001101100000100",
			4066 => "0000001011111111111001",
			4067 => "0000010011111111111001",
			4068 => "0010110011010000000100",
			4069 => "0000010011111111111001",
			4070 => "0000010011111111111001",
			4071 => "0000111100101100000100",
			4072 => "1111111011111111111001",
			4073 => "0000001011111111111001",
			4074 => "0011011010100100001100",
			4075 => "0001100010000000000100",
			4076 => "1111111011111111111001",
			4077 => "0001101000101100000100",
			4078 => "0000010011111111111001",
			4079 => "1111111011111111111001",
			4080 => "0001101010011000000100",
			4081 => "1111111011111111111001",
			4082 => "0000010011111111111001",
			4083 => "0001111000101000010100",
			4084 => "0001011001101100001100",
			4085 => "0001000101111000000100",
			4086 => "1111111011111111111001",
			4087 => "0010110011010000000100",
			4088 => "0000000011111111111001",
			4089 => "1111111011111111111001",
			4090 => "0000000000100100000100",
			4091 => "0000010011111111111001",
			4092 => "0000000011111111111001",
			4093 => "1111111011111111111001",
			4094 => "0000000111000001001100",
			4095 => "0011101001101100110000",
			4096 => "0000000111001000100000",
			4097 => "0010010110000000010100",
			4098 => "0001010110001100001100",
			4099 => "0001000000011000000100",
			4100 => "0000000100000011100101",
			4101 => "0001001000011000000100",
			4102 => "0000000100000011100101",
			4103 => "0000000100000011100101",
			4104 => "0010001001001100000100",
			4105 => "0000000100000011100101",
			4106 => "0000000100000011100101",
			4107 => "0000011110011000001000",
			4108 => "0011011011101100000100",
			4109 => "0000000100000011100101",
			4110 => "0000000100000011100101",
			4111 => "0000000100000011100101",
			4112 => "0000011000011000001000",
			4113 => "0010000101011100000100",
			4114 => "0000000100000011100101",
			4115 => "0000000100000011100101",
			4116 => "0010001010000100000100",
			4117 => "0000000100000011100101",
			4118 => "0000000100000011100101",
			4119 => "0010001111011000011000",
			4120 => "0010001111111100010000",
			4121 => "0001010001111100001100",
			4122 => "0001011110001100001000",
			4123 => "0001011101101000000100",
			4124 => "0000000100000011100101",
			4125 => "0000000100000011100101",
			4126 => "0000000100000011100101",
			4127 => "0000000100000011100101",
			4128 => "0011001100101000000100",
			4129 => "0000000100000011100101",
			4130 => "0000000100000011100101",
			4131 => "0000000100000011100101",
			4132 => "0011011010100100001100",
			4133 => "0011111111010100000100",
			4134 => "0000000100000011100101",
			4135 => "0001101101100000000100",
			4136 => "0000000100000011100101",
			4137 => "0000000100000011100101",
			4138 => "0010101100001100010100",
			4139 => "0010010101101100000100",
			4140 => "0000000100000011100101",
			4141 => "0001111001010000001000",
			4142 => "0011010101010100000100",
			4143 => "0000000100000011100101",
			4144 => "0000000100000011100101",
			4145 => "0001011110010100000100",
			4146 => "0000000100000011100101",
			4147 => "0000000100000011100101",
			4148 => "0001011101101100000100",
			4149 => "0000000100000011100101",
			4150 => "0001011010001100000100",
			4151 => "0000000100000011100101",
			4152 => "0000000100000011100101",
			4153 => "0010001001000101001000",
			4154 => "0011100100000000100100",
			4155 => "0000111011000000100000",
			4156 => "0011100010001100011000",
			4157 => "0000010110010000001100",
			4158 => "0000100110101100001000",
			4159 => "0011011011101100000100",
			4160 => "0000000100000111000001",
			4161 => "0000000100000111000001",
			4162 => "0000000100000111000001",
			4163 => "0010111010100100001000",
			4164 => "0000011001100000000100",
			4165 => "0000000100000111000001",
			4166 => "0000000100000111000001",
			4167 => "0000000100000111000001",
			4168 => "0000000001111000000100",
			4169 => "0000000100000111000001",
			4170 => "0000000100000111000001",
			4171 => "0000000100000111000001",
			4172 => "0001010011000100001100",
			4173 => "0000011000011000000100",
			4174 => "1111111100000111000001",
			4175 => "0001111100110000000100",
			4176 => "0000000100000111000001",
			4177 => "0000000100000111000001",
			4178 => "0010101100110100010100",
			4179 => "0001001110111000010000",
			4180 => "0010011010000100001000",
			4181 => "0011100010011100000100",
			4182 => "0000000100000111000001",
			4183 => "0000000100000111000001",
			4184 => "0000100111010000000100",
			4185 => "0000000100000111000001",
			4186 => "0000000100000111000001",
			4187 => "0000000100000111000001",
			4188 => "0000000100000111000001",
			4189 => "0000100100001000010100",
			4190 => "0011010101011100001000",
			4191 => "0001010101011100000100",
			4192 => "0000000100000111000001",
			4193 => "0000001100000111000001",
			4194 => "0001111100010000001000",
			4195 => "0001101100001100000100",
			4196 => "0000000100000111000001",
			4197 => "0000000100000111000001",
			4198 => "0000000100000111000001",
			4199 => "0001011001010100010000",
			4200 => "0001011100010000001100",
			4201 => "0001111000101000000100",
			4202 => "0000000100000111000001",
			4203 => "0000110011100100000100",
			4204 => "0000000100000111000001",
			4205 => "0000000100000111000001",
			4206 => "0000000100000111000001",
			4207 => "0000000100000111000001",
			4208 => "0000000010010000101100",
			4209 => "0001000011110100101000",
			4210 => "0001000110011100100000",
			4211 => "0010110111011100011000",
			4212 => "0011011011101100001100",
			4213 => "0011000110110100000100",
			4214 => "0000000100001010010101",
			4215 => "0010001111111100000100",
			4216 => "0000000100001010010101",
			4217 => "0000000100001010010101",
			4218 => "0001100011000100001000",
			4219 => "0011101000000100000100",
			4220 => "0000000100001010010101",
			4221 => "0000000100001010010101",
			4222 => "0000000100001010010101",
			4223 => "0000010011010000000100",
			4224 => "0000000100001010010101",
			4225 => "0000000100001010010101",
			4226 => "0011101111100000000100",
			4227 => "0000000100001010010101",
			4228 => "0000000100001010010101",
			4229 => "0000000100001010010101",
			4230 => "0011101010011000010100",
			4231 => "0000010110001100010000",
			4232 => "0010110101010100001000",
			4233 => "0001001110111000000100",
			4234 => "0000000100001010010101",
			4235 => "0000000100001010010101",
			4236 => "0000001100111100000100",
			4237 => "0000000100001010010101",
			4238 => "0000000100001010010101",
			4239 => "0000000100001010010101",
			4240 => "0001100011010100010000",
			4241 => "0011110101110100001000",
			4242 => "0011110010001000000100",
			4243 => "0000000100001010010101",
			4244 => "0000000100001010010101",
			4245 => "0011001001001000000100",
			4246 => "0000000100001010010101",
			4247 => "0000000100001010010101",
			4248 => "0001111101001000010000",
			4249 => "0001011100010000000100",
			4250 => "0000000100001010010101",
			4251 => "0011011011101100001000",
			4252 => "0011010110001100000100",
			4253 => "0000000100001010010101",
			4254 => "0000000100001010010101",
			4255 => "0000000100001010010101",
			4256 => "0001011111011000001000",
			4257 => "0010111110011000000100",
			4258 => "0000000100001010010101",
			4259 => "0000000100001010010101",
			4260 => "0000000100001010010101",
			4261 => "0011011011101100011100",
			4262 => "0000001110100100010000",
			4263 => "0001010110001100001000",
			4264 => "0000101100010000000100",
			4265 => "0000000100001101100001",
			4266 => "0000000100001101100001",
			4267 => "0011010110110100000100",
			4268 => "0000000100001101100001",
			4269 => "0000000100001101100001",
			4270 => "0001100100010000000100",
			4271 => "0000000100001101100001",
			4272 => "0000000011111000000100",
			4273 => "0000000100001101100001",
			4274 => "0000000100001101100001",
			4275 => "0011010101011101000000",
			4276 => "0010001111111100010100",
			4277 => "0011010111011100010000",
			4278 => "0010011010000100001100",
			4279 => "0001001100010000001000",
			4280 => "0001110011000000000100",
			4281 => "0000000100001101100001",
			4282 => "0000000100001101100001",
			4283 => "0000000100001101100001",
			4284 => "0000000100001101100001",
			4285 => "0000000100001101100001",
			4286 => "0001111000000000010100",
			4287 => "0000111101001000010000",
			4288 => "0011000101010100001000",
			4289 => "0001001001000100000100",
			4290 => "0000000100001101100001",
			4291 => "0000000100001101100001",
			4292 => "0001100011110100000100",
			4293 => "0000000100001101100001",
			4294 => "0000000100001101100001",
			4295 => "0000000100001101100001",
			4296 => "0000101000010100001000",
			4297 => "0001101010100000000100",
			4298 => "0000000100001101100001",
			4299 => "0000000100001101100001",
			4300 => "0011101010011000001000",
			4301 => "0010110101010100000100",
			4302 => "0000000100001101100001",
			4303 => "0000000100001101100001",
			4304 => "0010001111001000000100",
			4305 => "0000000100001101100001",
			4306 => "0000000100001101100001",
			4307 => "0001111100010000001000",
			4308 => "0001101110001100000100",
			4309 => "0000000100001101100001",
			4310 => "0000000100001101100001",
			4311 => "0000000100001101100001",
			4312 => "0000000000001101000000",
			4313 => "0011101010100000101100",
			4314 => "0010110110001100001000",
			4315 => "0000001110010100000100",
			4316 => "0000000100010001010101",
			4317 => "0000000100010001010101",
			4318 => "0000011000011000010000",
			4319 => "0001001100101100001100",
			4320 => "0010001001000100000100",
			4321 => "0000000100010001010101",
			4322 => "0010001111001000000100",
			4323 => "0000000100010001010101",
			4324 => "0000000100010001010101",
			4325 => "0000000100010001010101",
			4326 => "0001000111011100001100",
			4327 => "0001010101010100000100",
			4328 => "0000000100010001010101",
			4329 => "0001011001001000000100",
			4330 => "0000000100010001010101",
			4331 => "0000000100010001010101",
			4332 => "0011001001001000000100",
			4333 => "0000000100010001010101",
			4334 => "0000000100010001010101",
			4335 => "0001001111011000001000",
			4336 => "0011001010100100000100",
			4337 => "0000000100010001010101",
			4338 => "0000000100010001010101",
			4339 => "0001011111100000001000",
			4340 => "0001000110011100000100",
			4341 => "0000000100010001010101",
			4342 => "0000000100010001010101",
			4343 => "0000000100010001010101",
			4344 => "0011101010011000011100",
			4345 => "0001001110001100010100",
			4346 => "0000010110001100010000",
			4347 => "0010000011010000000100",
			4348 => "0000000100010001010101",
			4349 => "0001111001010100001000",
			4350 => "0011001001001000000100",
			4351 => "0000000100010001010101",
			4352 => "0000000100010001010101",
			4353 => "0000000100010001010101",
			4354 => "0000000100010001010101",
			4355 => "0001111000101000000100",
			4356 => "0000000100010001010101",
			4357 => "0000000100010001010101",
			4358 => "0000001011011000001100",
			4359 => "0011111110100000000100",
			4360 => "0000000100010001010101",
			4361 => "0001111001010000000100",
			4362 => "0000000100010001010101",
			4363 => "0000000100010001010101",
			4364 => "0001111101001000010000",
			4365 => "0000111111101000001100",
			4366 => "0001110110101100000100",
			4367 => "0000000100010001010101",
			4368 => "0000010111110000000100",
			4369 => "0000000100010001010101",
			4370 => "0000000100010001010101",
			4371 => "0000000100010001010101",
			4372 => "0000000100010001010101",
			4373 => "0011011010100101000000",
			4374 => "0000111011000000101100",
			4375 => "0001011110001100100100",
			4376 => "0010111110011000010000",
			4377 => "0010000011010000000100",
			4378 => "0000000100010101100001",
			4379 => "0001000001100100000100",
			4380 => "0000000100010101100001",
			4381 => "0011101100100000000100",
			4382 => "0000000100010101100001",
			4383 => "0000000100010101100001",
			4384 => "0011011011101100000100",
			4385 => "0000000100010101100001",
			4386 => "0001111000111000001000",
			4387 => "0000011000011000000100",
			4388 => "0000000100010101100001",
			4389 => "0000000100010101100001",
			4390 => "0011101110111100000100",
			4391 => "0000000100010101100001",
			4392 => "0000000100010101100001",
			4393 => "0010001111111100000100",
			4394 => "0000000100010101100001",
			4395 => "0000000100010101100001",
			4396 => "0010110101010100001000",
			4397 => "0001110110101100000100",
			4398 => "0000000100010101100001",
			4399 => "0000000100010101100001",
			4400 => "0001000001011000000100",
			4401 => "0000000100010101100001",
			4402 => "0011001001001000000100",
			4403 => "0000000100010101100001",
			4404 => "0000000100010101100001",
			4405 => "0001111100010000100000",
			4406 => "0011001100101000010000",
			4407 => "0000110101111000001000",
			4408 => "0001111101101000000100",
			4409 => "0000000100010101100001",
			4410 => "0000000100010101100001",
			4411 => "0011100010001100000100",
			4412 => "0000000100010101100001",
			4413 => "0000000100010101100001",
			4414 => "0000001010101100001100",
			4415 => "0010010011000000000100",
			4416 => "0000000100010101100001",
			4417 => "0010010101111000000100",
			4418 => "0000000100010101100001",
			4419 => "0000000100010101100001",
			4420 => "0000000100010101100001",
			4421 => "0001001110111000011000",
			4422 => "0011110100101000010000",
			4423 => "0000000010010000001000",
			4424 => "0000000100011100000100",
			4425 => "0000000100010101100001",
			4426 => "0000000100010101100001",
			4427 => "0001101111000100000100",
			4428 => "0000000100010101100001",
			4429 => "0000000100010101100001",
			4430 => "0001111001010000000100",
			4431 => "0000000100010101100001",
			4432 => "0000000100010101100001",
			4433 => "0010100001101000000100",
			4434 => "0000000100010101100001",
			4435 => "0001000010001100000100",
			4436 => "0000000100010101100001",
			4437 => "0001001111100100000100",
			4438 => "0000000100010101100001",
			4439 => "0000000100010101100001",
			4440 => "0010101100001101011000",
			4441 => "0001001100101100111100",
			4442 => "0010110111011100101100",
			4443 => "0011011011101100010100",
			4444 => "0000101001111100001000",
			4445 => "0011001110011000000100",
			4446 => "0000000100011000101101",
			4447 => "0000000100011000101101",
			4448 => "0001100100010000000100",
			4449 => "0000000100011000101101",
			4450 => "0011111010101100000100",
			4451 => "0000000100011000101101",
			4452 => "0000000100011000101101",
			4453 => "0011010011010000010000",
			4454 => "0001100010110000001000",
			4455 => "0000010110010000000100",
			4456 => "0000000100011000101101",
			4457 => "0000000100011000101101",
			4458 => "0000111000101000000100",
			4459 => "0000000100011000101101",
			4460 => "0000000100011000101101",
			4461 => "0000001011101000000100",
			4462 => "0000000100011000101101",
			4463 => "0000000100011000101101",
			4464 => "0001001111101000001000",
			4465 => "0010000101011100000100",
			4466 => "0000000100011000101101",
			4467 => "0000000100011000101101",
			4468 => "0001000100101100000100",
			4469 => "0000000100011000101101",
			4470 => "0000000100011000101101",
			4471 => "0011000101010100000100",
			4472 => "0000000100011000101101",
			4473 => "0000000000001100001000",
			4474 => "0010101110111000000100",
			4475 => "0000000100011000101101",
			4476 => "0000000100011000101101",
			4477 => "0011100000100000001000",
			4478 => "0011000101011100000100",
			4479 => "0000000100011000101101",
			4480 => "0000000100011000101101",
			4481 => "0010010101111000000100",
			4482 => "0000000100011000101101",
			4483 => "0000000100011000101101",
			4484 => "0011101001110000001000",
			4485 => "0000000010111100000100",
			4486 => "0000000100011000101101",
			4487 => "0000000100011000101101",
			4488 => "0000010110010000000100",
			4489 => "0000000100011000101101",
			4490 => "0000000100011000101101",
			4491 => "0000001011011101001100",
			4492 => "0011101010100000110100",
			4493 => "0000000111001000100100",
			4494 => "0010010110000000011000",
			4495 => "0001010110001100001100",
			4496 => "0001000000011000000100",
			4497 => "0000000100011100101001",
			4498 => "0011011011101100000100",
			4499 => "0000000100011100101001",
			4500 => "0000000100011100101001",
			4501 => "0011000101011100001000",
			4502 => "0000010001110000000100",
			4503 => "0000000100011100101001",
			4504 => "0000000100011100101001",
			4505 => "0000000100011100101001",
			4506 => "0000010011010000001000",
			4507 => "0011011011101100000100",
			4508 => "0000000100011100101001",
			4509 => "0000000100011100101001",
			4510 => "0000000100011100101001",
			4511 => "0000010001100100001000",
			4512 => "0011100010001100000100",
			4513 => "0000000100011100101001",
			4514 => "0000000100011100101001",
			4515 => "0011100010111000000100",
			4516 => "0000000100011100101001",
			4517 => "0000000100011100101001",
			4518 => "0010001111011000010100",
			4519 => "0010001111111100001100",
			4520 => "0000111011000000001000",
			4521 => "0011110011010100000100",
			4522 => "0000000100011100101001",
			4523 => "0000000100011100101001",
			4524 => "0000000100011100101001",
			4525 => "0011001100101000000100",
			4526 => "0000000100011100101001",
			4527 => "0000000100011100101001",
			4528 => "0000000100011100101001",
			4529 => "0001100000110100010100",
			4530 => "0000010110001100010000",
			4531 => "0011100000010100001100",
			4532 => "0011010111011100000100",
			4533 => "0000000100011100101001",
			4534 => "0001011101101100000100",
			4535 => "0000000100011100101001",
			4536 => "0000000100011100101001",
			4537 => "0000000100011100101001",
			4538 => "0000000100011100101001",
			4539 => "0001001111101000011000",
			4540 => "0001111100010000001000",
			4541 => "0010101000111000000100",
			4542 => "0000000100011100101001",
			4543 => "0000000100011100101001",
			4544 => "0010101000000000000100",
			4545 => "0000000100011100101001",
			4546 => "0000010111110000001000",
			4547 => "0000011001100100000100",
			4548 => "0000000100011100101001",
			4549 => "0000000100011100101001",
			4550 => "0000000100011100101001",
			4551 => "0011001001001000000100",
			4552 => "0000000100011100101001",
			4553 => "0000000100011100101001",
			4554 => "0000100100011100110000",
			4555 => "0011100001101000100000",
			4556 => "0001110111011100000100",
			4557 => "0000000100100000011101",
			4558 => "0010001001000100010000",
			4559 => "0000010111100100000100",
			4560 => "0000000100100000011101",
			4561 => "0000011001100000001000",
			4562 => "0000011000011000000100",
			4563 => "0000000100100000011101",
			4564 => "0000000100100000011101",
			4565 => "0000000100100000011101",
			4566 => "0001010110000000000100",
			4567 => "0000000100100000011101",
			4568 => "0011001100101000000100",
			4569 => "0000000100100000011101",
			4570 => "0000000100100000011101",
			4571 => "0000010110001100001100",
			4572 => "0010000101011100000100",
			4573 => "0000000100100000011101",
			4574 => "0001111000000100000100",
			4575 => "0000000100100000011101",
			4576 => "0000000100100000011101",
			4577 => "0000000100100000011101",
			4578 => "0011101111100100011000",
			4579 => "0011011010100100001100",
			4580 => "0000111011000000001000",
			4581 => "0000010001110000000100",
			4582 => "0000000100100000011101",
			4583 => "0000000100100000011101",
			4584 => "0000000100100000011101",
			4585 => "0011001100101000000100",
			4586 => "0000000100100000011101",
			4587 => "0010100000111100000100",
			4588 => "0000000100100000011101",
			4589 => "0000000100100000011101",
			4590 => "0000101110000100001100",
			4591 => "0000111000101000001000",
			4592 => "0011101110111100000100",
			4593 => "0000000100100000011101",
			4594 => "0000000100100000011101",
			4595 => "0000000100100000011101",
			4596 => "0001111100010000001100",
			4597 => "0010101000111000000100",
			4598 => "0000000100100000011101",
			4599 => "0010101011111000000100",
			4600 => "0000000100100000011101",
			4601 => "0000000100100000011101",
			4602 => "0000010000011000010000",
			4603 => "0000100011111100001000",
			4604 => "0001101100100000000100",
			4605 => "0000000100100000011101",
			4606 => "0000000100100000011101",
			4607 => "0000111011111000000100",
			4608 => "0000000100100000011101",
			4609 => "0000000100100000011101",
			4610 => "0010101000000000000100",
			4611 => "0000000100100000011101",
			4612 => "0001000001111100000100",
			4613 => "0000000100100000011101",
			4614 => "0000000100100000011101",
			4615 => "0000001100111100111000",
			4616 => "0000001000000100000100",
			4617 => "1111111100100011000001",
			4618 => "0000010001110000010100",
			4619 => "0000011001100100000100",
			4620 => "1111111100100011000001",
			4621 => "0000001010101100001100",
			4622 => "0011100010001100001000",
			4623 => "0000000001011100000100",
			4624 => "0000001100100011000001",
			4625 => "1111111100100011000001",
			4626 => "0000001100100011000001",
			4627 => "1111111100100011000001",
			4628 => "0010111100101000011000",
			4629 => "0011001010100100001100",
			4630 => "0010000101011100000100",
			4631 => "0000001100100011000001",
			4632 => "0011101010011100000100",
			4633 => "0000001100100011000001",
			4634 => "0000010100100011000001",
			4635 => "0001011000000100000100",
			4636 => "1111111100100011000001",
			4637 => "0011011011101100000100",
			4638 => "0000000100100011000001",
			4639 => "0000001100100011000001",
			4640 => "0001001000111000000100",
			4641 => "1111111100100011000001",
			4642 => "0000001100100011000001",
			4643 => "0011101110111100011000",
			4644 => "0011110010011000000100",
			4645 => "1111111100100011000001",
			4646 => "0001111000101000010000",
			4647 => "0011101010011000000100",
			4648 => "1111111100100011000001",
			4649 => "0010110011010000000100",
			4650 => "0000000100100011000001",
			4651 => "0011100000010100000100",
			4652 => "0000001100100011000001",
			4653 => "0000010100100011000001",
			4654 => "1111111100100011000001",
			4655 => "1111111100100011000001",
			4656 => "0011011011101100100100",
			4657 => "0000111011000000100000",
			4658 => "0000111011111000011100",
			4659 => "0011000110110100001000",
			4660 => "0000001010011100000100",
			4661 => "0000000100100110100101",
			4662 => "0000000100100110100101",
			4663 => "0001101110001100001100",
			4664 => "0011101001010100000100",
			4665 => "0000000100100110100101",
			4666 => "0000101101000100000100",
			4667 => "0000000100100110100101",
			4668 => "0000000100100110100101",
			4669 => "0000011000011000000100",
			4670 => "0000000100100110100101",
			4671 => "0000000100100110100101",
			4672 => "0000000100100110100101",
			4673 => "1111111100100110100101",
			4674 => "0000000000001100101100",
			4675 => "0011101101111100100000",
			4676 => "0000011000011000010100",
			4677 => "0010110111011100001000",
			4678 => "0010101100010000000100",
			4679 => "0000000100100110100101",
			4680 => "0000000100100110100101",
			4681 => "0000010111110000001000",
			4682 => "0000010001110000000100",
			4683 => "0000000100100110100101",
			4684 => "0000000100100110100101",
			4685 => "1111111100100110100101",
			4686 => "0011001001001000001000",
			4687 => "0001010011010000000100",
			4688 => "0000000100100110100101",
			4689 => "0000000100100110100101",
			4690 => "0000000100100110100101",
			4691 => "0001011011000000000100",
			4692 => "0000000100100110100101",
			4693 => "0001110110101100000100",
			4694 => "0000001100100110100101",
			4695 => "0000000100100110100101",
			4696 => "0001101010011000001000",
			4697 => "0010101010011100000100",
			4698 => "1111111100100110100101",
			4699 => "0000000100100110100101",
			4700 => "0010010101101100001100",
			4701 => "0001000101010100001000",
			4702 => "0011001010100100000100",
			4703 => "0000000100100110100101",
			4704 => "0000000100100110100101",
			4705 => "0000000100100110100101",
			4706 => "0001110001010000001100",
			4707 => "0010011001000100000100",
			4708 => "0000000100100110100101",
			4709 => "0001001000100000000100",
			4710 => "0000000100100110100101",
			4711 => "0000000100100110100101",
			4712 => "0000000100100110100101",
			4713 => "0000001100000100101100",
			4714 => "0010000011010000000100",
			4715 => "0000000100101010001001",
			4716 => "0001100100000000100100",
			4717 => "0000000111001000011000",
			4718 => "0011000101011100010000",
			4719 => "0001010110001100001000",
			4720 => "0010100110010000000100",
			4721 => "0000000100101010001001",
			4722 => "0000000100101010001001",
			4723 => "0000010001110000000100",
			4724 => "0000000100101010001001",
			4725 => "0000000100101010001001",
			4726 => "0000010011010000000100",
			4727 => "0000000100101010001001",
			4728 => "0000000100101010001001",
			4729 => "0000011000011000001000",
			4730 => "0000000011101000000100",
			4731 => "0000000100101010001001",
			4732 => "0000000100101010001001",
			4733 => "0000000100101010001001",
			4734 => "0000000100101010001001",
			4735 => "0001001110111000110100",
			4736 => "0011101010011000010000",
			4737 => "0011010111011100001000",
			4738 => "0001011111100000000100",
			4739 => "0000000100101010001001",
			4740 => "0000000100101010001001",
			4741 => "0001011001011000000100",
			4742 => "0000000100101010001001",
			4743 => "0000000100101010001001",
			4744 => "0000110011001000010000",
			4745 => "0001011000111000001100",
			4746 => "0011100010011000000100",
			4747 => "0000000100101010001001",
			4748 => "0000001000100100000100",
			4749 => "0000000100101010001001",
			4750 => "0000000100101010001001",
			4751 => "0000000100101010001001",
			4752 => "0011010110001100001000",
			4753 => "0001101110010000000100",
			4754 => "0000000100101010001001",
			4755 => "0000000100101010001001",
			4756 => "0001000000111100001000",
			4757 => "0001001111101000000100",
			4758 => "0000000100101010001001",
			4759 => "0000000100101010001001",
			4760 => "0000000100101010001001",
			4761 => "0010100001101000001000",
			4762 => "0000111110111000000100",
			4763 => "0000000100101010001001",
			4764 => "0000000100101010001001",
			4765 => "0001000010001100000100",
			4766 => "0000000100101010001001",
			4767 => "0001001111100100000100",
			4768 => "0000000100101010001001",
			4769 => "0000000100101010001001",
			4770 => "0001000010111001001000",
			4771 => "0001000011110101000000",
			4772 => "0000111110111000110100",
			4773 => "0001001100101100100000",
			4774 => "0010110111011100010000",
			4775 => "0010001111111100001000",
			4776 => "0011000110110100000100",
			4777 => "0000000100101100111101",
			4778 => "0000000100101100111101",
			4779 => "0010101001011000000100",
			4780 => "0000000100101100111101",
			4781 => "1111111100101100111101",
			4782 => "0001001111101000001000",
			4783 => "0010000101011100000100",
			4784 => "0000000100101100111101",
			4785 => "1111111100101100111101",
			4786 => "0000111011000000000100",
			4787 => "0000000100101100111101",
			4788 => "0000000100101100111101",
			4789 => "0001001011000000000100",
			4790 => "0000001100101100111101",
			4791 => "0000000000001100001000",
			4792 => "0011111010110100000100",
			4793 => "0000000100101100111101",
			4794 => "0000001100101100111101",
			4795 => "0011100010011100000100",
			4796 => "1111111100101100111101",
			4797 => "0000000100101100111101",
			4798 => "0011001001001000000100",
			4799 => "1111111100101100111101",
			4800 => "0011101111000000000100",
			4801 => "0000000100101100111101",
			4802 => "0000000100101100111101",
			4803 => "0010000101101100000100",
			4804 => "1111111100101100111101",
			4805 => "0000000100101100111101",
			4806 => "0011011010100100000100",
			4807 => "0000000100101100111101",
			4808 => "0001011111111000000100",
			4809 => "0000001100101100111101",
			4810 => "0011111110111100001000",
			4811 => "0001100010010100000100",
			4812 => "0000000100101100111101",
			4813 => "0000000100101100111101",
			4814 => "0000000100101100111101",
			4815 => "0000000111001000011000",
			4816 => "0001010110001100001000",
			4817 => "0001110101010100000100",
			4818 => "0000000100110000001001",
			4819 => "0000000100110000001001",
			4820 => "0011000101011100001000",
			4821 => "0010001001001100000100",
			4822 => "0000000100110000001001",
			4823 => "0000000100110000001001",
			4824 => "0000010011010000000100",
			4825 => "0000000100110000001001",
			4826 => "0000000100110000001001",
			4827 => "0011100010001100001000",
			4828 => "0010001111001000000100",
			4829 => "0000000100110000001001",
			4830 => "0000000100110000001001",
			4831 => "0001010011000100101000",
			4832 => "0000011000011000001100",
			4833 => "0001010101111000001000",
			4834 => "0001010011000000000100",
			4835 => "0000000100110000001001",
			4836 => "0000000100110000001001",
			4837 => "1111111100110000001001",
			4838 => "0011010011010000001100",
			4839 => "0001010101111000000100",
			4840 => "0000000100110000001001",
			4841 => "0010101001010100000100",
			4842 => "0000001100110000001001",
			4843 => "0000000100110000001001",
			4844 => "0000001011101000001000",
			4845 => "0011111010011000000100",
			4846 => "0000000100110000001001",
			4847 => "0000000100110000001001",
			4848 => "0000100111000100000100",
			4849 => "0000000100110000001001",
			4850 => "0000000100110000001001",
			4851 => "0000001100000100000100",
			4852 => "0000000100110000001001",
			4853 => "0001100000110100010000",
			4854 => "0000001100111100001000",
			4855 => "0011101001111100000100",
			4856 => "0000000100110000001001",
			4857 => "0000000100110000001001",
			4858 => "0010001111001000000100",
			4859 => "0000000100110000001001",
			4860 => "0000000100110000001001",
			4861 => "0010001111001000001000",
			4862 => "0011001001001000000100",
			4863 => "0000000100110000001001",
			4864 => "0000000100110000001001",
			4865 => "0000000100110000001001",
			4866 => "0011101110111101000000",
			4867 => "0011000110000000111100",
			4868 => "0010001001001100010000",
			4869 => "0010010110000000001000",
			4870 => "0001000111100100000100",
			4871 => "0000000100110010001101",
			4872 => "1111111100110010001101",
			4873 => "0010110111011100000100",
			4874 => "0000001100110010001101",
			4875 => "1111111100110010001101",
			4876 => "0011000011010000010000",
			4877 => "0000001110100000001000",
			4878 => "0001011011101100000100",
			4879 => "0000000100110010001101",
			4880 => "0000001100110010001101",
			4881 => "0011011011101100000100",
			4882 => "1111111100110010001101",
			4883 => "0000000100110010001101",
			4884 => "0001011001011000010000",
			4885 => "0010110011010000001000",
			4886 => "0000011000011000000100",
			4887 => "1111111100110010001101",
			4888 => "0000000100110010001101",
			4889 => "0001011111101000000100",
			4890 => "1111111100110010001101",
			4891 => "0000000100110010001101",
			4892 => "0011100010001100000100",
			4893 => "0000000100110010001101",
			4894 => "0000001100000100000100",
			4895 => "0000001100110010001101",
			4896 => "0000000100110010001101",
			4897 => "1111111100110010001101",
			4898 => "1111111100110010001101",
			4899 => "0000000010010001000000",
			4900 => "0011101010100000110000",
			4901 => "0000000111001000011100",
			4902 => "0001010110001100001000",
			4903 => "0001110111011100000100",
			4904 => "0000000100110110010001",
			4905 => "0000000100110110010001",
			4906 => "0011001100101000010000",
			4907 => "0011100011000100001000",
			4908 => "0011001010100100000100",
			4909 => "0000000100110110010001",
			4910 => "0000000100110110010001",
			4911 => "0010010101101100000100",
			4912 => "0000000100110110010001",
			4913 => "0000001100110110010001",
			4914 => "0000000100110110010001",
			4915 => "0011011010100100001100",
			4916 => "0001010010111000001000",
			4917 => "0001011010011100000100",
			4918 => "0000000100110110010001",
			4919 => "0000000100110110010001",
			4920 => "1111111100110110010001",
			4921 => "0011111010100000000100",
			4922 => "0000000100110110010001",
			4923 => "0000000100110110010001",
			4924 => "0001000110011100001100",
			4925 => "0010100100101100001000",
			4926 => "0011011011101100000100",
			4927 => "0000000100110110010001",
			4928 => "0000000100110110010001",
			4929 => "0000000100110110010001",
			4930 => "0000001100110110010001",
			4931 => "0001100100100100001100",
			4932 => "0010011111011000000100",
			4933 => "1111111100110110010001",
			4934 => "0010001111011000000100",
			4935 => "0000000100110110010001",
			4936 => "0000000100110110010001",
			4937 => "0001101111000100011000",
			4938 => "0011011110011000001000",
			4939 => "0001010111010100000100",
			4940 => "0000000100110110010001",
			4941 => "0000000100110110010001",
			4942 => "0010101100110100000100",
			4943 => "0000001100110110010001",
			4944 => "0001101101000100000100",
			4945 => "0000000100110110010001",
			4946 => "0011100100100100000100",
			4947 => "0000000100110110010001",
			4948 => "0000000100110110010001",
			4949 => "0011101010011000000100",
			4950 => "1111111100110110010001",
			4951 => "0001111101001000001100",
			4952 => "0001011000111000000100",
			4953 => "0000000100110110010001",
			4954 => "0000100111000100000100",
			4955 => "0000000100110110010001",
			4956 => "0000000100110110010001",
			4957 => "0001000001011000001000",
			4958 => "0011001110011000000100",
			4959 => "0000000100110110010001",
			4960 => "1111111100110110010001",
			4961 => "0011110011101100000100",
			4962 => "0000000100110110010001",
			4963 => "0000000100110110010001",
			4964 => "0000001100000100101100",
			4965 => "0010000011010000000100",
			4966 => "0000000100111001011101",
			4967 => "0001000110011100100100",
			4968 => "0011000011010000001100",
			4969 => "0001000001100100000100",
			4970 => "0000000100111001011101",
			4971 => "0000100010110000000100",
			4972 => "0000000100111001011101",
			4973 => "0000000100111001011101",
			4974 => "0011011010100100001100",
			4975 => "0000011000011000001000",
			4976 => "0010011010000100000100",
			4977 => "0000000100111001011101",
			4978 => "0000000100111001011101",
			4979 => "0000000100111001011101",
			4980 => "0001011000101000001000",
			4981 => "0010010110000000000100",
			4982 => "0000000100111001011101",
			4983 => "0000000100111001011101",
			4984 => "0000000100111001011101",
			4985 => "0000000100111001011101",
			4986 => "0001001000000100010100",
			4987 => "0011101010011000000100",
			4988 => "0000000100111001011101",
			4989 => "0011111101100100000100",
			4990 => "0000000100111001011101",
			4991 => "0011000111011100000100",
			4992 => "0000000100111001011101",
			4993 => "0000110011001000000100",
			4994 => "0000000100111001011101",
			4995 => "0000000100111001011101",
			4996 => "0011101010100000000100",
			4997 => "0000000100111001011101",
			4998 => "0000000000001100001000",
			4999 => "0010101110111000000100",
			5000 => "0000000100111001011101",
			5001 => "0000000100111001011101",
			5002 => "0001001110111000001100",
			5003 => "0011100010011100000100",
			5004 => "0000000100111001011101",
			5005 => "0000110000111100000100",
			5006 => "0000000100111001011101",
			5007 => "0000000100111001011101",
			5008 => "0011011010100100001000",
			5009 => "0010000101011100000100",
			5010 => "0000000100111001011101",
			5011 => "0000000100111001011101",
			5012 => "0001111000101000000100",
			5013 => "0000000100111001011101",
			5014 => "0000000100111001011101",
			5015 => "0011011011101100100100",
			5016 => "0000111011000000100000",
			5017 => "0000111011111000011100",
			5018 => "0000001110100100010100",
			5019 => "0001010110001100001000",
			5020 => "0001001000011000000100",
			5021 => "0000000100111100100001",
			5022 => "0000000100111100100001",
			5023 => "0011000011010000001000",
			5024 => "0010001001001100000100",
			5025 => "0000000100111100100001",
			5026 => "0000001100111100100001",
			5027 => "0000000100111100100001",
			5028 => "0010101011000000000100",
			5029 => "1111111100111100100001",
			5030 => "0000000100111100100001",
			5031 => "0000000100111100100001",
			5032 => "1111111100111100100001",
			5033 => "0001110001010000111100",
			5034 => "0010010011000000100100",
			5035 => "0001010001010100011100",
			5036 => "0011111110000000001100",
			5037 => "0011101001101100001000",
			5038 => "0010110111011100000100",
			5039 => "0000000100111100100001",
			5040 => "1111111100111100100001",
			5041 => "0000001100111100100001",
			5042 => "0011101111000100001000",
			5043 => "0000111100101100000100",
			5044 => "0000000100111100100001",
			5045 => "0000000100111100100001",
			5046 => "0001100110111000000100",
			5047 => "0000000100111100100001",
			5048 => "0000000100111100100001",
			5049 => "0000110011110100000100",
			5050 => "0000000100111100100001",
			5051 => "0000000100111100100001",
			5052 => "0010101110111000010000",
			5053 => "0001110110101100001100",
			5054 => "0000000111101000001000",
			5055 => "0010101001010100000100",
			5056 => "0000000100111100100001",
			5057 => "0000000100111100100001",
			5058 => "0000000100111100100001",
			5059 => "0000000100111100100001",
			5060 => "0010100001101000000100",
			5061 => "0000001100111100100001",
			5062 => "0000000100111100100001",
			5063 => "0000000100111100100001",
			5064 => "0011101110111100111100",
			5065 => "0001000010111000110100",
			5066 => "0001001100001100110000",
			5067 => "0000000000001100011100",
			5068 => "0011101101111100010000",
			5069 => "0000001100000100001000",
			5070 => "0011001100101000000100",
			5071 => "0000000100111110011101",
			5072 => "1111111100111110011101",
			5073 => "0011010111011100000100",
			5074 => "1111111100111110011101",
			5075 => "0000000100111110011101",
			5076 => "0001000110011100001000",
			5077 => "0011111010011000000100",
			5078 => "0000001100111110011101",
			5079 => "0000000100111110011101",
			5080 => "0000001100111110011101",
			5081 => "0011100010011100000100",
			5082 => "1111111100111110011101",
			5083 => "0000111110111000001000",
			5084 => "0001011000111000000100",
			5085 => "1111111100111110011101",
			5086 => "0000000100111110011101",
			5087 => "0000000101000100000100",
			5088 => "0000000100111110011101",
			5089 => "1111111100111110011101",
			5090 => "1111111100111110011101",
			5091 => "0000110001101000000100",
			5092 => "0000001100111110011101",
			5093 => "1111111100111110011101",
			5094 => "1111111100111110011101",
			5095 => "0010001111111100100100",
			5096 => "0011000110110100000100",
			5097 => "0000000101000001110001",
			5098 => "0011111100000100011000",
			5099 => "0001011110001100000100",
			5100 => "0000000101000001110001",
			5101 => "0001010001111100001000",
			5102 => "0000001110101100000100",
			5103 => "0000000101000001110001",
			5104 => "0000000101000001110001",
			5105 => "0000111010011100000100",
			5106 => "0000000101000001110001",
			5107 => "0000110010111000000100",
			5108 => "0000000101000001110001",
			5109 => "0000000101000001110001",
			5110 => "0001001000111000000100",
			5111 => "0000000101000001110001",
			5112 => "0000000101000001110001",
			5113 => "0001101111010101000000",
			5114 => "0011010101011100110100",
			5115 => "0001111000000000011000",
			5116 => "0010111010100100001000",
			5117 => "0001010100101100000100",
			5118 => "0000000101000001110001",
			5119 => "0000000101000001110001",
			5120 => "0011011010100100001000",
			5121 => "0010110101010100000100",
			5122 => "0000000101000001110001",
			5123 => "0000000101000001110001",
			5124 => "0010010110000000000100",
			5125 => "0000000101000001110001",
			5126 => "0000000101000001110001",
			5127 => "0010110101011100001100",
			5128 => "0011011011101100000100",
			5129 => "0000000101000001110001",
			5130 => "0001010101111000000100",
			5131 => "0000000101000001110001",
			5132 => "0000000101000001110001",
			5133 => "0000101101010100001000",
			5134 => "0000100001100000000100",
			5135 => "0000000101000001110001",
			5136 => "0000000101000001110001",
			5137 => "0011101001110000000100",
			5138 => "0000000101000001110001",
			5139 => "0000000101000001110001",
			5140 => "0001111100010000001000",
			5141 => "0001101110001100000100",
			5142 => "0000000101000001110001",
			5143 => "0000000101000001110001",
			5144 => "0000000101000001110001",
			5145 => "0000010000011000000100",
			5146 => "0000000101000001110001",
			5147 => "0000000101000001110001",
			5148 => "0001101111010101100100",
			5149 => "0010001111111100100000",
			5150 => "0000001101001100011100",
			5151 => "0001011110001100001100",
			5152 => "0011000110110100000100",
			5153 => "0000000101000101001101",
			5154 => "0000010111100100000100",
			5155 => "1111111101000101001101",
			5156 => "0000000101000101001101",
			5157 => "0001010001111100001000",
			5158 => "0000000000010000000100",
			5159 => "0000001101000101001101",
			5160 => "0000000101000101001101",
			5161 => "0011110010010100000100",
			5162 => "1111111101000101001101",
			5163 => "0000000101000101001101",
			5164 => "1111111101000101001101",
			5165 => "0011101001101100100100",
			5166 => "0011000011010000001000",
			5167 => "0011111010100000000100",
			5168 => "0000001101000101001101",
			5169 => "0000000101000101001101",
			5170 => "0010001111001000010000",
			5171 => "0001111000000000001000",
			5172 => "0011011010100100000100",
			5173 => "1111111101000101001101",
			5174 => "0000000101000101001101",
			5175 => "0010001001000100000100",
			5176 => "0000000101000101001101",
			5177 => "0000000101000101001101",
			5178 => "0001100011110100000100",
			5179 => "0000000101000101001101",
			5180 => "0010111001001000000100",
			5181 => "0000000101000101001101",
			5182 => "0000000101000101001101",
			5183 => "0011010101010100010100",
			5184 => "0000000100110000000100",
			5185 => "0000001101000101001101",
			5186 => "0011101111100100001000",
			5187 => "0011100101110000000100",
			5188 => "0000000101000101001101",
			5189 => "0000000101000101001101",
			5190 => "0000100000001100000100",
			5191 => "0000001101000101001101",
			5192 => "0000000101000101001101",
			5193 => "0011100010011100001000",
			5194 => "0010000011001000000100",
			5195 => "0000000101000101001101",
			5196 => "0000000101000101001101",
			5197 => "1111111101000101001101",
			5198 => "0000010111110000001000",
			5199 => "0010110011010000000100",
			5200 => "0000000101000101001101",
			5201 => "0000000101000101001101",
			5202 => "1111111101000101001101",
			5203 => "0001100100010001010000",
			5204 => "0011010101011101000100",
			5205 => "0000011000011000100100",
			5206 => "0000000111110100100000",
			5207 => "0001011110001100010000",
			5208 => "0001110011000000001000",
			5209 => "0011000111011100000100",
			5210 => "0000000101000111110001",
			5211 => "1111111101000111110001",
			5212 => "0010010101101100000100",
			5213 => "0000000101000111110001",
			5214 => "1111111101000111110001",
			5215 => "0000111011000000001000",
			5216 => "0010001111111100000100",
			5217 => "0000001101000111110001",
			5218 => "0000000101000111110001",
			5219 => "0011011110011000000100",
			5220 => "1111111101000111110001",
			5221 => "0000000101000111110001",
			5222 => "0000001101000111110001",
			5223 => "0000101000110100010100",
			5224 => "0011001100101000001100",
			5225 => "0001000001100100000100",
			5226 => "0000000101000111110001",
			5227 => "0011010110001100000100",
			5228 => "0000000101000111110001",
			5229 => "0000001101000111110001",
			5230 => "0001101001010100000100",
			5231 => "1111111101000111110001",
			5232 => "0000000101000111110001",
			5233 => "0011100010011100000100",
			5234 => "1111111101000111110001",
			5235 => "0000101011010100000100",
			5236 => "0000000101000111110001",
			5237 => "0000000101000111110001",
			5238 => "0001111100010000001000",
			5239 => "0001100011110100000100",
			5240 => "1111111101000111110001",
			5241 => "0000001101000111110001",
			5242 => "1111111101000111110001",
			5243 => "1111111101000111110001",
			5244 => "0001000010111001100000",
			5245 => "0000001100000100011100",
			5246 => "0010000011010000000100",
			5247 => "1111111101001010111101",
			5248 => "0001100100000000010000",
			5249 => "0010110110001100000100",
			5250 => "0000001101001010111101",
			5251 => "0001000110001100000100",
			5252 => "1111111101001010111101",
			5253 => "0000000111001000000100",
			5254 => "0000000101001010111101",
			5255 => "0000000101001010111101",
			5256 => "0011000101010100000100",
			5257 => "0000000101001010111101",
			5258 => "0000001101001010111101",
			5259 => "0011101111100100010100",
			5260 => "0000000000001100010000",
			5261 => "0000001010101100001100",
			5262 => "0010001111111100000100",
			5263 => "0000000101001010111101",
			5264 => "0011010111011100000100",
			5265 => "1111111101001010111101",
			5266 => "0000000101001010111101",
			5267 => "0000000101001010111101",
			5268 => "1111111101001010111101",
			5269 => "0001011001011000011000",
			5270 => "0000110011001000001100",
			5271 => "0010010101101100001000",
			5272 => "0000101100111000000100",
			5273 => "0000000101001010111101",
			5274 => "1111111101001010111101",
			5275 => "0000001101001010111101",
			5276 => "0001001001001000001000",
			5277 => "0011110100100000000100",
			5278 => "0000000101001010111101",
			5279 => "0000000101001010111101",
			5280 => "1111111101001010111101",
			5281 => "0000100111010000001100",
			5282 => "0011011110011000000100",
			5283 => "0000000101001010111101",
			5284 => "0001100100100100000100",
			5285 => "0000000101001010111101",
			5286 => "0000001101001010111101",
			5287 => "0011111110100100000100",
			5288 => "1111111101001010111101",
			5289 => "0000010110010000000100",
			5290 => "0000001101001010111101",
			5291 => "0000000101001010111101",
			5292 => "0001111000101000000100",
			5293 => "0000001101001010111101",
			5294 => "1111111101001010111101",
			5295 => "0001110001010001010100",
			5296 => "0001001100110101001100",
			5297 => "0000111011000000110000",
			5298 => "0010011101101000100000",
			5299 => "0001001000000100010000",
			5300 => "0010001111111100001000",
			5301 => "0011000110110100000100",
			5302 => "0000000101001101101001",
			5303 => "1111111101001101101001",
			5304 => "0010101101001000000100",
			5305 => "0000000101001101101001",
			5306 => "0000000101001101101001",
			5307 => "0001111000000100001000",
			5308 => "0011111010100000000100",
			5309 => "0000000101001101101001",
			5310 => "0000000101001101101001",
			5311 => "0000100111000100000100",
			5312 => "0000001101001101101001",
			5313 => "0000000101001101101001",
			5314 => "0010110111011100000100",
			5315 => "0000000101001101101001",
			5316 => "0000001000110100001000",
			5317 => "0000100100101000000100",
			5318 => "0000000101001101101001",
			5319 => "0000000101001101101001",
			5320 => "1111111101001101101001",
			5321 => "0011011110011000001100",
			5322 => "0001000110011100000100",
			5323 => "1111111101001101101001",
			5324 => "0000000010010000000100",
			5325 => "0000000101001101101001",
			5326 => "0000000101001101101001",
			5327 => "0010000101101100001000",
			5328 => "0001101010011000000100",
			5329 => "0000000101001101101001",
			5330 => "0000000101001101101001",
			5331 => "0000001000001000000100",
			5332 => "0000001101001101101001",
			5333 => "0000000101001101101001",
			5334 => "0000110010111000000100",
			5335 => "0000000101001101101001",
			5336 => "0000000101001101101001",
			5337 => "0000000101001101101001",
			5338 => "0001110001010001001100",
			5339 => "0001000010111001001000",
			5340 => "0000001100000100100000",
			5341 => "0010001111111100001100",
			5342 => "0011000110110100000100",
			5343 => "0000000101010000000101",
			5344 => "0001011001010100000100",
			5345 => "1111111101010000000101",
			5346 => "0000000101010000000101",
			5347 => "0001100100000000010000",
			5348 => "0010111010100100001000",
			5349 => "0001010101010100000100",
			5350 => "0000000101010000000101",
			5351 => "0000001101010000000101",
			5352 => "0010001111001000000100",
			5353 => "1111111101010000000101",
			5354 => "0000000101010000000101",
			5355 => "0000001101010000000101",
			5356 => "0011101111100100010100",
			5357 => "0000000100100000010000",
			5358 => "0011101101111100001000",
			5359 => "0011010111011100000100",
			5360 => "1111111101010000000101",
			5361 => "0000000101010000000101",
			5362 => "0001001100101100000100",
			5363 => "0000000101010000000101",
			5364 => "0000000101010000000101",
			5365 => "1111111101010000000101",
			5366 => "0000100001111000000100",
			5367 => "0000001101010000000101",
			5368 => "0001011000111000001000",
			5369 => "0001111001010000000100",
			5370 => "1111111101010000000101",
			5371 => "0000000101010000000101",
			5372 => "0001111100010000000100",
			5373 => "0000000101010000000101",
			5374 => "0000000101010000000101",
			5375 => "0000000101010000000101",
			5376 => "1111111101010000000101",
			5377 => "0010001001001100001000",
			5378 => "0000110110001100000100",
			5379 => "0000000101010011000001",
			5380 => "0000000101010011000001",
			5381 => "0001110001010001010100",
			5382 => "0000011000011000110000",
			5383 => "0001001100101100011100",
			5384 => "0011010110001100001100",
			5385 => "0001000011110000000100",
			5386 => "0000000101010011000001",
			5387 => "0001111100010000000100",
			5388 => "0000000101010011000001",
			5389 => "0000000101010011000001",
			5390 => "0001111010000100001000",
			5391 => "0011000111011100000100",
			5392 => "0000000101010011000001",
			5393 => "0000000101010011000001",
			5394 => "0011101111000100000100",
			5395 => "0000000101010011000001",
			5396 => "0000000101010011000001",
			5397 => "0011000101010100000100",
			5398 => "0000000101010011000001",
			5399 => "0011001100101000001000",
			5400 => "0010101100001100000100",
			5401 => "0000000101010011000001",
			5402 => "0000000101010011000001",
			5403 => "0010101010011100000100",
			5404 => "0000000101010011000001",
			5405 => "0000000101010011000001",
			5406 => "0011010101011100011000",
			5407 => "0001011000111000001100",
			5408 => "0011001110011000000100",
			5409 => "0000000101010011000001",
			5410 => "0000101000110100000100",
			5411 => "0000000101010011000001",
			5412 => "0000000101010011000001",
			5413 => "0010101000101000000100",
			5414 => "0000000101010011000001",
			5415 => "0001011001011000000100",
			5416 => "0000000101010011000001",
			5417 => "0000000101010011000001",
			5418 => "0001111100010000001000",
			5419 => "0001101100011100000100",
			5420 => "0000000101010011000001",
			5421 => "0000000101010011000001",
			5422 => "0000000101010011000001",
			5423 => "0000000101010011000001",
			5424 => "0001100100010001101000",
			5425 => "0011001100101000111100",
			5426 => "0010101100001100111000",
			5427 => "0000000011101100011100",
			5428 => "0000010001110000001100",
			5429 => "0010001001001100000100",
			5430 => "1111111101010110010111",
			5431 => "0010110011010000000100",
			5432 => "0000000101010110010111",
			5433 => "1111111101010110010111",
			5434 => "0011101000100000001000",
			5435 => "0010111010100100000100",
			5436 => "0000001101010110010111",
			5437 => "1111111101010110010111",
			5438 => "0001010110101100000100",
			5439 => "0000001101010110010111",
			5440 => "0000001101010110010111",
			5441 => "0011101001101100001100",
			5442 => "0000011000011000001000",
			5443 => "0000010000011000000100",
			5444 => "0000000101010110010111",
			5445 => "1111111101010110010111",
			5446 => "0000001101010110010111",
			5447 => "0001001000000100001000",
			5448 => "0001011101001000000100",
			5449 => "0000000101010110010111",
			5450 => "1111111101010110010111",
			5451 => "0000111000100000000100",
			5452 => "0000001101010110010111",
			5453 => "0000000101010110010111",
			5454 => "1111111101010110010111",
			5455 => "0000110001001000011000",
			5456 => "0011100101110000010000",
			5457 => "0000000111101000001000",
			5458 => "0000000110000100000100",
			5459 => "1111111101010110010111",
			5460 => "0000000101010110010111",
			5461 => "0000000000010000000100",
			5462 => "1111111101010110010111",
			5463 => "1111111101010110010111",
			5464 => "0001101111111000000100",
			5465 => "0000000101010110010111",
			5466 => "1111111101010110010111",
			5467 => "0000000100111100010000",
			5468 => "0011101111111000001100",
			5469 => "0000000010111100001000",
			5470 => "0010101100110100000100",
			5471 => "0000001101010110010111",
			5472 => "0000000101010110010111",
			5473 => "1111111101010110010111",
			5474 => "0000001101010110010111",
			5475 => "1111111101010110010111",
			5476 => "1111111101010110010111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1757, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3651, initial_addr_3'length));
	end generate gen_rom_7;

	gen_rom_8: if SELECT_ROM = 8 generate
		bank <= (
			0 => "0001001011111000011100",
			1 => "0001001001010000010000",
			2 => "0001011010011100001100",
			3 => "0001000110101100000100",
			4 => "1101101000000010010101",
			5 => "0000010111100100000100",
			6 => "1101110000000010010101",
			7 => "1101101000000010010101",
			8 => "1101110000000010010101",
			9 => "0010000101101100000100",
			10 => "1110010000000010010101",
			11 => "0000000111110100000100",
			12 => "1101101000000010010101",
			13 => "1101101000000010010101",
			14 => "0010110110000000100100",
			15 => "0000001011011100010100",
			16 => "0011011110011000001100",
			17 => "0001111000000100000100",
			18 => "1110101000000010010101",
			19 => "0000001010111100000100",
			20 => "1110000000000010010101",
			21 => "1110010000000010010101",
			22 => "0001111100010000000100",
			23 => "1101111000000010010101",
			24 => "1101101000000010010101",
			25 => "0000010001100100001100",
			26 => "0010101100110100001000",
			27 => "0011011110011000000100",
			28 => "1110101000000010010101",
			29 => "1110001000000010010101",
			30 => "1110101000000010010101",
			31 => "1101111000000010010101",
			32 => "0010111101101000000100",
			33 => "1101111000000010010101",
			34 => "0010111010000100000100",
			35 => "1101101000000010010101",
			36 => "1101101000000010010101",
			37 => "0011101101000100110100",
			38 => "0011000101010100010000",
			39 => "0011010110110100001000",
			40 => "0000010001110000000100",
			41 => "0000000000000100101001",
			42 => "0000000000000100101001",
			43 => "0001010001011000000100",
			44 => "0000000000000100101001",
			45 => "0000001000000100101001",
			46 => "0000001100000100001000",
			47 => "0010000101011100000100",
			48 => "0000000000000100101001",
			49 => "1111111000000100101001",
			50 => "0011011011101100001000",
			51 => "0010011010000100000100",
			52 => "1111111000000100101001",
			53 => "0000001000000100101001",
			54 => "0011100101110000001000",
			55 => "0010101001011000000100",
			56 => "0000000000000100101001",
			57 => "0000001000000100101001",
			58 => "0000000000001100000100",
			59 => "1111111000000100101001",
			60 => "0000001101001100000100",
			61 => "0000000000000100101001",
			62 => "0000001000000100101001",
			63 => "0011001001001000001100",
			64 => "0010000101011100001000",
			65 => "0010001001001100000100",
			66 => "0000000000000100101001",
			67 => "0000000000000100101001",
			68 => "1111111000000100101001",
			69 => "0000011101000000001000",
			70 => "0000110010010100000100",
			71 => "0000001000000100101001",
			72 => "0000000000000100101001",
			73 => "0000000000000100101001",
			74 => "0000001011100000110100",
			75 => "0010110111011100010100",
			76 => "0001000110101100000100",
			77 => "0000000000000110101101",
			78 => "0001001110111000001100",
			79 => "0001011110010100001000",
			80 => "0001011110001100000100",
			81 => "0000000000000110101101",
			82 => "0000000000000110101101",
			83 => "0000000000000110101101",
			84 => "0000000000000110101101",
			85 => "0000100100011100000100",
			86 => "0000000000000110101101",
			87 => "0000001010111100001000",
			88 => "0010001001000100000100",
			89 => "0000000000000110101101",
			90 => "0000000000000110101101",
			91 => "0011000101011100001000",
			92 => "0001110110101100000100",
			93 => "0000000000000110101101",
			94 => "0000000000000110101101",
			95 => "0000000100100000000100",
			96 => "0000000000000110101101",
			97 => "0011100101001000000100",
			98 => "0000000000000110101101",
			99 => "0000000000000110101101",
			100 => "0001011111100000001000",
			101 => "0000111001000000000100",
			102 => "0000000000000110101101",
			103 => "0000000000000110101101",
			104 => "0010100111010100000100",
			105 => "0000000000000110101101",
			106 => "0000000000000110101101",
			107 => "0001000110101100000100",
			108 => "1111111000000111111001",
			109 => "0000101010000000100000",
			110 => "0010101001111100011100",
			111 => "0010100000111000010000",
			112 => "0001111000000100000100",
			113 => "0000001000000111111001",
			114 => "0000100100011100000100",
			115 => "1111111000000111111001",
			116 => "0000010110010000000100",
			117 => "0000000000000111111001",
			118 => "0000000000000111111001",
			119 => "0010001001000100000100",
			120 => "0000001000000111111001",
			121 => "0001100010000000000100",
			122 => "0000000000000111111001",
			123 => "0000001000000111111001",
			124 => "1111111000000111111001",
			125 => "1111111000000111111001",
			126 => "0011010011010000111000",
			127 => "0001101001111100001100",
			128 => "0001111000000100001000",
			129 => "0001010001011000000100",
			130 => "0000000000001010000101",
			131 => "0000000000001010000101",
			132 => "0000000000001010000101",
			133 => "0011101001111100010000",
			134 => "0000000111101000000100",
			135 => "0000000000001010000101",
			136 => "0010101000100000000100",
			137 => "0000000000001010000101",
			138 => "0010101010011100000100",
			139 => "0000000000001010000101",
			140 => "0000000000001010000101",
			141 => "0000100111010000001000",
			142 => "0001010001101000000100",
			143 => "0000000000001010000101",
			144 => "0000000000001010000101",
			145 => "0010011010000100001100",
			146 => "0011101010011000000100",
			147 => "0000000000001010000101",
			148 => "0010110111011100000100",
			149 => "0000000000001010000101",
			150 => "0000000000001010000101",
			151 => "0010001001000100000100",
			152 => "0000000000001010000101",
			153 => "0000000000001010000101",
			154 => "0000010001110000000100",
			155 => "0000000000001010000101",
			156 => "0011110011101100000100",
			157 => "0000000000001010000101",
			158 => "0000101110110100000100",
			159 => "0000000000001010000101",
			160 => "0000000000001010000101",
			161 => "0001010001011000000100",
			162 => "1111111000001011111001",
			163 => "0011011010100100011100",
			164 => "0000111011000000001000",
			165 => "0000110100101100000100",
			166 => "0000000000001011111001",
			167 => "1111111000001011111001",
			168 => "0000010110010000001100",
			169 => "0011111010011000000100",
			170 => "0000000000001011111001",
			171 => "0011000101010100000100",
			172 => "0000000000001011111001",
			173 => "0000001000001011111001",
			174 => "0000000010111100000100",
			175 => "0000000000001011111001",
			176 => "0000001000001011111001",
			177 => "0010110101011100001000",
			178 => "0010001111111100000100",
			179 => "0000000000001011111001",
			180 => "1111111000001011111001",
			181 => "0001000110011100000100",
			182 => "1111111000001011111001",
			183 => "0000111001000000000100",
			184 => "0000001000001011111001",
			185 => "0000100010111100000100",
			186 => "1111111000001011111001",
			187 => "0000011000011000000100",
			188 => "0000001000001011111001",
			189 => "0000000000001011111001",
			190 => "0011101010011000111100",
			191 => "0000000111101000011000",
			192 => "0010011001000100001000",
			193 => "0001010001011000000100",
			194 => "0000000000001110111101",
			195 => "0000000000001110111101",
			196 => "0011000101010100001000",
			197 => "0011101110010100000100",
			198 => "0000000000001110111101",
			199 => "0000000000001110111101",
			200 => "0010000101011100000100",
			201 => "0000000000001110111101",
			202 => "0000000000001110111101",
			203 => "0001011100110100001100",
			204 => "0001101110000000001000",
			205 => "0000111111101000000100",
			206 => "0000000000001110111101",
			207 => "0000000000001110111101",
			208 => "0000000000001110111101",
			209 => "0011010111011100001100",
			210 => "0001111101001000001000",
			211 => "0001001001011000000100",
			212 => "0000000000001110111101",
			213 => "0000000000001110111101",
			214 => "0000000000001110111101",
			215 => "0000100010111100000100",
			216 => "0000000000001110111101",
			217 => "0001000100100100000100",
			218 => "0000000000001110111101",
			219 => "0000000000001110111101",
			220 => "0000001011011000001000",
			221 => "0001110001010000000100",
			222 => "0000000000001110111101",
			223 => "0000000000001110111101",
			224 => "0000000111110100010000",
			225 => "0000111011000000001000",
			226 => "0000101000100100000100",
			227 => "0000000000001110111101",
			228 => "0000000000001110111101",
			229 => "0000111001111100000100",
			230 => "0000000000001110111101",
			231 => "0000000000001110111101",
			232 => "0001011111100000001000",
			233 => "0000111001000000000100",
			234 => "0000000000001110111101",
			235 => "0000000000001110111101",
			236 => "0000111010100000000100",
			237 => "0000000000001110111101",
			238 => "0000000000001110111101",
			239 => "0001010001011000000100",
			240 => "1111111000010000011001",
			241 => "0000011101000000100100",
			242 => "0000111001111100100000",
			243 => "0010101100110100010100",
			244 => "0001111000000100001000",
			245 => "0000111011111000000100",
			246 => "0000001000010000011001",
			247 => "0000001000010000011001",
			248 => "0000100100011100000100",
			249 => "1111111000010000011001",
			250 => "0011010111011100000100",
			251 => "0000001000010000011001",
			252 => "0000000000010000011001",
			253 => "0001011010011000001000",
			254 => "0010001001000100000100",
			255 => "0000001000010000011001",
			256 => "0000000000010000011001",
			257 => "0000001000010000011001",
			258 => "1111111000010000011001",
			259 => "0010000000110000000100",
			260 => "0000000000010000011001",
			261 => "1111111000010000011001",
			262 => "0010001001000100111100",
			263 => "0010101100110100110100",
			264 => "0001101010011000011100",
			265 => "0001011100110100010000",
			266 => "0010110011010000001000",
			267 => "0001010001011000000100",
			268 => "0000000000010010111101",
			269 => "0000000000010010111101",
			270 => "0010010101101100000100",
			271 => "0000000000010010111101",
			272 => "0000000000010010111101",
			273 => "0001101101101100000100",
			274 => "0000000000010010111101",
			275 => "0011011110011000000100",
			276 => "0000000000010010111101",
			277 => "0000000000010010111101",
			278 => "0000100111010000001000",
			279 => "0011011011101100000100",
			280 => "0000000000010010111101",
			281 => "0000000000010010111101",
			282 => "0010011010000100001100",
			283 => "0001100010000000000100",
			284 => "0000000000010010111101",
			285 => "0000011001100100000100",
			286 => "0000000000010010111101",
			287 => "0000000000010010111101",
			288 => "0000000000010010111101",
			289 => "0010011000000100000100",
			290 => "0000000000010010111101",
			291 => "0000000000010010111101",
			292 => "0010011101101000001000",
			293 => "0010101011000000000100",
			294 => "0000000000010010111101",
			295 => "0000000000010010111101",
			296 => "0001011010001100001000",
			297 => "0000110000111000000100",
			298 => "0000000000010010111101",
			299 => "0000000000010010111101",
			300 => "0010101101101100000100",
			301 => "0000000000010010111101",
			302 => "0000000000010010111101",
			303 => "0001000110101100000100",
			304 => "1111111000010100011001",
			305 => "0000100111000100100100",
			306 => "0010101001111100100000",
			307 => "0001111000101000011000",
			308 => "0011010111011100010000",
			309 => "0011101010011000001000",
			310 => "0000001110101100000100",
			311 => "0000000000010100011001",
			312 => "0000001000010100011001",
			313 => "0001000001011000000100",
			314 => "0000000000010100011001",
			315 => "0000000000010100011001",
			316 => "0000100010111100000100",
			317 => "1111111000010100011001",
			318 => "0000000000010100011001",
			319 => "0001101111110000000100",
			320 => "0000001000010100011001",
			321 => "0000001000010100011001",
			322 => "1111111000010100011001",
			323 => "0001011010100000000100",
			324 => "1111111000010100011001",
			325 => "0000000000010100011001",
			326 => "0010001111001001000000",
			327 => "0010101011000000010100",
			328 => "0001111000000100001000",
			329 => "0001010000111100000100",
			330 => "0000000000010110101101",
			331 => "0000000000010110101101",
			332 => "0010011010000100000100",
			333 => "0000000000010110101101",
			334 => "0010010011000000000100",
			335 => "0000000000010110101101",
			336 => "0000000000010110101101",
			337 => "0010101010011100011000",
			338 => "0011010111011100010100",
			339 => "0011111111111000001000",
			340 => "0000010111110000000100",
			341 => "0000000000010110101101",
			342 => "0000000000010110101101",
			343 => "0010001001001100000100",
			344 => "0000000000010110101101",
			345 => "0010100000111100000100",
			346 => "0000000000010110101101",
			347 => "0000000000010110101101",
			348 => "0000000000010110101101",
			349 => "0010101100001100000100",
			350 => "0000000000010110101101",
			351 => "0000011000111100000100",
			352 => "0000000000010110101101",
			353 => "0000000100011000000100",
			354 => "0000000000010110101101",
			355 => "0000110100000000000100",
			356 => "0000000000010110101101",
			357 => "0000000000010110101101",
			358 => "0001001110010100000100",
			359 => "0000000000010110101101",
			360 => "0001010011101100000100",
			361 => "0000000000010110101101",
			362 => "0000000000010110101101",
			363 => "0000010110010000111000",
			364 => "0010001111111100011100",
			365 => "0001011110010100011000",
			366 => "0001111100010000010000",
			367 => "0001111111011000001000",
			368 => "0010011100101000000100",
			369 => "0000000000011001100001",
			370 => "0000000000011001100001",
			371 => "0001101011110000000100",
			372 => "0000000000011001100001",
			373 => "0000000000011001100001",
			374 => "0000001011001000000100",
			375 => "0000000000011001100001",
			376 => "0000000000011001100001",
			377 => "0000000000011001100001",
			378 => "0001010010001100010100",
			379 => "0011111010011000001100",
			380 => "0000010111110000001000",
			381 => "0010000101101100000100",
			382 => "0000000000011001100001",
			383 => "0000000000011001100001",
			384 => "0000000000011001100001",
			385 => "0001011010011100000100",
			386 => "0000000000011001100001",
			387 => "0000000000011001100001",
			388 => "0011001001001000000100",
			389 => "0000000000011001100001",
			390 => "0000000000011001100001",
			391 => "0010010110000000001000",
			392 => "0001011100011100000100",
			393 => "0000000000011001100001",
			394 => "0000000000011001100001",
			395 => "0001001100001100010100",
			396 => "0000001101001100000100",
			397 => "0000000000011001100001",
			398 => "0000101110110100001100",
			399 => "0000110001001000001000",
			400 => "0000000000011100000100",
			401 => "0000000000011001100001",
			402 => "0000000000011001100001",
			403 => "0000000000011001100001",
			404 => "0000000000011001100001",
			405 => "0010101101101100000100",
			406 => "0000000000011001100001",
			407 => "0000000000011001100001",
			408 => "0011011010100100111000",
			409 => "0001011110010100100100",
			410 => "0011011011101100010000",
			411 => "0001111111011000001000",
			412 => "0001010001011000000100",
			413 => "0000000000011100101101",
			414 => "0000000000011100101101",
			415 => "0001111101001000000100",
			416 => "0000000000011100101101",
			417 => "0000000000011100101101",
			418 => "0000001100000100001100",
			419 => "0011100001010100001000",
			420 => "0001110101111000000100",
			421 => "0000000000011100101101",
			422 => "0000000000011100101101",
			423 => "0000000000011100101101",
			424 => "0001001001010100000100",
			425 => "0000000000011100101101",
			426 => "0000000000011100101101",
			427 => "0011011110011000001100",
			428 => "0001001110111000000100",
			429 => "0000000000011100101101",
			430 => "0000010001110000000100",
			431 => "0000000000011100101101",
			432 => "0000000000011100101101",
			433 => "0010001111111100000100",
			434 => "0000000000011100101101",
			435 => "0000000000011100101101",
			436 => "0001101111111000001000",
			437 => "0011000011010000000100",
			438 => "0000000000011100101101",
			439 => "0000000000011100101101",
			440 => "0010110101011100001100",
			441 => "0010110111011100001000",
			442 => "0001101111010100000100",
			443 => "0000000000011100101101",
			444 => "0000000000011100101101",
			445 => "0000000000011100101101",
			446 => "0001000001010100001100",
			447 => "0010000000110000001000",
			448 => "0010100000111100000100",
			449 => "0000000000011100101101",
			450 => "0000000000011100101101",
			451 => "0000000000011100101101",
			452 => "0011101100100000001000",
			453 => "0000010111100100000100",
			454 => "0000000000011100101101",
			455 => "0000000000011100101101",
			456 => "0001110001011000000100",
			457 => "0000000000011100101101",
			458 => "0000000000011100101101",
			459 => "0010001001000100111100",
			460 => "0010101011000000010100",
			461 => "0001110011001000001100",
			462 => "0001111010000100000100",
			463 => "0000000000011111010001",
			464 => "0010011100101000000100",
			465 => "0000000000011111010001",
			466 => "0000000000011111010001",
			467 => "0010011010000100000100",
			468 => "0000000000011111010001",
			469 => "0000000000011111010001",
			470 => "0011010111011100100000",
			471 => "0010010011000000011000",
			472 => "0000010111110000010000",
			473 => "0000110000111100001000",
			474 => "0010100000111100000100",
			475 => "0000000000011111010001",
			476 => "0000000000011111010001",
			477 => "0001001110111000000100",
			478 => "0000000000011111010001",
			479 => "0000000000011111010001",
			480 => "0001101010011000000100",
			481 => "0000000000011111010001",
			482 => "0000000000011111010001",
			483 => "0000100101111100000100",
			484 => "0000000000011111010001",
			485 => "0000000000011111010001",
			486 => "0000111010011100000100",
			487 => "0000000000011111010001",
			488 => "0000000000011111010001",
			489 => "0011011011101100000100",
			490 => "0000000000011111010001",
			491 => "0011111110111100000100",
			492 => "0000000000011111010001",
			493 => "0011101010011000000100",
			494 => "0000000000011111010001",
			495 => "0001011010001100000100",
			496 => "0000000000011111010001",
			497 => "0001010011101100000100",
			498 => "0000000000011111010001",
			499 => "0000000000011111010001",
			500 => "0001000110101100000100",
			501 => "1111111000100000110101",
			502 => "0000011101000000101000",
			503 => "0001000100100100100100",
			504 => "0010101100110100010100",
			505 => "0001111000000100001000",
			506 => "0010101011000000000100",
			507 => "0000001000100000110101",
			508 => "0000001000100000110101",
			509 => "0000100100011100000100",
			510 => "1111111000100000110101",
			511 => "0000001011100000000100",
			512 => "0000001000100000110101",
			513 => "0000000000100000110101",
			514 => "0000100101000100001000",
			515 => "0010000101101100000100",
			516 => "0000001000100000110101",
			517 => "0000000000100000110101",
			518 => "0001110110011100000100",
			519 => "0000001000100000110101",
			520 => "0000001000100000110101",
			521 => "1111111000100000110101",
			522 => "0010000000110000000100",
			523 => "0000000000100000110101",
			524 => "1111111000100000110101",
			525 => "0001010001011000000100",
			526 => "1111111000100010001001",
			527 => "0000101010000000100100",
			528 => "0010111010000100100000",
			529 => "0010100001101000011000",
			530 => "0010011001000100001000",
			531 => "0001011110001100000100",
			532 => "0000001000100010001001",
			533 => "0000001000100010001001",
			534 => "0000001110101100001000",
			535 => "0001000011000100000100",
			536 => "1111111000100010001001",
			537 => "0000000000100010001001",
			538 => "0011101111111000000100",
			539 => "0000001000100010001001",
			540 => "0000000000100010001001",
			541 => "0011111110111100000100",
			542 => "0000000000100010001001",
			543 => "0000001000100010001001",
			544 => "1111111000100010001001",
			545 => "1111111000100010001001",
			546 => "0001011110111000000100",
			547 => "1111111000100100011101",
			548 => "0010001001000100100100",
			549 => "0011101111100100010000",
			550 => "0001011110010100001000",
			551 => "0010011001000100000100",
			552 => "0000001000100100011101",
			553 => "0000000000100100011101",
			554 => "0011100101110000000100",
			555 => "0000001000100100011101",
			556 => "0000001000100100011101",
			557 => "0000000100011000000100",
			558 => "1111111000100100011101",
			559 => "0011101111111000000100",
			560 => "0000001000100100011101",
			561 => "0001111101001000000100",
			562 => "1111111000100100011101",
			563 => "0000101011010100000100",
			564 => "0000000000100100011101",
			565 => "0000001000100100011101",
			566 => "0001010001011100010000",
			567 => "0010100000111100001000",
			568 => "0010101000100000000100",
			569 => "1111111000100100011101",
			570 => "0000000000100100011101",
			571 => "0000110011110100000100",
			572 => "1111111000100100011101",
			573 => "0000000000100100011101",
			574 => "0011110010001000001000",
			575 => "0001001110010100000100",
			576 => "0000000000100100011101",
			577 => "1111111000100100011101",
			578 => "0010101101101100001000",
			579 => "0011100001101100000100",
			580 => "0000001000100100011101",
			581 => "0000000000100100011101",
			582 => "1111111000100100011101",
			583 => "0001000110101100000100",
			584 => "1111111000100110011001",
			585 => "0010010110000000001100",
			586 => "0001010010111000001000",
			587 => "0001111000000100000100",
			588 => "0000000000100110011001",
			589 => "0000000000100110011001",
			590 => "0000001000100110011001",
			591 => "0010001111111100010000",
			592 => "0001010001111100001000",
			593 => "0000000100011000000100",
			594 => "1111111000100110011001",
			595 => "0000000000100110011001",
			596 => "0011001001001000000100",
			597 => "0000001000100110011001",
			598 => "0000000000100110011001",
			599 => "0000010111110000001000",
			600 => "0001000001011000000100",
			601 => "0000000000100110011001",
			602 => "1111111000100110011001",
			603 => "0001000000111100001100",
			604 => "0000001011011100000100",
			605 => "1111111000100110011001",
			606 => "0001001100101100000100",
			607 => "0000000000100110011001",
			608 => "0000000000100110011001",
			609 => "0000010110010000000100",
			610 => "0000001000100110011001",
			611 => "0001001100001100000100",
			612 => "0000000000100110011001",
			613 => "0000000000100110011001",
			614 => "0000001011100001000100",
			615 => "0010010110000000001100",
			616 => "0001010001011000000100",
			617 => "0000000000101000111101",
			618 => "0011010110001100000100",
			619 => "0000000000101000111101",
			620 => "0000001000101000111101",
			621 => "0000001110101100011100",
			622 => "0011100100000000010100",
			623 => "0001010001010100010000",
			624 => "0001110110101100001000",
			625 => "0000011001100100000100",
			626 => "0000000000101000111101",
			627 => "1111111000101000111101",
			628 => "0000011001100000000100",
			629 => "0000000000101000111101",
			630 => "0000000000101000111101",
			631 => "0000000000101000111101",
			632 => "0001010010111000000100",
			633 => "0000000000101000111101",
			634 => "1111111000101000111101",
			635 => "0011101011110000001100",
			636 => "0011010111011100000100",
			637 => "0000001000101000111101",
			638 => "0001111101001000000100",
			639 => "0000000000101000111101",
			640 => "0000000000101000111101",
			641 => "0000001101001100000100",
			642 => "0000000000101000111101",
			643 => "0001110110101100000100",
			644 => "0000000000101000111101",
			645 => "0011010101010100000100",
			646 => "0000001000101000111101",
			647 => "0000000000101000111101",
			648 => "0001011111100000001000",
			649 => "0000111001000000000100",
			650 => "0000000000101000111101",
			651 => "0000000000101000111101",
			652 => "0000111010100000000100",
			653 => "0000000000101000111101",
			654 => "0000000000101000111101",
			655 => "0001000110101100000100",
			656 => "1111111000101010100001",
			657 => "0010001111011000101100",
			658 => "0001011110010100010100",
			659 => "0001111000000100001000",
			660 => "0010000101011100000100",
			661 => "0000001000101010100001",
			662 => "0000001000101010100001",
			663 => "0011011011101100000100",
			664 => "1111111000101010100001",
			665 => "0000000000001100000100",
			666 => "0000000000101010100001",
			667 => "0000000000101010100001",
			668 => "0011100101110000000100",
			669 => "0000001000101010100001",
			670 => "0000000010010000000100",
			671 => "1111111000101010100001",
			672 => "0011101011110000001000",
			673 => "0001010111010100000100",
			674 => "0000001000101010100001",
			675 => "0000001000101010100001",
			676 => "0000001101001100000100",
			677 => "1111111000101010100001",
			678 => "0000001000101010100001",
			679 => "1111111000101010100001",
			680 => "0000101011100001001100",
			681 => "0000001101001100100100",
			682 => "0001100010010100011100",
			683 => "0010011001000100001000",
			684 => "0001010001011000000100",
			685 => "0000000000101101001101",
			686 => "0000001000101101001101",
			687 => "0000001011011100001100",
			688 => "0011101111100100001000",
			689 => "0000101000101100000100",
			690 => "0000000000101101001101",
			691 => "0000000000101101001101",
			692 => "1111111000101101001101",
			693 => "0001101011110000000100",
			694 => "0000000000101101001101",
			695 => "0000001000101101001101",
			696 => "0011011011101100000100",
			697 => "0000000000101101001101",
			698 => "1111111000101101001101",
			699 => "0000000000011100010100",
			700 => "0011010101010100001000",
			701 => "0001001001010100000100",
			702 => "0000000000101101001101",
			703 => "0000001000101101001101",
			704 => "0000011000011000000100",
			705 => "0000000000101101001101",
			706 => "0001110100101100000100",
			707 => "0000000000101101001101",
			708 => "0000000000101101001101",
			709 => "0001110110101100000100",
			710 => "1111111000101101001101",
			711 => "0000111101101100001100",
			712 => "0000011101000000001000",
			713 => "0001001111101000000100",
			714 => "0000000000101101001101",
			715 => "0000001000101101001101",
			716 => "0000000000101101001101",
			717 => "0000000000101101001101",
			718 => "0000111001000000000100",
			719 => "1111111000101101001101",
			720 => "0000011101000000000100",
			721 => "0000000000101101001101",
			722 => "0000000000101101001101",
			723 => "0001001111101000001100",
			724 => "0001000110101100000100",
			725 => "1111111000101111000001",
			726 => "0000001000011100000100",
			727 => "0000001000101111000001",
			728 => "1111111000101111000001",
			729 => "0011011001001000101100",
			730 => "0001000000100000101000",
			731 => "0001011110010100001100",
			732 => "0001111000000100000100",
			733 => "0000010000101111000001",
			734 => "0011110101001000000100",
			735 => "1111111000101111000001",
			736 => "0000001000101111000001",
			737 => "0000000010111100001100",
			738 => "0000010110010000001000",
			739 => "0010001111111100000100",
			740 => "0000010000101111000001",
			741 => "0000001000101111000001",
			742 => "0000000000101111000001",
			743 => "0010011111011000001000",
			744 => "0011101111111000000100",
			745 => "0000010000101111000001",
			746 => "0000001000101111000001",
			747 => "0000011001100000000100",
			748 => "0000010000101111000001",
			749 => "0000010000101111000001",
			750 => "1111111000101111000001",
			751 => "1111111000101111000001",
			752 => "0001011010011100001100",
			753 => "0001010001011000000100",
			754 => "1111111000110001001101",
			755 => "0000000111001100000100",
			756 => "0000010000110001001101",
			757 => "1111111000110001001101",
			758 => "0011011001001000110000",
			759 => "0000111001111100101100",
			760 => "0000001110101100010100",
			761 => "0011000101010100001000",
			762 => "0010111010100100000100",
			763 => "0000100000110001001101",
			764 => "0000011000110001001101",
			765 => "0011011110011000000100",
			766 => "0000010000110001001101",
			767 => "0001111100010000000100",
			768 => "0000000000110001001101",
			769 => "1111111000110001001101",
			770 => "0000011001100000010000",
			771 => "0000100010111100001000",
			772 => "0011100010011100000100",
			773 => "0000100000110001001101",
			774 => "0000001000110001001101",
			775 => "0010011010000100000100",
			776 => "0000011000110001001101",
			777 => "0000011000110001001101",
			778 => "0001011010100000000100",
			779 => "0000001000110001001101",
			780 => "0000011000110001001101",
			781 => "1111111000110001001101",
			782 => "0010111101101000001000",
			783 => "0001101000010100000100",
			784 => "0000000000110001001101",
			785 => "1111111000110001001101",
			786 => "1111111000110001001101",
			787 => "0001000110101100000100",
			788 => "1111111000110011011001",
			789 => "0010110111011100010100",
			790 => "0001011110010100001100",
			791 => "0000111011111000000100",
			792 => "0000001000110011011001",
			793 => "0010100000111100000100",
			794 => "0000000000110011011001",
			795 => "0000000000110011011001",
			796 => "0001111100010000000100",
			797 => "0000001000110011011001",
			798 => "0000000000110011011001",
			799 => "0001010001011100010100",
			800 => "0000000000001100000100",
			801 => "1111111000110011011001",
			802 => "0011100010011100000100",
			803 => "0000001000110011011001",
			804 => "0001111101001000000100",
			805 => "1111111000110011011001",
			806 => "0010101010011100000100",
			807 => "0000000000110011011001",
			808 => "1111111000110011011001",
			809 => "0010010011000000001000",
			810 => "0011111001011100000100",
			811 => "0000001000110011011001",
			812 => "0000000000110011011001",
			813 => "0011110011101100001100",
			814 => "0011100000010100001000",
			815 => "0000100010111100000100",
			816 => "0000000000110011011001",
			817 => "0000000000110011011001",
			818 => "1111111000110011011001",
			819 => "0000011101000000000100",
			820 => "0000001000110011011001",
			821 => "1111111000110011011001",
			822 => "0011011010100100110100",
			823 => "0000111000100000100000",
			824 => "0001111000000100001000",
			825 => "0001010001011000000100",
			826 => "0000000000110110101101",
			827 => "0000000000110110101101",
			828 => "0000001011011100001100",
			829 => "0010011001000100000100",
			830 => "0000000000110110101101",
			831 => "0011001001001000000100",
			832 => "0000000000110110101101",
			833 => "0000000000110110101101",
			834 => "0000000111001100001000",
			835 => "0001001001010100000100",
			836 => "0000000000110110101101",
			837 => "0000000000110110101101",
			838 => "0000000000110110101101",
			839 => "0010010011000000001100",
			840 => "0011101010110100000100",
			841 => "0000000000110110101101",
			842 => "0001100110100000000100",
			843 => "0000000000110110101101",
			844 => "0000000000110110101101",
			845 => "0010001111111100000100",
			846 => "0000000000110110101101",
			847 => "0000000000110110101101",
			848 => "0000010001110000001000",
			849 => "0010001001000100000100",
			850 => "0000000000110110101101",
			851 => "0000000000110110101101",
			852 => "0010100000111000100100",
			853 => "0000100001100000010000",
			854 => "0001111100010000001100",
			855 => "0001111000111000001000",
			856 => "0010011001000100000100",
			857 => "0000000000110110101101",
			858 => "0000000000110110101101",
			859 => "0000000000110110101101",
			860 => "0000000000110110101101",
			861 => "0010110011010000001000",
			862 => "0010010110000000000100",
			863 => "0000000000110110101101",
			864 => "0000000000110110101101",
			865 => "0001100010011000000100",
			866 => "0000000000110110101101",
			867 => "0010010011000000000100",
			868 => "0000000000110110101101",
			869 => "0000000000110110101101",
			870 => "0010101101101100001000",
			871 => "0011110111101000000100",
			872 => "0000000000110110101101",
			873 => "0000000000110110101101",
			874 => "0000000000110110101101",
			875 => "0010110111011100100000",
			876 => "0001011110010100011000",
			877 => "0001111000000100001000",
			878 => "0001010001011000000100",
			879 => "0000000000111001111001",
			880 => "0000000000111001111001",
			881 => "0000100100100000000100",
			882 => "0000000000111001111001",
			883 => "0000100011100000001000",
			884 => "0000111100010000000100",
			885 => "0000000000111001111001",
			886 => "0000000000111001111001",
			887 => "0000000000111001111001",
			888 => "0001010001011100000100",
			889 => "0000000000111001111001",
			890 => "0000000000111001111001",
			891 => "0001011101111100100100",
			892 => "0000000000001100001100",
			893 => "0010011001000100000100",
			894 => "0000000000111001111001",
			895 => "0000111001000000000100",
			896 => "1111111000111001111001",
			897 => "0000000000111001111001",
			898 => "0011100010011100001000",
			899 => "0000100111000000000100",
			900 => "0000000000111001111001",
			901 => "0000000000111001111001",
			902 => "0011110001101100000100",
			903 => "0000000000111001111001",
			904 => "0000110001001000000100",
			905 => "0000000000111001111001",
			906 => "0010101010011100000100",
			907 => "0000000000111001111001",
			908 => "0000000000111001111001",
			909 => "0010010011000000001000",
			910 => "0011101010110100000100",
			911 => "0000000000111001111001",
			912 => "0000000000111001111001",
			913 => "0000100010111100000100",
			914 => "0000000000111001111001",
			915 => "0011101110000000001100",
			916 => "0010001111001000000100",
			917 => "0000000000111001111001",
			918 => "0000011000011000000100",
			919 => "0000000000111001111001",
			920 => "0000000000111001111001",
			921 => "0011110011101100000100",
			922 => "0000000000111001111001",
			923 => "0010101101101100000100",
			924 => "0000000000111001111001",
			925 => "0000000000111001111001",
			926 => "0011011010100101000100",
			927 => "0001011110010100110000",
			928 => "0011011011101100011100",
			929 => "0001111111011000001000",
			930 => "0001010001011000000100",
			931 => "0000000000111101011101",
			932 => "0000000000111101011101",
			933 => "0001111101001000001100",
			934 => "0001011001000000001000",
			935 => "0001011100101100000100",
			936 => "0000000000111101011101",
			937 => "0000000000111101011101",
			938 => "0000000000111101011101",
			939 => "0000111001010000000100",
			940 => "0000000000111101011101",
			941 => "0000000000111101011101",
			942 => "0000001100000100001100",
			943 => "0011100001010100001000",
			944 => "0001110101111000000100",
			945 => "0000000000111101011101",
			946 => "0000000000111101011101",
			947 => "0000000000111101011101",
			948 => "0001001001010100000100",
			949 => "0000000000111101011101",
			950 => "0000000000111101011101",
			951 => "0011011110011000001100",
			952 => "0001001110111000000100",
			953 => "0000000000111101011101",
			954 => "0000010001110000000100",
			955 => "0000000000111101011101",
			956 => "0000000000111101011101",
			957 => "0010001111111100000100",
			958 => "0000000000111101011101",
			959 => "0000000000111101011101",
			960 => "0001101111111000001000",
			961 => "0011000011010000000100",
			962 => "0000000000111101011101",
			963 => "0000000000111101011101",
			964 => "0010110101011100001100",
			965 => "0010110111011100001000",
			966 => "0001101111010100000100",
			967 => "0000000000111101011101",
			968 => "0000000000111101011101",
			969 => "0000000000111101011101",
			970 => "0001000001010100001100",
			971 => "0010000000110000001000",
			972 => "0010100000111100000100",
			973 => "0000000000111101011101",
			974 => "0000000000111101011101",
			975 => "0000000000111101011101",
			976 => "0011101100100000001000",
			977 => "0000010111100100000100",
			978 => "0000000000111101011101",
			979 => "0000000000111101011101",
			980 => "0001110001011000000100",
			981 => "0000000000111101011101",
			982 => "0000000000111101011101",
			983 => "0001000110101100000100",
			984 => "1111111000111111010001",
			985 => "0000000001110100101000",
			986 => "0010011001000100000100",
			987 => "0000001000111111010001",
			988 => "0000101000101100001000",
			989 => "0010011101101000000100",
			990 => "0000000000111111010001",
			991 => "1111111000111111010001",
			992 => "0010101010011100001100",
			993 => "0010000101011100000100",
			994 => "0000000000111111010001",
			995 => "0011010111011100000100",
			996 => "0000001000111111010001",
			997 => "0000000000111111010001",
			998 => "0000001011011000001000",
			999 => "0011101010011000000100",
			1000 => "0000000000111111010001",
			1001 => "1111111000111111010001",
			1002 => "0011110010000000000100",
			1003 => "0000000000111111010001",
			1004 => "0000001000111111010001",
			1005 => "0000111001000000000100",
			1006 => "1111111000111111010001",
			1007 => "0000010001100100000100",
			1008 => "0000001000111111010001",
			1009 => "0010100001101000000100",
			1010 => "0000000000111111010001",
			1011 => "0000000000111111010001",
			1012 => "0001011010011100010100",
			1013 => "0001001001010000001100",
			1014 => "0001011110111000000100",
			1015 => "1111111001000001011101",
			1016 => "0000111011111000000100",
			1017 => "0000000001000001011101",
			1018 => "1111111001000001011101",
			1019 => "0000111011111000000100",
			1020 => "0000001001000001011101",
			1021 => "1111111001000001011101",
			1022 => "0010111010000100110000",
			1023 => "0000101010000000101100",
			1024 => "0001010001011100010100",
			1025 => "0010011001000100000100",
			1026 => "0000001001000001011101",
			1027 => "0000001110101100001000",
			1028 => "0011101111100100000100",
			1029 => "0000000001000001011101",
			1030 => "1111111001000001011101",
			1031 => "0010110111011100000100",
			1032 => "0000001001000001011101",
			1033 => "0000000001000001011101",
			1034 => "0011110011101100010000",
			1035 => "0010000101101100001000",
			1036 => "0011101111100100000100",
			1037 => "0000001001000001011101",
			1038 => "0000001001000001011101",
			1039 => "0000001011110100000100",
			1040 => "0000000001000001011101",
			1041 => "0000001001000001011101",
			1042 => "0011010101011100000100",
			1043 => "0000001001000001011101",
			1044 => "0000001001000001011101",
			1045 => "1111111001000001011101",
			1046 => "1111111001000001011101",
			1047 => "0011011010100100111100",
			1048 => "0000111000100000101000",
			1049 => "0001111000000100001000",
			1050 => "0001010001011000000100",
			1051 => "0000000001000100111001",
			1052 => "0000000001000100111001",
			1053 => "0001111000111000001100",
			1054 => "0010011001000100001000",
			1055 => "0011101101000100000100",
			1056 => "0000000001000100111001",
			1057 => "0000000001000100111001",
			1058 => "0000000001000100111001",
			1059 => "0000000111001100010000",
			1060 => "0000100001111000001000",
			1061 => "0001101010110100000100",
			1062 => "0000000001000100111001",
			1063 => "0000000001000100111001",
			1064 => "0000111000101000000100",
			1065 => "0000000001000100111001",
			1066 => "0000000001000100111001",
			1067 => "0000000001000100111001",
			1068 => "0010010011000000001100",
			1069 => "0011101010110100000100",
			1070 => "0000000001000100111001",
			1071 => "0001100110100000000100",
			1072 => "0000000001000100111001",
			1073 => "0000000001000100111001",
			1074 => "0010001111111100000100",
			1075 => "0000000001000100111001",
			1076 => "0000000001000100111001",
			1077 => "0000010001110000001000",
			1078 => "0010001001000100000100",
			1079 => "0000000001000100111001",
			1080 => "0000000001000100111001",
			1081 => "0010100000111000100000",
			1082 => "0000100001100000001100",
			1083 => "0001111100010000001000",
			1084 => "0000000100111000000100",
			1085 => "0000000001000100111001",
			1086 => "0000000001000100111001",
			1087 => "0000000001000100111001",
			1088 => "0010110011010000001000",
			1089 => "0010010110000000000100",
			1090 => "0000000001000100111001",
			1091 => "0000000001000100111001",
			1092 => "0001100010011000000100",
			1093 => "0000000001000100111001",
			1094 => "0001100110110000000100",
			1095 => "0000000001000100111001",
			1096 => "0000000001000100111001",
			1097 => "0010101101101100001000",
			1098 => "0011110111101000000100",
			1099 => "0000000001000100111001",
			1100 => "0000000001000100111001",
			1101 => "0000000001000100111001",
			1102 => "0010001001000101000000",
			1103 => "0010101011000000010100",
			1104 => "0001110011001000001100",
			1105 => "0001111010000100000100",
			1106 => "0000000001000111110101",
			1107 => "0010011100101000000100",
			1108 => "0000000001000111110101",
			1109 => "0000000001000111110101",
			1110 => "0010011010000100000100",
			1111 => "0000000001000111110101",
			1112 => "0000000001000111110101",
			1113 => "0011010111011100100100",
			1114 => "0010110111011100001100",
			1115 => "0010000011010000000100",
			1116 => "0000000001000111110101",
			1117 => "0000000111000100000100",
			1118 => "0000000001000111110101",
			1119 => "0000000001000111110101",
			1120 => "0001011010100000010000",
			1121 => "0011100010011100001000",
			1122 => "0011000101011100000100",
			1123 => "0000000001000111110101",
			1124 => "0000000001000111110101",
			1125 => "0000000100111100000100",
			1126 => "0000000001000111110101",
			1127 => "0000000001000111110101",
			1128 => "0010001111111100000100",
			1129 => "0000000001000111110101",
			1130 => "0000000001000111110101",
			1131 => "0000111010011100000100",
			1132 => "0000000001000111110101",
			1133 => "0000000001000111110101",
			1134 => "0011011011101100000100",
			1135 => "0000000001000111110101",
			1136 => "0011111110111100000100",
			1137 => "0000000001000111110101",
			1138 => "0011101010011000000100",
			1139 => "0000000001000111110101",
			1140 => "0001011010001100001100",
			1141 => "0011000110000000000100",
			1142 => "0000000001000111110101",
			1143 => "0011001101101000000100",
			1144 => "0000000001000111110101",
			1145 => "0000000001000111110101",
			1146 => "0011000011000000000100",
			1147 => "0000000001000111110101",
			1148 => "0000000001000111110101",
			1149 => "0001010001011000000100",
			1150 => "1111111001001001100001",
			1151 => "0000011101000000101100",
			1152 => "0000111001111100101000",
			1153 => "0010100001101000011100",
			1154 => "0011011010100100001100",
			1155 => "0000001011001000001000",
			1156 => "0010011001000100000100",
			1157 => "0000001001001001100001",
			1158 => "0000001001001001100001",
			1159 => "0000000001001001100001",
			1160 => "0010110101011100001000",
			1161 => "0001010001010100000100",
			1162 => "0000000001001001100001",
			1163 => "1111111001001001100001",
			1164 => "0000000100110100000100",
			1165 => "0000000001001001100001",
			1166 => "0000001001001001100001",
			1167 => "0000000000100100000100",
			1168 => "0000001001001001100001",
			1169 => "0001011010011000000100",
			1170 => "0000001001001001100001",
			1171 => "0000001001001001100001",
			1172 => "1111111001001001100001",
			1173 => "0001111111101000000100",
			1174 => "0000000001001001100001",
			1175 => "1111111001001001100001",
			1176 => "0001000110101100000100",
			1177 => "1111111001001011110101",
			1178 => "0011101010011000101100",
			1179 => "0011011010100100010100",
			1180 => "0000000010010000001100",
			1181 => "0001111000000000001000",
			1182 => "0010001111111100000100",
			1183 => "0000000001001011110101",
			1184 => "0000001001001011110101",
			1185 => "0000000001001011110101",
			1186 => "0010011101101000000100",
			1187 => "0000000001001011110101",
			1188 => "0000001001001011110101",
			1189 => "0001000001011000001000",
			1190 => "0001000100101100000100",
			1191 => "0000000001001011110101",
			1192 => "1111111001001011110101",
			1193 => "0000111110111000000100",
			1194 => "0000001001001011110101",
			1195 => "0000100111000000000100",
			1196 => "1111111001001011110101",
			1197 => "0011111001011100000100",
			1198 => "0000000001001011110101",
			1199 => "0000001001001011110101",
			1200 => "0001110110101100000100",
			1201 => "1111111001001011110101",
			1202 => "0000001011011000000100",
			1203 => "1111111001001011110101",
			1204 => "0000001001110100001100",
			1205 => "0011000101111000001000",
			1206 => "0000000001110100000100",
			1207 => "0000001001001011110101",
			1208 => "0000000001001011110101",
			1209 => "1111111001001011110101",
			1210 => "0001010001011100000100",
			1211 => "1111111001001011110101",
			1212 => "0000000001001011110101",
			1213 => "0001000110101100000100",
			1214 => "1111111001001101111001",
			1215 => "0011011010100100100000",
			1216 => "0000101000100100011100",
			1217 => "0011110001101100011000",
			1218 => "0001111000000000001100",
			1219 => "0000111000100000001000",
			1220 => "0001001100101100000100",
			1221 => "0000001001001101111001",
			1222 => "0000000001001101111001",
			1223 => "0000001001001101111001",
			1224 => "0000000010010000000100",
			1225 => "0000000001001101111001",
			1226 => "0011100000100000000100",
			1227 => "0000001001001101111001",
			1228 => "0000000001001101111001",
			1229 => "0000001001001101111001",
			1230 => "0000000001001101111001",
			1231 => "0010110101011100001000",
			1232 => "0010000101101100000100",
			1233 => "0000000001001101111001",
			1234 => "1111111001001101111001",
			1235 => "0010100000111100000100",
			1236 => "1111111001001101111001",
			1237 => "0000110000111100001000",
			1238 => "0001001011000000000100",
			1239 => "1111111001001101111001",
			1240 => "0000001001001101111001",
			1241 => "0000001001111000000100",
			1242 => "1111111001001101111001",
			1243 => "0011011001001000000100",
			1244 => "0000000001001101111001",
			1245 => "1111111001001101111001",
			1246 => "0001000110101100000100",
			1247 => "1111111001010000001101",
			1248 => "0010001001000100101100",
			1249 => "0010101100110100100100",
			1250 => "0001101010011000010100",
			1251 => "0000010111110000001000",
			1252 => "0011101010100000000100",
			1253 => "0000000001010000001101",
			1254 => "0000000001010000001101",
			1255 => "0010010110000000000100",
			1256 => "0000001001010000001101",
			1257 => "0001101111000000000100",
			1258 => "0000000001010000001101",
			1259 => "0000000001010000001101",
			1260 => "0000000100011000000100",
			1261 => "1111111001010000001101",
			1262 => "0000000011100000001000",
			1263 => "0001011111100000000100",
			1264 => "0000001001010000001101",
			1265 => "0000000001010000001101",
			1266 => "0000000001010000001101",
			1267 => "0010011000000100000100",
			1268 => "0000001001010000001101",
			1269 => "0000000001010000001101",
			1270 => "0011001100101000000100",
			1271 => "0000000001010000001101",
			1272 => "0001011010001100001100",
			1273 => "0001111011111000000100",
			1274 => "1111111001010000001101",
			1275 => "0000001001110100000100",
			1276 => "0000000001010000001101",
			1277 => "0000000001010000001101",
			1278 => "0010101101101100000100",
			1279 => "0000000001010000001101",
			1280 => "0011011001001000000100",
			1281 => "0000000001010000001101",
			1282 => "0000000001010000001101",
			1283 => "0010110111011100010100",
			1284 => "0001011110010100001100",
			1285 => "0001011110001100001000",
			1286 => "0001010001011000000100",
			1287 => "0000000001010010111001",
			1288 => "0000000001010010111001",
			1289 => "0000000001010010111001",
			1290 => "0001010001011100000100",
			1291 => "0000000001010010111001",
			1292 => "0000000001010010111001",
			1293 => "0010001001001100000100",
			1294 => "0000000001010010111001",
			1295 => "0011000101011100010100",
			1296 => "0010011001000100000100",
			1297 => "0000000001010010111001",
			1298 => "0001111101001000001000",
			1299 => "0011111001111100000100",
			1300 => "0000000001010010111001",
			1301 => "0000000001010010111001",
			1302 => "0001100001100000000100",
			1303 => "0000000001010010111001",
			1304 => "0000000001010010111001",
			1305 => "0000110000111100010000",
			1306 => "0001001000100000001100",
			1307 => "0010110101010100001000",
			1308 => "0011110110100000000100",
			1309 => "0000000001010010111001",
			1310 => "0000000001010010111001",
			1311 => "0000000001010010111001",
			1312 => "0000000001010010111001",
			1313 => "0001111000101000001100",
			1314 => "0010100001101000001000",
			1315 => "0001000001011000000100",
			1316 => "0000000001010010111001",
			1317 => "0000000001010010111001",
			1318 => "0000000001010010111001",
			1319 => "0011011001001000001000",
			1320 => "0000111001111100000100",
			1321 => "0000000001010010111001",
			1322 => "0000000001010010111001",
			1323 => "0000000111101100000100",
			1324 => "0000000001010010111001",
			1325 => "0000000001010010111001",
			1326 => "0000101011100001010100",
			1327 => "0001011101111100111100",
			1328 => "0010101010011100110100",
			1329 => "0010000101011100011000",
			1330 => "0001110110101100010000",
			1331 => "0010111010100100001000",
			1332 => "0011011101000000000100",
			1333 => "0000000001010101110101",
			1334 => "0000000001010101110101",
			1335 => "0010011001000100000100",
			1336 => "0000000001010101110101",
			1337 => "1111111001010101110101",
			1338 => "0000000101000100000100",
			1339 => "0000000001010101110101",
			1340 => "0000000001010101110101",
			1341 => "0000000000001100001100",
			1342 => "0001111000000000001000",
			1343 => "0001010000111000000100",
			1344 => "0000000001010101110101",
			1345 => "0000001001010101110101",
			1346 => "1111111001010101110101",
			1347 => "0011100010011100001000",
			1348 => "0000001011110100000100",
			1349 => "0000001001010101110101",
			1350 => "0000000001010101110101",
			1351 => "0000001011110100000100",
			1352 => "0000000001010101110101",
			1353 => "0000001001010101110101",
			1354 => "0010001111111100000100",
			1355 => "0000000001010101110101",
			1356 => "1111111001010101110101",
			1357 => "0010000101101100001100",
			1358 => "0010010011000000000100",
			1359 => "0000001001010101110101",
			1360 => "0001101111000100000100",
			1361 => "0000000001010101110101",
			1362 => "0000000001010101110101",
			1363 => "0000001011110100000100",
			1364 => "1111111001010101110101",
			1365 => "0000111001111100000100",
			1366 => "0000001001010101110101",
			1367 => "0000000001010101110101",
			1368 => "0000111001000000000100",
			1369 => "1111111001010101110101",
			1370 => "0000011101000000000100",
			1371 => "0000000001010101110101",
			1372 => "0000000001010101110101",
			1373 => "0011101010011000111100",
			1374 => "0010010110000000011000",
			1375 => "0001011100110100010100",
			1376 => "0001111000000100010000",
			1377 => "0001011110111000001100",
			1378 => "0011001010100100001000",
			1379 => "0001011100010000000100",
			1380 => "0000000001011001101001",
			1381 => "0000000001011001101001",
			1382 => "0000000001011001101001",
			1383 => "0000001001011001101001",
			1384 => "0000000001011001101001",
			1385 => "0000001001011001101001",
			1386 => "0001100101110000000100",
			1387 => "1111111001011001101001",
			1388 => "0000100010111100010100",
			1389 => "0001101010011000001100",
			1390 => "0010001001000100001000",
			1391 => "0011000101011100000100",
			1392 => "0000000001011001101001",
			1393 => "0000000001011001101001",
			1394 => "1111111001011001101001",
			1395 => "0000010110010000000100",
			1396 => "0000000001011001101001",
			1397 => "1111111001011001101001",
			1398 => "0010110101101100001000",
			1399 => "0000101011010100000100",
			1400 => "0000001001011001101001",
			1401 => "0000000001011001101001",
			1402 => "0000000001011001101001",
			1403 => "0001110110101100001100",
			1404 => "0000111111101000001000",
			1405 => "0000111101001000000100",
			1406 => "0000000001011001101001",
			1407 => "0000000001011001101001",
			1408 => "1111111001011001101001",
			1409 => "0010001001000100011100",
			1410 => "0000000101100100000100",
			1411 => "1111111001011001101001",
			1412 => "0000101011100000001100",
			1413 => "0001001100001100001000",
			1414 => "0000111111101000000100",
			1415 => "0000000001011001101001",
			1416 => "0000001001011001101001",
			1417 => "0000000001011001101001",
			1418 => "0001111011111000000100",
			1419 => "0000000001011001101001",
			1420 => "0010000101101100000100",
			1421 => "0000000001011001101001",
			1422 => "0000000001011001101001",
			1423 => "0000110000111000001100",
			1424 => "0011000110000000000100",
			1425 => "1111111001011001101001",
			1426 => "0011001101101000000100",
			1427 => "0000000001011001101001",
			1428 => "0000000001011001101001",
			1429 => "0010101101101100000100",
			1430 => "0000000001011001101001",
			1431 => "0000011000011000000100",
			1432 => "0000000001011001101001",
			1433 => "0000000001011001101001",
			1434 => "0001010001011000000100",
			1435 => "1111111001011100000111",
			1436 => "0010011001000100001000",
			1437 => "0000001110101100000100",
			1438 => "0000001001011100000111",
			1439 => "0000000001011100000111",
			1440 => "0001011101111100100100",
			1441 => "0010101010011100011000",
			1442 => "0000111000100000001100",
			1443 => "0001001000100000001000",
			1444 => "0001011100001100000100",
			1445 => "0000000001011100000111",
			1446 => "1111111001011100000111",
			1447 => "0000000001011100000111",
			1448 => "0010001111001000001000",
			1449 => "0010110101010100000100",
			1450 => "0000001001011100000111",
			1451 => "0000000001011100000111",
			1452 => "1111111001011100000111",
			1453 => "0010001111111100000100",
			1454 => "0000000001011100000111",
			1455 => "0001100110110000000100",
			1456 => "1111111001011100000111",
			1457 => "0000000001011100000111",
			1458 => "0010000101101100001100",
			1459 => "0010010011000000000100",
			1460 => "0000001001011100000111",
			1461 => "0001000010111000000100",
			1462 => "0000000001011100000111",
			1463 => "0000000001011100000111",
			1464 => "0000001011110100000100",
			1465 => "1111111001011100000111",
			1466 => "0010101101101100001000",
			1467 => "0001001100011100000100",
			1468 => "0000000001011100000111",
			1469 => "0000001001011100000111",
			1470 => "0000011000011000000100",
			1471 => "0000000001011100000111",
			1472 => "0000000001011100000111",
			1473 => "0001001001010000010000",
			1474 => "0001011010011100001100",
			1475 => "0001000110101100000100",
			1476 => "1111111001011101111001",
			1477 => "0010011101101000000100",
			1478 => "0000000001011101111001",
			1479 => "1111111001011101111001",
			1480 => "0000000001011101111001",
			1481 => "0011011001001000100000",
			1482 => "0001000000100000011100",
			1483 => "0010101100110100010000",
			1484 => "0011010101010100001100",
			1485 => "0001111000000100000100",
			1486 => "0000001001011101111001",
			1487 => "0000001110101100000100",
			1488 => "0000000001011101111001",
			1489 => "0000001001011101111001",
			1490 => "1111111001011101111001",
			1491 => "0010001001000100000100",
			1492 => "0000001001011101111001",
			1493 => "0010011000000100000100",
			1494 => "0000000001011101111001",
			1495 => "0000001001011101111001",
			1496 => "1111111001011101111001",
			1497 => "0000010011110000001000",
			1498 => "0000100011111100000100",
			1499 => "1111111001011101111001",
			1500 => "0000001001011101111001",
			1501 => "1111111001011101111001",
			1502 => "0010000101101100110000",
			1503 => "0010011010000100011000",
			1504 => "0001001100101100001100",
			1505 => "0000000111001100001000",
			1506 => "0001000110101100000100",
			1507 => "0000000001100000100101",
			1508 => "0000000001100000100101",
			1509 => "0000000001100000100101",
			1510 => "0010101100110100001000",
			1511 => "0011111010110100000100",
			1512 => "0000000001100000100101",
			1513 => "0000000001100000100101",
			1514 => "0000000001100000100101",
			1515 => "0010010011000000001000",
			1516 => "0011001001001000000100",
			1517 => "0000000001100000100101",
			1518 => "0000000001100000100101",
			1519 => "0000101000001000001100",
			1520 => "0010010101111000000100",
			1521 => "0000000001100000100101",
			1522 => "0000010111110000000100",
			1523 => "0000000001100000100101",
			1524 => "0000000001100000100101",
			1525 => "0000000001100000100101",
			1526 => "0000001101010000010000",
			1527 => "0001100111010100001100",
			1528 => "0010011101101000001000",
			1529 => "0000001110100100000100",
			1530 => "0000000001100000100101",
			1531 => "0000000001100000100101",
			1532 => "0000000001100000100101",
			1533 => "0000000001100000100101",
			1534 => "0011011010100100001000",
			1535 => "0001011110001100000100",
			1536 => "0000000001100000100101",
			1537 => "0000000001100000100101",
			1538 => "0001011010001100001000",
			1539 => "0000110000111000000100",
			1540 => "0000000001100000100101",
			1541 => "0000000001100000100101",
			1542 => "0010101101101100000100",
			1543 => "0000000001100000100101",
			1544 => "0000000001100000100101",
			1545 => "0011011010100100101100",
			1546 => "0000111000100000011100",
			1547 => "0001111000000100001000",
			1548 => "0001010001011000000100",
			1549 => "0000000001100011010001",
			1550 => "0000001001100011010001",
			1551 => "0000100001111000000100",
			1552 => "1111111001100011010001",
			1553 => "0000000111001100001100",
			1554 => "0000001011011100000100",
			1555 => "0000000001100011010001",
			1556 => "0001001001010100000100",
			1557 => "0000000001100011010001",
			1558 => "0000001001100011010001",
			1559 => "1111111001100011010001",
			1560 => "0001000001011000001000",
			1561 => "0010000101011100000100",
			1562 => "0000000001100011010001",
			1563 => "0000001001100011010001",
			1564 => "0001011010100000000100",
			1565 => "0000000001100011010001",
			1566 => "0000001001100011010001",
			1567 => "0010110101011100010000",
			1568 => "0010110011010000001000",
			1569 => "0000011000011000000100",
			1570 => "0000000001100011010001",
			1571 => "0000000001100011010001",
			1572 => "0000010001110000000100",
			1573 => "0000000001100011010001",
			1574 => "1111111001100011010001",
			1575 => "0000110000111100001000",
			1576 => "0001001011000000000100",
			1577 => "0000000001100011010001",
			1578 => "0000001001100011010001",
			1579 => "0010101100001100000100",
			1580 => "1111111001100011010001",
			1581 => "0010001111001000001000",
			1582 => "0001000010001100000100",
			1583 => "0000000001100011010001",
			1584 => "0000000001100011010001",
			1585 => "0000011000011000000100",
			1586 => "0000000001100011010001",
			1587 => "0000000001100011010001",
			1588 => "0011101101000100111000",
			1589 => "0011000101010100010000",
			1590 => "0011010110110100001000",
			1591 => "0000010001110000000100",
			1592 => "0000000001100101101101",
			1593 => "0000000001100101101101",
			1594 => "0001010001011000000100",
			1595 => "0000000001100101101101",
			1596 => "0000001001100101101101",
			1597 => "0000001100000100001000",
			1598 => "0010000101011100000100",
			1599 => "0000000001100101101101",
			1600 => "1111111001100101101101",
			1601 => "0011011011101100001000",
			1602 => "0010011010000100000100",
			1603 => "1111111001100101101101",
			1604 => "0000001001100101101101",
			1605 => "0000010001110000001000",
			1606 => "0010110101010100000100",
			1607 => "0000001001100101101101",
			1608 => "0000000001100101101101",
			1609 => "0011101101111100001000",
			1610 => "0000100100000100000100",
			1611 => "0000001001100101101101",
			1612 => "0000000001100101101101",
			1613 => "0011001100101000000100",
			1614 => "0000000001100101101101",
			1615 => "0000000001100101101101",
			1616 => "0011001001001000001100",
			1617 => "0010000101011100001000",
			1618 => "0010001001001100000100",
			1619 => "0000000001100101101101",
			1620 => "0000000001100101101101",
			1621 => "1111111001100101101101",
			1622 => "0000011101000000001000",
			1623 => "0000110010010100000100",
			1624 => "0000000001100101101101",
			1625 => "0000000001100101101101",
			1626 => "0000000001100101101101",
			1627 => "0000111011000000010100",
			1628 => "0001111000000100001000",
			1629 => "0001010001011000000100",
			1630 => "0000000001101000001001",
			1631 => "0000000001101000001001",
			1632 => "0000011001100100001000",
			1633 => "0000000011100000000100",
			1634 => "0000000001101000001001",
			1635 => "0000000001101000001001",
			1636 => "0000000001101000001001",
			1637 => "0010000101101100011000",
			1638 => "0000000011011100010100",
			1639 => "0010010011000000001100",
			1640 => "0010011010000100001000",
			1641 => "0010011101101000000100",
			1642 => "0000000001101000001001",
			1643 => "0000000001101000001001",
			1644 => "0000000001101000001001",
			1645 => "0000101000001000000100",
			1646 => "0000000001101000001001",
			1647 => "0000000001101000001001",
			1648 => "0000000001101000001001",
			1649 => "0011111110111100010000",
			1650 => "0010101001000000000100",
			1651 => "0000000001101000001001",
			1652 => "0000100100001000000100",
			1653 => "0000000001101000001001",
			1654 => "0000100010101000000100",
			1655 => "0000000001101000001001",
			1656 => "0000000001101000001001",
			1657 => "0011101010011000000100",
			1658 => "0000000001101000001001",
			1659 => "0011110011101100000100",
			1660 => "0000000001101000001001",
			1661 => "0000000011111000001000",
			1662 => "0000110101001000000100",
			1663 => "0000000001101000001001",
			1664 => "0000000001101000001001",
			1665 => "0000000001101000001001",
			1666 => "0011011010100100110000",
			1667 => "0000111011000000011100",
			1668 => "0001111000000100001000",
			1669 => "0001010001011000000100",
			1670 => "0000000001101010111101",
			1671 => "0000000001101010111101",
			1672 => "0000011001100100001000",
			1673 => "0010010110000000000100",
			1674 => "0000000001101010111101",
			1675 => "0000000001101010111101",
			1676 => "0011000101011100000100",
			1677 => "0000000001101010111101",
			1678 => "0010011010000100000100",
			1679 => "0000000001101010111101",
			1680 => "0000000001101010111101",
			1681 => "0010010011000000001100",
			1682 => "0010000101101100001000",
			1683 => "0011000101011100000100",
			1684 => "0000000001101010111101",
			1685 => "0000000001101010111101",
			1686 => "0000000001101010111101",
			1687 => "0000001101001100000100",
			1688 => "0000000001101010111101",
			1689 => "0000000001101010111101",
			1690 => "0010110101011100010000",
			1691 => "0000010001110000000100",
			1692 => "0000000001101010111101",
			1693 => "0010110011010000001000",
			1694 => "0001011011111000000100",
			1695 => "0000000001101010111101",
			1696 => "0000000001101010111101",
			1697 => "0000000001101010111101",
			1698 => "0010100000111100000100",
			1699 => "0000000001101010111101",
			1700 => "0000111110111000001000",
			1701 => "0001000110011100000100",
			1702 => "0000000001101010111101",
			1703 => "0000000001101010111101",
			1704 => "0000100010111100000100",
			1705 => "0000000001101010111101",
			1706 => "0010101101101100001000",
			1707 => "0000001011111100000100",
			1708 => "0000000001101010111101",
			1709 => "0000000001101010111101",
			1710 => "0000000001101010111101",
			1711 => "0011101010011000111100",
			1712 => "0000000111101000011000",
			1713 => "0010011001000100001000",
			1714 => "0001010001011000000100",
			1715 => "0000000001101110001001",
			1716 => "0000000001101110001001",
			1717 => "0011000101010100001000",
			1718 => "0011101110010100000100",
			1719 => "0000000001101110001001",
			1720 => "0000000001101110001001",
			1721 => "0010000101011100000100",
			1722 => "0000000001101110001001",
			1723 => "0000000001101110001001",
			1724 => "0001011100110100001100",
			1725 => "0001101110000000001000",
			1726 => "0000111111101000000100",
			1727 => "0000000001101110001001",
			1728 => "0000000001101110001001",
			1729 => "0000000001101110001001",
			1730 => "0011010111011100001100",
			1731 => "0001111101001000001000",
			1732 => "0010001001001100000100",
			1733 => "0000000001101110001001",
			1734 => "0000000001101110001001",
			1735 => "0000000001101110001001",
			1736 => "0000100010111100000100",
			1737 => "0000000001101110001001",
			1738 => "0001111011111000000100",
			1739 => "0000000001101110001001",
			1740 => "0000000001101110001001",
			1741 => "0000001011011000001100",
			1742 => "0001010010001100001000",
			1743 => "0001111001010000000100",
			1744 => "0000000001101110001001",
			1745 => "0000000001101110001001",
			1746 => "0000000001101110001001",
			1747 => "0000000111110100010000",
			1748 => "0000111011000000001000",
			1749 => "0000101000100100000100",
			1750 => "0000000001101110001001",
			1751 => "0000000001101110001001",
			1752 => "0000111001111100000100",
			1753 => "0000000001101110001001",
			1754 => "0000000001101110001001",
			1755 => "0001011111100000001000",
			1756 => "0000111001000000000100",
			1757 => "0000000001101110001001",
			1758 => "0000000001101110001001",
			1759 => "0000111010100000000100",
			1760 => "0000000001101110001001",
			1761 => "0000000001101110001001",
			1762 => "0001001001010000010000",
			1763 => "0001011010011100001100",
			1764 => "0001000110101100000100",
			1765 => "1111111001110000001101",
			1766 => "0010110111011100000100",
			1767 => "0000000001110000001101",
			1768 => "1111111001110000001101",
			1769 => "0000000001110000001101",
			1770 => "0011011001001000101000",
			1771 => "0001000000100000100100",
			1772 => "0010100000111000011000",
			1773 => "0011011010100100001100",
			1774 => "0011101010011000001000",
			1775 => "0010110101010100000100",
			1776 => "0000001001110000001101",
			1777 => "0000001001110000001101",
			1778 => "0000001001110000001101",
			1779 => "0000000100111100001000",
			1780 => "0000111001000000000100",
			1781 => "0000000001110000001101",
			1782 => "1111111001110000001101",
			1783 => "0000001001110000001101",
			1784 => "0011000110000000001000",
			1785 => "0010100001101000000100",
			1786 => "0000001001110000001101",
			1787 => "0000001001110000001101",
			1788 => "0000001001110000001101",
			1789 => "1111111001110000001101",
			1790 => "0000010011110000001000",
			1791 => "0011110010001000000100",
			1792 => "1111111001110000001101",
			1793 => "0000001001110000001101",
			1794 => "1111111001110000001101",
			1795 => "0001010001010100101100",
			1796 => "0001111000000100001000",
			1797 => "0001011110111000000100",
			1798 => "0000000001110010110001",
			1799 => "0000000001110010110001",
			1800 => "0000000000010000001100",
			1801 => "0010011001000100000100",
			1802 => "0000000001110010110001",
			1803 => "0000011001100100000100",
			1804 => "0000000001110010110001",
			1805 => "0000000001110010110001",
			1806 => "0000100100110100001100",
			1807 => "0011111010011000000100",
			1808 => "0000000001110010110001",
			1809 => "0001001001010100000100",
			1810 => "0000000001110010110001",
			1811 => "0000000001110010110001",
			1812 => "0000011001100100000100",
			1813 => "0000000001110010110001",
			1814 => "0010101010011100000100",
			1815 => "0000000001110010110001",
			1816 => "0000000001110010110001",
			1817 => "0010001111111100001100",
			1818 => "0000111010011100000100",
			1819 => "0000000001110010110001",
			1820 => "0000111100110100000100",
			1821 => "0000000001110010110001",
			1822 => "0000000001110010110001",
			1823 => "0001101010110100000100",
			1824 => "0000000001110010110001",
			1825 => "0000001011011100000100",
			1826 => "0000000001110010110001",
			1827 => "0011101010011000001000",
			1828 => "0001000010001100000100",
			1829 => "0000000001110010110001",
			1830 => "0000000001110010110001",
			1831 => "0000100101100100000100",
			1832 => "0000000001110010110001",
			1833 => "0011011001001000000100",
			1834 => "0000000001110010110001",
			1835 => "0000000001110010110001",
			1836 => "0001011110111000001000",
			1837 => "0001010001011000000100",
			1838 => "1111111001110100011101",
			1839 => "0000000001110100011101",
			1840 => "0011011001001000100100",
			1841 => "0000001001110100100000",
			1842 => "0010011001000100000100",
			1843 => "0000001001110100011101",
			1844 => "0000001110101100010000",
			1845 => "0011100100000000001000",
			1846 => "0001010001010100000100",
			1847 => "0000000001110100011101",
			1848 => "0000001001110100011101",
			1849 => "0011001100101000000100",
			1850 => "1111111001110100011101",
			1851 => "0000000001110100011101",
			1852 => "0000111001111100001000",
			1853 => "0010100000111000000100",
			1854 => "0000001001110100011101",
			1855 => "0000001001110100011101",
			1856 => "1111111001110100011101",
			1857 => "1111111001110100011101",
			1858 => "0000010001100100001000",
			1859 => "0000110001101100000100",
			1860 => "0000001001110100011101",
			1861 => "1111111001110100011101",
			1862 => "1111111001110100011101",
			1863 => "0010001001000100101100",
			1864 => "0010101100110100100100",
			1865 => "0010101010011100011100",
			1866 => "0001011110010100010100",
			1867 => "0000000111001100010000",
			1868 => "0011110100100100001000",
			1869 => "0010011001000100000100",
			1870 => "0000000001110110111001",
			1871 => "0000000001110110111001",
			1872 => "0000010110010000000100",
			1873 => "0000000001110110111001",
			1874 => "0000000001110110111001",
			1875 => "0000000001110110111001",
			1876 => "0011101001111100000100",
			1877 => "0000000001110110111001",
			1878 => "0000000001110110111001",
			1879 => "0010001111111100000100",
			1880 => "0000000001110110111001",
			1881 => "0000000001110110111001",
			1882 => "0010011000000100000100",
			1883 => "0000000001110110111001",
			1884 => "0000000001110110111001",
			1885 => "0010011101101000001000",
			1886 => "0010101011000000000100",
			1887 => "0000000001110110111001",
			1888 => "0000000001110110111001",
			1889 => "0001011010001100010100",
			1890 => "0001111000101000000100",
			1891 => "0000000001110110111001",
			1892 => "0000110001001000000100",
			1893 => "0000000001110110111001",
			1894 => "0000110001101000001000",
			1895 => "0001111001011000000100",
			1896 => "0000000001110110111001",
			1897 => "0000000001110110111001",
			1898 => "0000000001110110111001",
			1899 => "0010101101101100000100",
			1900 => "0000000001110110111001",
			1901 => "0000000001110110111001",
			1902 => "0011101010011000110000",
			1903 => "0000000010111100011100",
			1904 => "0001101010011000011000",
			1905 => "0010001001000100010000",
			1906 => "0000000100100000001100",
			1907 => "0011100100000000001000",
			1908 => "0010001111111100000100",
			1909 => "0000000001111001111101",
			1910 => "0000000001111001111101",
			1911 => "0000000001111001111101",
			1912 => "0000000001111001111101",
			1913 => "0010011001000100000100",
			1914 => "0000000001111001111101",
			1915 => "1111111001111001111101",
			1916 => "1111111001111001111101",
			1917 => "0011110100100100000100",
			1918 => "0000000001111001111101",
			1919 => "0000100100111100001100",
			1920 => "0011010011010000000100",
			1921 => "0000001001111001111101",
			1922 => "0001111011000000000100",
			1923 => "0000000001111001111101",
			1924 => "0000000001111001111101",
			1925 => "0000000001111001111101",
			1926 => "0010100001101000100100",
			1927 => "0010001111111100010100",
			1928 => "0000000011100000001000",
			1929 => "0000000100111100000100",
			1930 => "0000000001111001111101",
			1931 => "0000001001111001111101",
			1932 => "0001110110101100000100",
			1933 => "1111111001111001111101",
			1934 => "0000010001110000000100",
			1935 => "0000000001111001111101",
			1936 => "0000000001111001111101",
			1937 => "0011001001001000001000",
			1938 => "0010110101011100000100",
			1939 => "1111111001111001111101",
			1940 => "0000000001111001111101",
			1941 => "0000001010101000000100",
			1942 => "0000000001111001111101",
			1943 => "0000000001111001111101",
			1944 => "0010101101101100001000",
			1945 => "0000001110110100000100",
			1946 => "0000000001111001111101",
			1947 => "0000000001111001111101",
			1948 => "0011011001001000000100",
			1949 => "0000000001111001111101",
			1950 => "0000000001111001111101",
			1951 => "0011011110011000101000",
			1952 => "0001011110010100100000",
			1953 => "0001111000000100001100",
			1954 => "0011011101000000000100",
			1955 => "0000000001111101000001",
			1956 => "0001000110101100000100",
			1957 => "0000000001111101000001",
			1958 => "0000000001111101000001",
			1959 => "0001101010001100000100",
			1960 => "0000000001111101000001",
			1961 => "0010110011010000001000",
			1962 => "0011011011101100000100",
			1963 => "0000000001111101000001",
			1964 => "0000000001111101000001",
			1965 => "0001100011101100000100",
			1966 => "0000000001111101000001",
			1967 => "0000000001111101000001",
			1968 => "0010010011000000000100",
			1969 => "0000000001111101000001",
			1970 => "0000000001111101000001",
			1971 => "0000000000100100011000",
			1972 => "0001111100000000001000",
			1973 => "0000000100111000000100",
			1974 => "0000000001111101000001",
			1975 => "0000000001111101000001",
			1976 => "0000111011111000001000",
			1977 => "0010011101101000000100",
			1978 => "0000000001111101000001",
			1979 => "0000000001111101000001",
			1980 => "0010100000111000000100",
			1981 => "0000000001111101000001",
			1982 => "0000000001111101000001",
			1983 => "0011101110000000001000",
			1984 => "0011110001001100000100",
			1985 => "0000000001111101000001",
			1986 => "0000000001111101000001",
			1987 => "0011001001001000001100",
			1988 => "0010101000100000001000",
			1989 => "0010101011000000000100",
			1990 => "0000000001111101000001",
			1991 => "0000000001111101000001",
			1992 => "0000000001111101000001",
			1993 => "0000100111000100001100",
			1994 => "0000111001111100001000",
			1995 => "0010101001000000000100",
			1996 => "0000000001111101000001",
			1997 => "0000000001111101000001",
			1998 => "0000000001111101000001",
			1999 => "0000000001111101000001",
			2000 => "0000001011100000111100",
			2001 => "0000001100000100001100",
			2002 => "0011000101010100001000",
			2003 => "0001010001011000000100",
			2004 => "0000000001111111001101",
			2005 => "0000000001111111001101",
			2006 => "1111111001111111001101",
			2007 => "0001000010111000100100",
			2008 => "0011011011101100010000",
			2009 => "0010011010000100001100",
			2010 => "0001011001101100001000",
			2011 => "0001011110001100000100",
			2012 => "0000000001111111001101",
			2013 => "0000000001111111001101",
			2014 => "0000000001111111001101",
			2015 => "0000000001111111001101",
			2016 => "0000010001110000000100",
			2017 => "0000000001111111001101",
			2018 => "0010010011000000001000",
			2019 => "0000010111110000000100",
			2020 => "0000000001111111001101",
			2021 => "0000000001111111001101",
			2022 => "0000100010111100000100",
			2023 => "0000000001111111001101",
			2024 => "0000000001111111001101",
			2025 => "0001110001010000000100",
			2026 => "0000000001111111001101",
			2027 => "0000111001111100000100",
			2028 => "0000000001111111001101",
			2029 => "0000000001111111001101",
			2030 => "0001011111100000000100",
			2031 => "0000000001111111001101",
			2032 => "0010100001011100000100",
			2033 => "0000000001111111001101",
			2034 => "0000000001111111001101",
			2035 => "0011011010100100111100",
			2036 => "0011101010011000100100",
			2037 => "0000001110101100011000",
			2038 => "0011100101110000010100",
			2039 => "0001010000111000001100",
			2040 => "0001111000000100001000",
			2041 => "0001010001011000000100",
			2042 => "0000000010000010011001",
			2043 => "0000000010000010011001",
			2044 => "0000000010000010011001",
			2045 => "0010011101101000000100",
			2046 => "0000000010000010011001",
			2047 => "0000000010000010011001",
			2048 => "0000000010000010011001",
			2049 => "0001111000000000001000",
			2050 => "0010010101101100000100",
			2051 => "0000000010000010011001",
			2052 => "0000000010000010011001",
			2053 => "0000000010000010011001",
			2054 => "0001110110101100001100",
			2055 => "0000111111101000001000",
			2056 => "0000111101001000000100",
			2057 => "0000000010000010011001",
			2058 => "0000000010000010011001",
			2059 => "0000000010000010011001",
			2060 => "0000000101100100000100",
			2061 => "0000000010000010011001",
			2062 => "0010010110000000000100",
			2063 => "0000000010000010011001",
			2064 => "0000000010000010011001",
			2065 => "0000010001110000001000",
			2066 => "0010000101101100000100",
			2067 => "0000000010000010011001",
			2068 => "0000000010000010011001",
			2069 => "0010100000111000010100",
			2070 => "0010110011010000001000",
			2071 => "0001101001011100000100",
			2072 => "0000000010000010011001",
			2073 => "0000000010000010011001",
			2074 => "0001110001010000000100",
			2075 => "0000000010000010011001",
			2076 => "0011110100110000000100",
			2077 => "0000000010000010011001",
			2078 => "0000000010000010011001",
			2079 => "0010101101101100001100",
			2080 => "0011111110111100000100",
			2081 => "0000000010000010011001",
			2082 => "0011110111101000000100",
			2083 => "0000000010000010011001",
			2084 => "0000000010000010011001",
			2085 => "0000000010000010011001",
			2086 => "0000010001110000011100",
			2087 => "0001011110010100010100",
			2088 => "0011110100100100000100",
			2089 => "0000000010000101000101",
			2090 => "0000000011100000001000",
			2091 => "0010101101001000000100",
			2092 => "0000000010000101000101",
			2093 => "0000000010000101000101",
			2094 => "0001111001010000000100",
			2095 => "0000000010000101000101",
			2096 => "0000000010000101000101",
			2097 => "0001001100001100000100",
			2098 => "0000000010000101000101",
			2099 => "0000000010000101000101",
			2100 => "0001111000000100001000",
			2101 => "0001010001011000000100",
			2102 => "0000000010000101000101",
			2103 => "0000000010000101000101",
			2104 => "0010100000111000100100",
			2105 => "0010100000111100001100",
			2106 => "0011100010001100001000",
			2107 => "0001100010001100000100",
			2108 => "0000000010000101000101",
			2109 => "0000000010000101000101",
			2110 => "0000000010000101000101",
			2111 => "0010010011000000001100",
			2112 => "0000010111110000000100",
			2113 => "0000000010000101000101",
			2114 => "0001000011000100000100",
			2115 => "0000000010000101000101",
			2116 => "0000000010000101000101",
			2117 => "0011110011011000000100",
			2118 => "0000000010000101000101",
			2119 => "0001001100101100000100",
			2120 => "0000000010000101000101",
			2121 => "0000000010000101000101",
			2122 => "0010101101101100001000",
			2123 => "0010001111011000000100",
			2124 => "0000000010000101000101",
			2125 => "0000000010000101000101",
			2126 => "0000011000011000000100",
			2127 => "0000000010000101000101",
			2128 => "0000000010000101000101",
			2129 => "0011011010100101000000",
			2130 => "0001011110010100101000",
			2131 => "0001111000000100010100",
			2132 => "0001011110111000010000",
			2133 => "0000010001110000000100",
			2134 => "0000000010001000011001",
			2135 => "0000010111110000001000",
			2136 => "0010000101011100000100",
			2137 => "0000000010001000011001",
			2138 => "0000000010001000011001",
			2139 => "0000000010001000011001",
			2140 => "0000000010001000011001",
			2141 => "0001101010001100000100",
			2142 => "1111111010001000011001",
			2143 => "0000000111001100001100",
			2144 => "0000010110010000001000",
			2145 => "0000111000101000000100",
			2146 => "0000000010001000011001",
			2147 => "0000001010001000011001",
			2148 => "0000000010001000011001",
			2149 => "0000000010001000011001",
			2150 => "0001000001011000001000",
			2151 => "0000001011011100000100",
			2152 => "0000000010001000011001",
			2153 => "0000001010001000011001",
			2154 => "0001011010100000001000",
			2155 => "0001001110111000000100",
			2156 => "0000000010001000011001",
			2157 => "0000000010001000011001",
			2158 => "0010010011000000000100",
			2159 => "0000000010001000011001",
			2160 => "0000000010001000011001",
			2161 => "0000100010111100001100",
			2162 => "0000010001110000000100",
			2163 => "0000000010001000011001",
			2164 => "0011000011010000000100",
			2165 => "0000000010001000011001",
			2166 => "1111111010001000011001",
			2167 => "0010110101011100001100",
			2168 => "0010110111011100001000",
			2169 => "0010110011010000000100",
			2170 => "0000000010001000011001",
			2171 => "0000000010001000011001",
			2172 => "0000000010001000011001",
			2173 => "0000010001100100001100",
			2174 => "0000110000100000001000",
			2175 => "0001001100101100000100",
			2176 => "0000000010001000011001",
			2177 => "0000001010001000011001",
			2178 => "0000000010001000011001",
			2179 => "0010001010000100000100",
			2180 => "0000000010001000011001",
			2181 => "0000000010001000011001",
			2182 => "0010101011000000010100",
			2183 => "0001111000000100010000",
			2184 => "0001111010000100000100",
			2185 => "0000000010001011000101",
			2186 => "0011000111011100001000",
			2187 => "0011001010100100000100",
			2188 => "0000000010001011000101",
			2189 => "0000000010001011000101",
			2190 => "0000000010001011000101",
			2191 => "0000000010001011000101",
			2192 => "0010001001000100101000",
			2193 => "0011010011010000100000",
			2194 => "0001011110010100010000",
			2195 => "0011011011101100001000",
			2196 => "0010101000100000000100",
			2197 => "0000000010001011000101",
			2198 => "0000000010001011000101",
			2199 => "0000000000001100000100",
			2200 => "0000000010001011000101",
			2201 => "0000000010001011000101",
			2202 => "0011100101110000000100",
			2203 => "0000000010001011000101",
			2204 => "0000001011011100000100",
			2205 => "0000000010001011000101",
			2206 => "0010011010000100000100",
			2207 => "0000000010001011000101",
			2208 => "0000000010001011000101",
			2209 => "0001100010011000000100",
			2210 => "0000000010001011000101",
			2211 => "0000000010001011000101",
			2212 => "0011111110111100001000",
			2213 => "0001101101101100000100",
			2214 => "0000000010001011000101",
			2215 => "0000000010001011000101",
			2216 => "0011100101001000000100",
			2217 => "0000000010001011000101",
			2218 => "0010111100101000000100",
			2219 => "0000000010001011000101",
			2220 => "0011010101101100001000",
			2221 => "0000110000100000000100",
			2222 => "0000000010001011000101",
			2223 => "0000000010001011000101",
			2224 => "0000000010001011000101",
			2225 => "0000001011100001000100",
			2226 => "0010010110000000001100",
			2227 => "0001010001011000000100",
			2228 => "0000000010001101101001",
			2229 => "0011010110001100000100",
			2230 => "0000000010001101101001",
			2231 => "0000000010001101101001",
			2232 => "0000001110101100011100",
			2233 => "0011100100000000010100",
			2234 => "0001010001010100010000",
			2235 => "0001110110101100001000",
			2236 => "0000011001100100000100",
			2237 => "0000000010001101101001",
			2238 => "1111111010001101101001",
			2239 => "0000011001100000000100",
			2240 => "0000000010001101101001",
			2241 => "0000000010001101101001",
			2242 => "0000000010001101101001",
			2243 => "0001010010111000000100",
			2244 => "0000000010001101101001",
			2245 => "1111111010001101101001",
			2246 => "0011101011110000001100",
			2247 => "0011010111011100000100",
			2248 => "0000001010001101101001",
			2249 => "0001111101001000000100",
			2250 => "0000000010001101101001",
			2251 => "0000000010001101101001",
			2252 => "0000001101001100000100",
			2253 => "0000000010001101101001",
			2254 => "0001110110101100000100",
			2255 => "0000000010001101101001",
			2256 => "0011010101010100000100",
			2257 => "0000001010001101101001",
			2258 => "0000000010001101101001",
			2259 => "0001011111100000001000",
			2260 => "0000111001000000000100",
			2261 => "0000000010001101101001",
			2262 => "0000000010001101101001",
			2263 => "0000111010100000000100",
			2264 => "0000000010001101101001",
			2265 => "0000000010001101101001",
			2266 => "0001011010100001001100",
			2267 => "0011100010011100100100",
			2268 => "0001101111111000011100",
			2269 => "0010010110000000010000",
			2270 => "0000000011101100000100",
			2271 => "0000000010010000101101",
			2272 => "0000011001100100000100",
			2273 => "0000000010010000101101",
			2274 => "0001010001011000000100",
			2275 => "0000000010010000101101",
			2276 => "0000000010010000101101",
			2277 => "0001010001010100001000",
			2278 => "0001101010110100000100",
			2279 => "0000000010010000101101",
			2280 => "0000000010010000101101",
			2281 => "0000000010010000101101",
			2282 => "0000000101111100000100",
			2283 => "0000000010010000101101",
			2284 => "0000000010010000101101",
			2285 => "0000011001100100001100",
			2286 => "0000000100111100000100",
			2287 => "0000000010010000101101",
			2288 => "0010101011000000000100",
			2289 => "0000000010010000101101",
			2290 => "0000000010010000101101",
			2291 => "0011011110011000001100",
			2292 => "0000111011000000001000",
			2293 => "0000010111100100000100",
			2294 => "0000000010010000101101",
			2295 => "0000000010010000101101",
			2296 => "0000000010010000101101",
			2297 => "0010100000111000001100",
			2298 => "0010110011010000001000",
			2299 => "0010111010100100000100",
			2300 => "0000000010010000101101",
			2301 => "0000000010010000101101",
			2302 => "0000000010010000101101",
			2303 => "0000000010010000101101",
			2304 => "0010000101101100001000",
			2305 => "0001100000110100000100",
			2306 => "0000000010010000101101",
			2307 => "0000000010010000101101",
			2308 => "0001111000101000000100",
			2309 => "0000000010010000101101",
			2310 => "0010101101101100000100",
			2311 => "0000000010010000101101",
			2312 => "0000011000011000000100",
			2313 => "0000000010010000101101",
			2314 => "0000000010010000101101",
			2315 => "0001010001011000000100",
			2316 => "1111111010010010101001",
			2317 => "0010010110000000001100",
			2318 => "0001010010111000001000",
			2319 => "0001111000000100000100",
			2320 => "0000001010010010101001",
			2321 => "0000000010010010101001",
			2322 => "0000001010010010101001",
			2323 => "0000001110101100010000",
			2324 => "0010100000111100000100",
			2325 => "1111111010010010101001",
			2326 => "0011100100000000000100",
			2327 => "0000000010010010101001",
			2328 => "0001101111111000000100",
			2329 => "1111111010010010101001",
			2330 => "0000000010010010101001",
			2331 => "0010110111011100001000",
			2332 => "0001000000111100000100",
			2333 => "0000001010010010101001",
			2334 => "0000000010010010101001",
			2335 => "0010011010000100001000",
			2336 => "0000000101000100000100",
			2337 => "0000000010010010101001",
			2338 => "1111111010010010101001",
			2339 => "0011011010100100001000",
			2340 => "0001111001010100000100",
			2341 => "0000001010010010101001",
			2342 => "0000000010010010101001",
			2343 => "0011110011101100000100",
			2344 => "0000000010010010101001",
			2345 => "0000000010010010101001",
			2346 => "0001010001011000000100",
			2347 => "1111111010010100010101",
			2348 => "0000100111000100101100",
			2349 => "0010010110000000001000",
			2350 => "0000010111110000000100",
			2351 => "0000000010010100010101",
			2352 => "0000001010010100010101",
			2353 => "0000001101001100010100",
			2354 => "0011101111111000010000",
			2355 => "0001010001010100001000",
			2356 => "0001101010110100000100",
			2357 => "1111111010010100010101",
			2358 => "0000000010010100010101",
			2359 => "0010010011000000000100",
			2360 => "0000001010010100010101",
			2361 => "0000000010010100010101",
			2362 => "1111111010010100010101",
			2363 => "0001110110101100000100",
			2364 => "0000000010010100010101",
			2365 => "0011010011010000000100",
			2366 => "0000001010010100010101",
			2367 => "0011110011011000000100",
			2368 => "0000000010010100010101",
			2369 => "0000001010010100010101",
			2370 => "0001011010100000000100",
			2371 => "1111111010010100010101",
			2372 => "0000000010010100010101",
			2373 => "0001011010011100001100",
			2374 => "0001010001011000000100",
			2375 => "1111111010010110100001",
			2376 => "0011011110011000000100",
			2377 => "0000001010010110100001",
			2378 => "1111111010010110100001",
			2379 => "0011011001001000110000",
			2380 => "0000111001111100101100",
			2381 => "0000001110101100010100",
			2382 => "0011000101010100001000",
			2383 => "0011110010011100000100",
			2384 => "0000010010010110100001",
			2385 => "0000001010010110100001",
			2386 => "0011011110011000000100",
			2387 => "0000001010010110100001",
			2388 => "0010110101011100000100",
			2389 => "1111111010010110100001",
			2390 => "0000000010010110100001",
			2391 => "0011011010100100001100",
			2392 => "0011101010011000001000",
			2393 => "0010110101010100000100",
			2394 => "0000010010010110100001",
			2395 => "0000001010010110100001",
			2396 => "0000001010010110100001",
			2397 => "0010110101011100000100",
			2398 => "0000000010010110100001",
			2399 => "0000101101001100000100",
			2400 => "0000001010010110100001",
			2401 => "0000010010010110100001",
			2402 => "1111111010010110100001",
			2403 => "0010111101101000001000",
			2404 => "0001101000010100000100",
			2405 => "0000000010010110100001",
			2406 => "1111111010010110100001",
			2407 => "1111111010010110100001",
			2408 => "0001010001011000000100",
			2409 => "1111111010011000101101",
			2410 => "0010110111011100010100",
			2411 => "0001011110010100001100",
			2412 => "0000111011111000000100",
			2413 => "0000001010011000101101",
			2414 => "0011011011101100000100",
			2415 => "1111111010011000101101",
			2416 => "0000000010011000101101",
			2417 => "0001010001011100000100",
			2418 => "0000001010011000101101",
			2419 => "0000000010011000101101",
			2420 => "0001010001011100010100",
			2421 => "0000010001110000000100",
			2422 => "0000000010011000101101",
			2423 => "0000001011011100000100",
			2424 => "1111111010011000101101",
			2425 => "0011100010011100000100",
			2426 => "0000000010011000101101",
			2427 => "0001011100110100000100",
			2428 => "0000000010011000101101",
			2429 => "1111111010011000101101",
			2430 => "0010010011000000001000",
			2431 => "0010110101010100000100",
			2432 => "0000001010011000101101",
			2433 => "0000000010011000101101",
			2434 => "0011110011101100001100",
			2435 => "0011100000010100001000",
			2436 => "0000100010111100000100",
			2437 => "1111111010011000101101",
			2438 => "0000000010011000101101",
			2439 => "1111111010011000101101",
			2440 => "0000011101000000000100",
			2441 => "0000001010011000101101",
			2442 => "0000000010011000101101",
			2443 => "0011011010100100110000",
			2444 => "0000111000100000100000",
			2445 => "0001111000000100001000",
			2446 => "0001011110111000000100",
			2447 => "0000000010011100000001",
			2448 => "0000000010011100000001",
			2449 => "0000001011011100001100",
			2450 => "0010011001000100000100",
			2451 => "0000000010011100000001",
			2452 => "0011001001001000000100",
			2453 => "0000000010011100000001",
			2454 => "0000000010011100000001",
			2455 => "0000000111001100001000",
			2456 => "0001001001010000000100",
			2457 => "0000000010011100000001",
			2458 => "0000000010011100000001",
			2459 => "0000000010011100000001",
			2460 => "0001000001011000000100",
			2461 => "0000000010011100000001",
			2462 => "0010001111111100001000",
			2463 => "0010011010000100000100",
			2464 => "0000000010011100000001",
			2465 => "0000000010011100000001",
			2466 => "0000000010011100000001",
			2467 => "0010110101011100010100",
			2468 => "0010110011010000001000",
			2469 => "0001101001011100000100",
			2470 => "0000000010011100000001",
			2471 => "0000000010011100000001",
			2472 => "0001001000101000001000",
			2473 => "0010101011000000000100",
			2474 => "0000000010011100000001",
			2475 => "0000000010011100000001",
			2476 => "0000000010011100000001",
			2477 => "0010100000111100000100",
			2478 => "0000000010011100000001",
			2479 => "0001000000111000010100",
			2480 => "0000010011110000001000",
			2481 => "0010001001000100000100",
			2482 => "0000000010011100000001",
			2483 => "0000000010011100000001",
			2484 => "0001101111000100000100",
			2485 => "0000000010011100000001",
			2486 => "0001101000110100000100",
			2487 => "0000000010011100000001",
			2488 => "0000000010011100000001",
			2489 => "0011111110111100000100",
			2490 => "0000000010011100000001",
			2491 => "0011100000010100000100",
			2492 => "0000000010011100000001",
			2493 => "0011101100100000000100",
			2494 => "0000000010011100000001",
			2495 => "0000000010011100000001",
			2496 => "0001000110101100000100",
			2497 => "1111111010011110000101",
			2498 => "0011101111100100011000",
			2499 => "0010001001000100010100",
			2500 => "0011111111111000001100",
			2501 => "0010011001000100000100",
			2502 => "0000001010011110000101",
			2503 => "0001100101110000000100",
			2504 => "0000000010011110000101",
			2505 => "0000000010011110000101",
			2506 => "0000111001000000000100",
			2507 => "0000001010011110000101",
			2508 => "0000000010011110000101",
			2509 => "0000000010011110000101",
			2510 => "0000000010111100001000",
			2511 => "0011001100101000000100",
			2512 => "1111111010011110000101",
			2513 => "0000000010011110000101",
			2514 => "0011101010011000010000",
			2515 => "0011011010100100000100",
			2516 => "0000001010011110000101",
			2517 => "0001100000010100000100",
			2518 => "1111111010011110000101",
			2519 => "0001101101000100000100",
			2520 => "0000001010011110000101",
			2521 => "0000000010011110000101",
			2522 => "0000001011011000000100",
			2523 => "0000000010011110000101",
			2524 => "0001111101001000000100",
			2525 => "0000000010011110000101",
			2526 => "0000101010000000000100",
			2527 => "0000001010011110000101",
			2528 => "1111111010011110000101",
			2529 => "0000010110010000111100",
			2530 => "0010001001000100101100",
			2531 => "0000001011100000100100",
			2532 => "0000111000100000011100",
			2533 => "0001111000111000001100",
			2534 => "0001111000000100001000",
			2535 => "0001010001011000000100",
			2536 => "0000000010100001100001",
			2537 => "0000000010100001100001",
			2538 => "0000000010100001100001",
			2539 => "0001100010000000001000",
			2540 => "0000000000001100000100",
			2541 => "0000000010100001100001",
			2542 => "0000000010100001100001",
			2543 => "0001111001010100000100",
			2544 => "0000000010100001100001",
			2545 => "0000000010100001100001",
			2546 => "0011001001001000000100",
			2547 => "0000000010100001100001",
			2548 => "0000000010100001100001",
			2549 => "0001110100101100000100",
			2550 => "0000000010100001100001",
			2551 => "0000000010100001100001",
			2552 => "0001111000000000000100",
			2553 => "0000000010100001100001",
			2554 => "0010101001000000001000",
			2555 => "0010010101111000000100",
			2556 => "0000000010100001100001",
			2557 => "0000000010100001100001",
			2558 => "0000000010100001100001",
			2559 => "0001001100001100100000",
			2560 => "0000100100011000010000",
			2561 => "0010010110000000001100",
			2562 => "0000001110100100000100",
			2563 => "0000000010100001100001",
			2564 => "0001100101110000000100",
			2565 => "0000000010100001100001",
			2566 => "0000000010100001100001",
			2567 => "0000000010100001100001",
			2568 => "0000100111000100001100",
			2569 => "0010100000111100000100",
			2570 => "0000000010100001100001",
			2571 => "0001100010010100000100",
			2572 => "0000000010100001100001",
			2573 => "0000000010100001100001",
			2574 => "0000000010100001100001",
			2575 => "0001000001010100001000",
			2576 => "0001110100101100000100",
			2577 => "0000000010100001100001",
			2578 => "0000000010100001100001",
			2579 => "0011101100100000000100",
			2580 => "0000000010100001100001",
			2581 => "0001111110111000000100",
			2582 => "0000000010100001100001",
			2583 => "0000000010100001100001",
			2584 => "0010001001000101001100",
			2585 => "0000010110010000101100",
			2586 => "0001011010100000100100",
			2587 => "0010101010011100100000",
			2588 => "0010000101011100010000",
			2589 => "0000000111001100001000",
			2590 => "0001111000111000000100",
			2591 => "0000000010100100101101",
			2592 => "0000000010100100101101",
			2593 => "0001110110101100000100",
			2594 => "0000000010100100101101",
			2595 => "0000000010100100101101",
			2596 => "0000000000001100001000",
			2597 => "0001111000000000000100",
			2598 => "0000000010100100101101",
			2599 => "0000000010100100101101",
			2600 => "0001010001011000000100",
			2601 => "0000000010100100101101",
			2602 => "0000001010100100101101",
			2603 => "0000000010100100101101",
			2604 => "0001011101101100000100",
			2605 => "0000001010100100101101",
			2606 => "0000000010100100101101",
			2607 => "0001111000000000001100",
			2608 => "0011111010100000000100",
			2609 => "0000000010100100101101",
			2610 => "0001011001011000000100",
			2611 => "0000000010100100101101",
			2612 => "0000000010100100101101",
			2613 => "0011001001001000001100",
			2614 => "0000010011110000001000",
			2615 => "0001110001010000000100",
			2616 => "1111111010100100101101",
			2617 => "0000000010100100101101",
			2618 => "0000000010100100101101",
			2619 => "0011111110000000000100",
			2620 => "0000000010100100101101",
			2621 => "0000000010100100101101",
			2622 => "0010011101101000001000",
			2623 => "0010101011000000000100",
			2624 => "0000000010100100101101",
			2625 => "0000000010100100101101",
			2626 => "0001011010001100001000",
			2627 => "0000110000111000000100",
			2628 => "1111111010100100101101",
			2629 => "0000000010100100101101",
			2630 => "0011111110111100000100",
			2631 => "0000000010100100101101",
			2632 => "0010101101101100000100",
			2633 => "0000000010100100101101",
			2634 => "0000000010100100101101",
			2635 => "0001010001011000000100",
			2636 => "1111111010100110011001",
			2637 => "0010001111011000101100",
			2638 => "0000111001111100101000",
			2639 => "0001010001011100010100",
			2640 => "0001111000000100001000",
			2641 => "0000111011111000000100",
			2642 => "0000001010100110011001",
			2643 => "0000001010100110011001",
			2644 => "0000001100000100000100",
			2645 => "1111111010100110011001",
			2646 => "0000000000011100000100",
			2647 => "0000000010100110011001",
			2648 => "1111111010100110011001",
			2649 => "0010010011000000001000",
			2650 => "0000000111000000000100",
			2651 => "0000001010100110011001",
			2652 => "0000001010100110011001",
			2653 => "0000001101001100000100",
			2654 => "0000000010100110011001",
			2655 => "0011001001001000000100",
			2656 => "0000000010100110011001",
			2657 => "0000001010100110011001",
			2658 => "1111111010100110011001",
			2659 => "0000011101000000000100",
			2660 => "0000000010100110011001",
			2661 => "1111111010100110011001",
			2662 => "0001011110111000000100",
			2663 => "1111111010101000001101",
			2664 => "0000100111000100110000",
			2665 => "0010010110000000001000",
			2666 => "0000010111110000000100",
			2667 => "0000000010101000001101",
			2668 => "0000001010101000001101",
			2669 => "0000010110010000010000",
			2670 => "0010101100110100001100",
			2671 => "0011101010011000001000",
			2672 => "0000000000001100000100",
			2673 => "0000000010101000001101",
			2674 => "0000001010101000001101",
			2675 => "0000000010101000001101",
			2676 => "0000001010101000001101",
			2677 => "0000001101001100001100",
			2678 => "0001001100001100001000",
			2679 => "0011101111100100000100",
			2680 => "0000000010101000001101",
			2681 => "1111111010101000001101",
			2682 => "0000000010101000001101",
			2683 => "0010101111100100001000",
			2684 => "0001111000101000000100",
			2685 => "0000000010101000001101",
			2686 => "0000001010101000001101",
			2687 => "1111111010101000001101",
			2688 => "0001011010100000000100",
			2689 => "1111111010101000001101",
			2690 => "0000000010101000001101",
			2691 => "0000001011100001011000",
			2692 => "0000010110010000101000",
			2693 => "0010001001000100100000",
			2694 => "0001100101110000001100",
			2695 => "0011000101010100001000",
			2696 => "0001010001011000000100",
			2697 => "0000000010101011011001",
			2698 => "0000000010101011011001",
			2699 => "0000000010101011011001",
			2700 => "0010010110000000001100",
			2701 => "0001101011110000000100",
			2702 => "0000000010101011011001",
			2703 => "0001111100010000000100",
			2704 => "0000000010101011011001",
			2705 => "0000000010101011011001",
			2706 => "0001001100001100000100",
			2707 => "0000000010101011011001",
			2708 => "0000000010101011011001",
			2709 => "0000010111110000000100",
			2710 => "0000000010101011011001",
			2711 => "0000000010101011011001",
			2712 => "0000100010111100011000",
			2713 => "0011101111100100010100",
			2714 => "0010000101101100001000",
			2715 => "0001011100011100000100",
			2716 => "0000000010101011011001",
			2717 => "0000000010101011011001",
			2718 => "0000101010111100001000",
			2719 => "0010010110000000000100",
			2720 => "0000000010101011011001",
			2721 => "0000000010101011011001",
			2722 => "0000000010101011011001",
			2723 => "0000000010101011011001",
			2724 => "0001000001111100010000",
			2725 => "0010001111001000001000",
			2726 => "0001001100101100000100",
			2727 => "0000000010101011011001",
			2728 => "0000000010101011011001",
			2729 => "0001110001010000000100",
			2730 => "0000000010101011011001",
			2731 => "0000000010101011011001",
			2732 => "0011100110100000000100",
			2733 => "0000000010101011011001",
			2734 => "0000000010101011011001",
			2735 => "0001011111100000001000",
			2736 => "0000111001000000000100",
			2737 => "0000000010101011011001",
			2738 => "0000000010101011011001",
			2739 => "0000111010100000000100",
			2740 => "0000000010101011011001",
			2741 => "0000000010101011011001",
			2742 => "0001010001011000000100",
			2743 => "1111111010101101000101",
			2744 => "0000011101000000101100",
			2745 => "0000111001111100101000",
			2746 => "0010100001101000011100",
			2747 => "0011011010100100001100",
			2748 => "0000001011001000001000",
			2749 => "0010011001000100000100",
			2750 => "0000001010101101000101",
			2751 => "0000001010101101000101",
			2752 => "0000000010101101000101",
			2753 => "0010110101011100001000",
			2754 => "0001010001010100000100",
			2755 => "0000000010101101000101",
			2756 => "1111111010101101000101",
			2757 => "0000000100110100000100",
			2758 => "0000000010101101000101",
			2759 => "0000001010101101000101",
			2760 => "0000000000100100000100",
			2761 => "0000001010101101000101",
			2762 => "0001111001011000000100",
			2763 => "0000001010101101000101",
			2764 => "0000001010101101000101",
			2765 => "1111111010101101000101",
			2766 => "0001111111101000000100",
			2767 => "0000000010101101000101",
			2768 => "1111111010101101000101",
			2769 => "0001010001011000000100",
			2770 => "1111111010101111000001",
			2771 => "0010011001000100001000",
			2772 => "0000000101100000000100",
			2773 => "0000001010101111000001",
			2774 => "0000000010101111000001",
			2775 => "0001011110010100010100",
			2776 => "0011110100100100000100",
			2777 => "1111111010101111000001",
			2778 => "0000000111001100000100",
			2779 => "0000000010101111000001",
			2780 => "0001011010011100001000",
			2781 => "0001010011110100000100",
			2782 => "0000000010101111000001",
			2783 => "0000000010101111000001",
			2784 => "1111111010101111000001",
			2785 => "0011101111100100001100",
			2786 => "0010010011000000001000",
			2787 => "0000010111110000000100",
			2788 => "0000000010101111000001",
			2789 => "0000001010101111000001",
			2790 => "0000000010101111000001",
			2791 => "0000000010111100000100",
			2792 => "1111111010101111000001",
			2793 => "0011101010011000001000",
			2794 => "0000100010111100000100",
			2795 => "0000000010101111000001",
			2796 => "0000001010101111000001",
			2797 => "0000100101000100000100",
			2798 => "1111111010101111000001",
			2799 => "0000000010101111000001",
			2800 => "0001010001011000000100",
			2801 => "1111111010110001000101",
			2802 => "0010011001000100001000",
			2803 => "0000000101100000000100",
			2804 => "0000001010110001000101",
			2805 => "0000000010110001000101",
			2806 => "0001011110010100010100",
			2807 => "0011110100100100001000",
			2808 => "0000010110010000000100",
			2809 => "1111111010110001000101",
			2810 => "1111111010110001000101",
			2811 => "0001010010111000001000",
			2812 => "0000001011001000000100",
			2813 => "0000001010110001000101",
			2814 => "1111111010110001000101",
			2815 => "1111111010110001000101",
			2816 => "0011101001111100010000",
			2817 => "0010001001000100001100",
			2818 => "0011011110011000001000",
			2819 => "0011101101101100000100",
			2820 => "0000001010110001000101",
			2821 => "0000000010110001000101",
			2822 => "0000000010110001000101",
			2823 => "0000000010110001000101",
			2824 => "0000001100111100000100",
			2825 => "1111111010110001000101",
			2826 => "0011101010011000001000",
			2827 => "0010011000000000000100",
			2828 => "0000001010110001000101",
			2829 => "0000000010110001000101",
			2830 => "0000100101000100000100",
			2831 => "0000000010110001000101",
			2832 => "0000000010110001000101",
			2833 => "0010110111011100010100",
			2834 => "0001010001011000000100",
			2835 => "0000000010110011111001",
			2836 => "0001001001000000001100",
			2837 => "0001011110010100001000",
			2838 => "0001011100110100000100",
			2839 => "0000000010110011111001",
			2840 => "0000000010110011111001",
			2841 => "0000000010110011111001",
			2842 => "0000000010110011111001",
			2843 => "0001010001011100100100",
			2844 => "0010011001000100000100",
			2845 => "0000000010110011111001",
			2846 => "0000000000001100001000",
			2847 => "0000011001100100000100",
			2848 => "0000000010110011111001",
			2849 => "0000000010110011111001",
			2850 => "0001101010011000001000",
			2851 => "0000101110000100000100",
			2852 => "0000000010110011111001",
			2853 => "0000000010110011111001",
			2854 => "0000011001100000001000",
			2855 => "0001111101001000000100",
			2856 => "0000000010110011111001",
			2857 => "0000000010110011111001",
			2858 => "0000011101000000000100",
			2859 => "0000000010110011111001",
			2860 => "0000000010110011111001",
			2861 => "0010010011000000000100",
			2862 => "0000000010110011111001",
			2863 => "0000001101001100001000",
			2864 => "0010101100110100000100",
			2865 => "0000000010110011111001",
			2866 => "0000000010110011111001",
			2867 => "0000011000011000001100",
			2868 => "0000110000100000001000",
			2869 => "0011101001110000000100",
			2870 => "0000000010110011111001",
			2871 => "0000000010110011111001",
			2872 => "0000000010110011111001",
			2873 => "0011110011101100000100",
			2874 => "0000000010110011111001",
			2875 => "0010001111011000000100",
			2876 => "0000000010110011111001",
			2877 => "0000000010110011111001",
			2878 => "0001000110101100000100",
			2879 => "1111111010110101011101",
			2880 => "0000101010000000101100",
			2881 => "0010101001111100101000",
			2882 => "0010101100110100011000",
			2883 => "0011010111011100010000",
			2884 => "0001111000000100001000",
			2885 => "0011010110001100000100",
			2886 => "0000001010110101011101",
			2887 => "0000001010110101011101",
			2888 => "0000100100011100000100",
			2889 => "1111111010110101011101",
			2890 => "0000000010110101011101",
			2891 => "0011001001001000000100",
			2892 => "1111111010110101011101",
			2893 => "0000000010110101011101",
			2894 => "0010001001000100000100",
			2895 => "0000001010110101011101",
			2896 => "0000001000100100000100",
			2897 => "0000000010110101011101",
			2898 => "0001010000100000000100",
			2899 => "0000001010110101011101",
			2900 => "0000001010110101011101",
			2901 => "1111111010110101011101",
			2902 => "1111111010110101011101",
			2903 => "0010110111011100100000",
			2904 => "0001011110010100011000",
			2905 => "0001111000000100001000",
			2906 => "0001010001011000000100",
			2907 => "0000000010111000100001",
			2908 => "0000000010111000100001",
			2909 => "0000001110101100000100",
			2910 => "0000000010111000100001",
			2911 => "0000100011100000001000",
			2912 => "0000111100010000000100",
			2913 => "0000000010111000100001",
			2914 => "0000000010111000100001",
			2915 => "0000000010111000100001",
			2916 => "0001010001011100000100",
			2917 => "0000000010111000100001",
			2918 => "0000000010111000100001",
			2919 => "0010001001001100000100",
			2920 => "0000000010111000100001",
			2921 => "0011000101011100010100",
			2922 => "0010011001000100000100",
			2923 => "0000000010111000100001",
			2924 => "0001111101001000001000",
			2925 => "0011111001111100000100",
			2926 => "0000000010111000100001",
			2927 => "0000000010111000100001",
			2928 => "0001100001100000000100",
			2929 => "0000000010111000100001",
			2930 => "0000000010111000100001",
			2931 => "0000110000111100010000",
			2932 => "0001001000100000001100",
			2933 => "0010110101010100001000",
			2934 => "0011110110100000000100",
			2935 => "0000000010111000100001",
			2936 => "0000000010111000100001",
			2937 => "0000000010111000100001",
			2938 => "0000000010111000100001",
			2939 => "0001111000101000001100",
			2940 => "0010100001101000001000",
			2941 => "0001000001011000000100",
			2942 => "0000000010111000100001",
			2943 => "0000000010111000100001",
			2944 => "0000000010111000100001",
			2945 => "0011011001001000001000",
			2946 => "0000111001111100000100",
			2947 => "0000000010111000100001",
			2948 => "0000000010111000100001",
			2949 => "0000000111101100000100",
			2950 => "0000000010111000100001",
			2951 => "0000000010111000100001",
			2952 => "0001010001011000000100",
			2953 => "1111111010111011001111",
			2954 => "0010110111011100010100",
			2955 => "0001011110010100001100",
			2956 => "0001111111011000000100",
			2957 => "0000001010111011001111",
			2958 => "0000001110000100000100",
			2959 => "1111111010111011001111",
			2960 => "0000000010111011001111",
			2961 => "0001111100010000000100",
			2962 => "0000001010111011001111",
			2963 => "0000000010111011001111",
			2964 => "0001011101111100100000",
			2965 => "0000111110111000011000",
			2966 => "0010101001000000001100",
			2967 => "0000010111110000000100",
			2968 => "0000000010111011001111",
			2969 => "0000000010111100000100",
			2970 => "1111111010111011001111",
			2971 => "0000000010111011001111",
			2972 => "0011001001001000000100",
			2973 => "1111111010111011001111",
			2974 => "0001101000110100000100",
			2975 => "0000000010111011001111",
			2976 => "0000000010111011001111",
			2977 => "0001000110011100000100",
			2978 => "0000001010111011001111",
			2979 => "0000000010111011001111",
			2980 => "0010000101101100001100",
			2981 => "0001000010111000001000",
			2982 => "0010010011000000000100",
			2983 => "0000001010111011001111",
			2984 => "0000000010111011001111",
			2985 => "0000000010111011001111",
			2986 => "0001111000101000000100",
			2987 => "1111111010111011001111",
			2988 => "0010101101101100001000",
			2989 => "0001100100010000000100",
			2990 => "0000001010111011001111",
			2991 => "0000000010111011001111",
			2992 => "0000011000011000000100",
			2993 => "0000000010111011001111",
			2994 => "1111111010111011001111",
			2995 => "0011011010100100101100",
			2996 => "0000111011000000011100",
			2997 => "0001111000000100001000",
			2998 => "0001010001011000000100",
			2999 => "0000000010111101110001",
			3000 => "0000000010111101110001",
			3001 => "0000011001100100001000",
			3002 => "0010010110000000000100",
			3003 => "0000000010111101110001",
			3004 => "0000000010111101110001",
			3005 => "0011000101011100000100",
			3006 => "0000000010111101110001",
			3007 => "0010011010000100000100",
			3008 => "0000000010111101110001",
			3009 => "0000000010111101110001",
			3010 => "0011001100101000001000",
			3011 => "0010000101101100000100",
			3012 => "0000000010111101110001",
			3013 => "0000000010111101110001",
			3014 => "0011001001001000000100",
			3015 => "0000000010111101110001",
			3016 => "0000000010111101110001",
			3017 => "0011001100101000001100",
			3018 => "0010110011010000001000",
			3019 => "0001101001011100000100",
			3020 => "0000000010111101110001",
			3021 => "0000000010111101110001",
			3022 => "0000000010111101110001",
			3023 => "0010001001000100010000",
			3024 => "0001001110010100001100",
			3025 => "0010100000111100001000",
			3026 => "0001111100110000000100",
			3027 => "0000000010111101110001",
			3028 => "0000000010111101110001",
			3029 => "0000000010111101110001",
			3030 => "0000000010111101110001",
			3031 => "0001011010001100000100",
			3032 => "0000000010111101110001",
			3033 => "0010101101101100000100",
			3034 => "0000000010111101110001",
			3035 => "0000000010111101110001",
			3036 => "0000010001110000011100",
			3037 => "0001011110010100010100",
			3038 => "0011110100100100000100",
			3039 => "0000000011000000000101",
			3040 => "0000000011100000001000",
			3041 => "0010101101001000000100",
			3042 => "0000000011000000000101",
			3043 => "0000000011000000000101",
			3044 => "0001111001010000000100",
			3045 => "0000000011000000000101",
			3046 => "0000000011000000000101",
			3047 => "0001001100001100000100",
			3048 => "0000000011000000000101",
			3049 => "0000000011000000000101",
			3050 => "0001111000000100001000",
			3051 => "0001010001011000000100",
			3052 => "0000000011000000000101",
			3053 => "0000000011000000000101",
			3054 => "0010100000111000011000",
			3055 => "0011111010110100001000",
			3056 => "0011111101101100000100",
			3057 => "0000000011000000000101",
			3058 => "0000000011000000000101",
			3059 => "0001000011110100001100",
			3060 => "0001111001010000000100",
			3061 => "0000000011000000000101",
			3062 => "0001111011000000000100",
			3063 => "0000000011000000000101",
			3064 => "0000000011000000000101",
			3065 => "0000000011000000000101",
			3066 => "0010101101101100001000",
			3067 => "0010001111011000000100",
			3068 => "0000000011000000000101",
			3069 => "0000000011000000000101",
			3070 => "0000011000011000000100",
			3071 => "0000000011000000000101",
			3072 => "0000000011000000000101",
			3073 => "0010110111011100100000",
			3074 => "0001011110010100011000",
			3075 => "0001111000000100001000",
			3076 => "0001010001011000000100",
			3077 => "0000000011000010110001",
			3078 => "0000000011000010110001",
			3079 => "0000100100100000000100",
			3080 => "0000000011000010110001",
			3081 => "0000100011100000001000",
			3082 => "0000111100010000000100",
			3083 => "0000000011000010110001",
			3084 => "0000000011000010110001",
			3085 => "0000000011000010110001",
			3086 => "0001010001011100000100",
			3087 => "0000000011000010110001",
			3088 => "0000000011000010110001",
			3089 => "0001010001011100011100",
			3090 => "0000000000001100001000",
			3091 => "0010011001000100000100",
			3092 => "0000000011000010110001",
			3093 => "1111111011000010110001",
			3094 => "0011100010011100001000",
			3095 => "0000100111000000000100",
			3096 => "0000000011000010110001",
			3097 => "0000000011000010110001",
			3098 => "0001111101001000000100",
			3099 => "0000000011000010110001",
			3100 => "0010000101101100000100",
			3101 => "0000000011000010110001",
			3102 => "0000000011000010110001",
			3103 => "0010010011000000001000",
			3104 => "0001101110000000000100",
			3105 => "0000000011000010110001",
			3106 => "0000000011000010110001",
			3107 => "0001111000101000001000",
			3108 => "0010100001101000000100",
			3109 => "0000000011000010110001",
			3110 => "0000000011000010110001",
			3111 => "0010101101101100001000",
			3112 => "0000001101110100000100",
			3113 => "0000000011000010110001",
			3114 => "0000000011000010110001",
			3115 => "0000000011000010110001",
			3116 => "0011011010100100111000",
			3117 => "0000111011000000011100",
			3118 => "0001111000000100001000",
			3119 => "0001011110111000000100",
			3120 => "0000000011000101110101",
			3121 => "0000000011000101110101",
			3122 => "0000011001100100001000",
			3123 => "0010010110000000000100",
			3124 => "0000000011000101110101",
			3125 => "0000000011000101110101",
			3126 => "0011000101011100000100",
			3127 => "1111111011000101110101",
			3128 => "0000001011011100000100",
			3129 => "0000000011000101110101",
			3130 => "0000000011000101110101",
			3131 => "0010010011000000010100",
			3132 => "0000011000111100001000",
			3133 => "0000001000001000000100",
			3134 => "0000000011000101110101",
			3135 => "0000000011000101110101",
			3136 => "0010110101010100001000",
			3137 => "0010011101101000000100",
			3138 => "0000001011000101110101",
			3139 => "0000000011000101110101",
			3140 => "0000000011000101110101",
			3141 => "0000001101001100000100",
			3142 => "0000000011000101110101",
			3143 => "0000000011000101110101",
			3144 => "0011001100101000010000",
			3145 => "0010110011010000001000",
			3146 => "0010100100101100000100",
			3147 => "0000000011000101110101",
			3148 => "0000000011000101110101",
			3149 => "0010010011000000000100",
			3150 => "1111111011000101110101",
			3151 => "0000000011000101110101",
			3152 => "0010001001000100010000",
			3153 => "0010100000111100001000",
			3154 => "0000010001110000000100",
			3155 => "0000000011000101110101",
			3156 => "0000000011000101110101",
			3157 => "0001001110010100000100",
			3158 => "0000001011000101110101",
			3159 => "0000000011000101110101",
			3160 => "0001000001101000000100",
			3161 => "0000000011000101110101",
			3162 => "0010101101101100000100",
			3163 => "0000000011000101110101",
			3164 => "0000000011000101110101",
			3165 => "0011011010100100100100",
			3166 => "0000111000100000010100",
			3167 => "0010101001000000010000",
			3168 => "0001000110101100000100",
			3169 => "0000000011001000011001",
			3170 => "0011100010001100000100",
			3171 => "0000001011001000011001",
			3172 => "0001111100010000000100",
			3173 => "0000000011001000011001",
			3174 => "0000000011001000011001",
			3175 => "0000000011001000011001",
			3176 => "0011011110011000001000",
			3177 => "0000011001100100000100",
			3178 => "0000000011001000011001",
			3179 => "0000001011001000011001",
			3180 => "0000101011110100000100",
			3181 => "0000000011001000011001",
			3182 => "0000000011001000011001",
			3183 => "0010110101011100010000",
			3184 => "0010110011010000001000",
			3185 => "0000011000011000000100",
			3186 => "0000000011001000011001",
			3187 => "0000000011001000011001",
			3188 => "0001111001010000000100",
			3189 => "1111111011001000011001",
			3190 => "0000000011001000011001",
			3191 => "0010100000111100000100",
			3192 => "0000000011001000011001",
			3193 => "0000110000111100001000",
			3194 => "0001001011000000000100",
			3195 => "0000000011001000011001",
			3196 => "0000001011001000011001",
			3197 => "0000100010111100000100",
			3198 => "0000000011001000011001",
			3199 => "0011011001001000001000",
			3200 => "0001000001111100000100",
			3201 => "0000000011001000011001",
			3202 => "0000000011001000011001",
			3203 => "0000010001100100000100",
			3204 => "0000000011001000011001",
			3205 => "0000000011001000011001",
			3206 => "0011011010100100110100",
			3207 => "0011101010011000011100",
			3208 => "0001010000111000010000",
			3209 => "0001101011110000001100",
			3210 => "0001110011001000001000",
			3211 => "0001011000100000000100",
			3212 => "0000000011001011010101",
			3213 => "0000000011001011010101",
			3214 => "0000000011001011010101",
			3215 => "0000000011001011010101",
			3216 => "0010110101010100000100",
			3217 => "0000000011001011010101",
			3218 => "0000000010111100000100",
			3219 => "0000000011001011010101",
			3220 => "0000000011001011010101",
			3221 => "0001110110101100001100",
			3222 => "0000111111101000001000",
			3223 => "0000111101001000000100",
			3224 => "0000000011001011010101",
			3225 => "0000000011001011010101",
			3226 => "0000000011001011010101",
			3227 => "0000000101100100000100",
			3228 => "0000000011001011010101",
			3229 => "0010010110000000000100",
			3230 => "0000000011001011010101",
			3231 => "0000000011001011010101",
			3232 => "0000010001110000001000",
			3233 => "0010000101101100000100",
			3234 => "0000000011001011010101",
			3235 => "0000000011001011010101",
			3236 => "0010100000111000010100",
			3237 => "0010110011010000001000",
			3238 => "0001101001011100000100",
			3239 => "0000000011001011010101",
			3240 => "0000000011001011010101",
			3241 => "0001110001010000000100",
			3242 => "0000000011001011010101",
			3243 => "0011110100110000000100",
			3244 => "0000000011001011010101",
			3245 => "0000000011001011010101",
			3246 => "0010101101101100001100",
			3247 => "0011111110111100000100",
			3248 => "0000000011001011010101",
			3249 => "0011110111101000000100",
			3250 => "0000000011001011010101",
			3251 => "0000000011001011010101",
			3252 => "0000000011001011010101",
			3253 => "0000001011100000111100",
			3254 => "0010110111011100011100",
			3255 => "0001011110010100010100",
			3256 => "0001111000000100001000",
			3257 => "0001010001011000000100",
			3258 => "0000000011001101100001",
			3259 => "0000000011001101100001",
			3260 => "0000001110101100000100",
			3261 => "0000000011001101100001",
			3262 => "0000111100010000000100",
			3263 => "0000000011001101100001",
			3264 => "0000000011001101100001",
			3265 => "0001001001000000000100",
			3266 => "0000001011001101100001",
			3267 => "0000000011001101100001",
			3268 => "0000100100011100000100",
			3269 => "0000000011001101100001",
			3270 => "0000001010111100001000",
			3271 => "0011010111011100000100",
			3272 => "0000000011001101100001",
			3273 => "0000000011001101100001",
			3274 => "0011000101011100001000",
			3275 => "0001110110101100000100",
			3276 => "0000000011001101100001",
			3277 => "0000000011001101100001",
			3278 => "0000000100100000000100",
			3279 => "0000000011001101100001",
			3280 => "0000110011110100000100",
			3281 => "0000000011001101100001",
			3282 => "0000000011001101100001",
			3283 => "0001011111100000000100",
			3284 => "0000000011001101100001",
			3285 => "0010100001011100000100",
			3286 => "0000000011001101100001",
			3287 => "0000000011001101100001",
			3288 => "0011011010100100110000",
			3289 => "0000111110111000100100",
			3290 => "0000000111001100100000",
			3291 => "0000001110101100010100",
			3292 => "0001111000000100001000",
			3293 => "0001010001011000000100",
			3294 => "0000000011010000000101",
			3295 => "0000000011010000000101",
			3296 => "0000011001100100000100",
			3297 => "0000000011010000000101",
			3298 => "0011001001001000000100",
			3299 => "0000000011010000000101",
			3300 => "0000000011010000000101",
			3301 => "0011011110011000001000",
			3302 => "0001001001010100000100",
			3303 => "0000000011010000000101",
			3304 => "0000001011010000000101",
			3305 => "0000000011010000000101",
			3306 => "1111111011010000000101",
			3307 => "0001001110111000000100",
			3308 => "0000001011010000000101",
			3309 => "0011001100101000000100",
			3310 => "0000000011010000000101",
			3311 => "0000000011010000000101",
			3312 => "0000100010111100001100",
			3313 => "0000010001110000000100",
			3314 => "0000000011010000000101",
			3315 => "0011000011010000000100",
			3316 => "0000000011010000000101",
			3317 => "1111111011010000000101",
			3318 => "0010110101011100000100",
			3319 => "0000000011010000000101",
			3320 => "0000010001100100001100",
			3321 => "0000110000100000001000",
			3322 => "0001001100101100000100",
			3323 => "0000000011010000000101",
			3324 => "0000001011010000000101",
			3325 => "0000000011010000000101",
			3326 => "0010001010000100000100",
			3327 => "0000000011010000000101",
			3328 => "0000000011010000000101",
			3329 => "0011011010100100110000",
			3330 => "0000111000100000100000",
			3331 => "0010101001000000011100",
			3332 => "0000111011000000011000",
			3333 => "0001111000000100001000",
			3334 => "0001010001011000000100",
			3335 => "0000000011010010110001",
			3336 => "0000000011010010110001",
			3337 => "0001111100110000001000",
			3338 => "0010011010000100000100",
			3339 => "1111111011010010110001",
			3340 => "0000000011010010110001",
			3341 => "0001100010110000000100",
			3342 => "0000000011010010110001",
			3343 => "0000000011010010110001",
			3344 => "0000000011010010110001",
			3345 => "0000000011010010110001",
			3346 => "0011011110011000001000",
			3347 => "0000000000101100000100",
			3348 => "0000001011010010110001",
			3349 => "0000000011010010110001",
			3350 => "0000101011110100000100",
			3351 => "0000000011010010110001",
			3352 => "0000000011010010110001",
			3353 => "0010110101011100010000",
			3354 => "0010110011010000001000",
			3355 => "0000011000011000000100",
			3356 => "0000000011010010110001",
			3357 => "0000000011010010110001",
			3358 => "0001111001010000000100",
			3359 => "1111111011010010110001",
			3360 => "0000000011010010110001",
			3361 => "0010100000111100000100",
			3362 => "1111111011010010110001",
			3363 => "0001011010100000001000",
			3364 => "0000010011110000000100",
			3365 => "0000001011010010110001",
			3366 => "0000000011010010110001",
			3367 => "0010100000111000000100",
			3368 => "0000000011010010110001",
			3369 => "0010101101101100000100",
			3370 => "0000000011010010110001",
			3371 => "0000000011010010110001",
			3372 => "0001010001011000000100",
			3373 => "1111111011010100100101",
			3374 => "0010010110000000001100",
			3375 => "0001010010111000001000",
			3376 => "0001111000000100000100",
			3377 => "0000001011010100100101",
			3378 => "0000000011010100100101",
			3379 => "0000001011010100100101",
			3380 => "0000001100111100010000",
			3381 => "0011100010011100001100",
			3382 => "0000000000001100001000",
			3383 => "0001010001010100000100",
			3384 => "1111111011010100100101",
			3385 => "0000000011010100100101",
			3386 => "0000001011010100100101",
			3387 => "1111111011010100100101",
			3388 => "0011101010011000001000",
			3389 => "0011010101011100000100",
			3390 => "0000001011010100100101",
			3391 => "0000000011010100100101",
			3392 => "0000111011111000001000",
			3393 => "0011111011110100000100",
			3394 => "0000001011010100100101",
			3395 => "0000000011010100100101",
			3396 => "0010011010000100000100",
			3397 => "1111111011010100100101",
			3398 => "0001000010111000000100",
			3399 => "0000000011010100100101",
			3400 => "0000000011010100100101",
			3401 => "0000010110010000111000",
			3402 => "0010001111111100011100",
			3403 => "0001010001101000011000",
			3404 => "0001111100010000010000",
			3405 => "0001111111011000001000",
			3406 => "0010011100101000000100",
			3407 => "0000000011010111011001",
			3408 => "0000000011010111011001",
			3409 => "0001101011110000000100",
			3410 => "0000000011010111011001",
			3411 => "0000000011010111011001",
			3412 => "0000001011001000000100",
			3413 => "0000000011010111011001",
			3414 => "0000000011010111011001",
			3415 => "0000000011010111011001",
			3416 => "0001010010001100010100",
			3417 => "0011111010011000001100",
			3418 => "0000010111110000001000",
			3419 => "0010000101101100000100",
			3420 => "0000000011010111011001",
			3421 => "0000000011010111011001",
			3422 => "0000000011010111011001",
			3423 => "0001011010011100000100",
			3424 => "0000000011010111011001",
			3425 => "0000000011010111011001",
			3426 => "0011001001001000000100",
			3427 => "0000000011010111011001",
			3428 => "0000000011010111011001",
			3429 => "0010010110000000001000",
			3430 => "0001011100011100000100",
			3431 => "0000000011010111011001",
			3432 => "0000000011010111011001",
			3433 => "0001001100001100010100",
			3434 => "0000001101001100000100",
			3435 => "0000000011010111011001",
			3436 => "0000101110110100001100",
			3437 => "0000110001001000001000",
			3438 => "0000000000011100000100",
			3439 => "0000000011010111011001",
			3440 => "0000000011010111011001",
			3441 => "0000000011010111011001",
			3442 => "0000000011010111011001",
			3443 => "0010101101101100000100",
			3444 => "0000000011010111011001",
			3445 => "0000000011010111011001",
			3446 => "0000010110010000110000",
			3447 => "0010001001000100100000",
			3448 => "0001000011000100011000",
			3449 => "0001000110011100010100",
			3450 => "0000000111001100001000",
			3451 => "0001000110101100000100",
			3452 => "0000000011011010011101",
			3453 => "0000000011011010011101",
			3454 => "0001111101001000000100",
			3455 => "0000000011011010011101",
			3456 => "0001111000101000000100",
			3457 => "0000000011011010011101",
			3458 => "0000000011011010011101",
			3459 => "0000000011011010011101",
			3460 => "0011001001001000000100",
			3461 => "0000000011011010011101",
			3462 => "0000000011011010011101",
			3463 => "0001111000000000000100",
			3464 => "0000000011011010011101",
			3465 => "0010101001000000001000",
			3466 => "0010010101111000000100",
			3467 => "0000000011011010011101",
			3468 => "0000000011011010011101",
			3469 => "0000000011011010011101",
			3470 => "0001001100001100100000",
			3471 => "0000100100011000010000",
			3472 => "0010010110000000001100",
			3473 => "0000001110100100000100",
			3474 => "0000000011011010011101",
			3475 => "0001100101110000000100",
			3476 => "0000000011011010011101",
			3477 => "0000000011011010011101",
			3478 => "0000000011011010011101",
			3479 => "0000100111000100001100",
			3480 => "0010100000111100000100",
			3481 => "0000000011011010011101",
			3482 => "0001100010010100000100",
			3483 => "0000000011011010011101",
			3484 => "0000000011011010011101",
			3485 => "0000000011011010011101",
			3486 => "0001000001010100001000",
			3487 => "0001110100101100000100",
			3488 => "0000000011011010011101",
			3489 => "0000000011011010011101",
			3490 => "0011101100100000000100",
			3491 => "0000000011011010011101",
			3492 => "0001111110111000000100",
			3493 => "0000000011011010011101",
			3494 => "0000000011011010011101",
			3495 => "0010001001000101001100",
			3496 => "0011101011110000101100",
			3497 => "0011000101011100011000",
			3498 => "0010011101101000010000",
			3499 => "0001010000111000001100",
			3500 => "0001111000000100001000",
			3501 => "0001011110111000000100",
			3502 => "0000000011011101011001",
			3503 => "0000000011011101011001",
			3504 => "0000000011011101011001",
			3505 => "0000001011011101011001",
			3506 => "0000001011011100000100",
			3507 => "0000000011011101011001",
			3508 => "0000000011011101011001",
			3509 => "0001001001011000001100",
			3510 => "0000110100101100001000",
			3511 => "0000000101000000000100",
			3512 => "0000000011011101011001",
			3513 => "0000000011011101011001",
			3514 => "0000000011011101011001",
			3515 => "0011001100101000000100",
			3516 => "0000000011011101011001",
			3517 => "0000001011011101011001",
			3518 => "0000000100111100001100",
			3519 => "0001000001011000001000",
			3520 => "0000001011110100000100",
			3521 => "0000000011011101011001",
			3522 => "0000000011011101011001",
			3523 => "1111111011011101011001",
			3524 => "0010011010000100010000",
			3525 => "0000011001100100001000",
			3526 => "0001011100101100000100",
			3527 => "0000000011011101011001",
			3528 => "0000000011011101011001",
			3529 => "0000000000011100000100",
			3530 => "0000000011011101011001",
			3531 => "1111111011011101011001",
			3532 => "0000001011011101011001",
			3533 => "0011011110011000001000",
			3534 => "0000011001100000000100",
			3535 => "0000000011011101011001",
			3536 => "0000000011011101011001",
			3537 => "0001011010001100000100",
			3538 => "1111111011011101011001",
			3539 => "0000111010100000000100",
			3540 => "0000000011011101011001",
			3541 => "0000000011011101011001",
			3542 => "0001000110101100000100",
			3543 => "1111111011011111010101",
			3544 => "0010001001000100100000",
			3545 => "0010101100110100011000",
			3546 => "0010101010011100010000",
			3547 => "0000000011100000001100",
			3548 => "0000001100111100001000",
			3549 => "0001101010011000000100",
			3550 => "0000000011011111010101",
			3551 => "1111111011011111010101",
			3552 => "0000001011011111010101",
			3553 => "0000000011011111010101",
			3554 => "0010110101010100000100",
			3555 => "0000000011011111010101",
			3556 => "1111111011011111010101",
			3557 => "0010011000000100000100",
			3558 => "0000001011011111010101",
			3559 => "0000000011011111010101",
			3560 => "0011001100101000000100",
			3561 => "0000000011011111010101",
			3562 => "0001011010001100001100",
			3563 => "0001111011111000000100",
			3564 => "1111111011011111010101",
			3565 => "0000001001110100000100",
			3566 => "0000000011011111010101",
			3567 => "0000000011011111010101",
			3568 => "0010101101101100000100",
			3569 => "0000000011011111010101",
			3570 => "0011011001001000000100",
			3571 => "0000000011011111010101",
			3572 => "0000000011011111010101",
			3573 => "0001011010100001001000",
			3574 => "0011100010011100100000",
			3575 => "0011110000010100011000",
			3576 => "0010011001000100001000",
			3577 => "0001010001011000000100",
			3578 => "0000000011100010010001",
			3579 => "0000000011100010010001",
			3580 => "0001010001010100001100",
			3581 => "0001101010110100001000",
			3582 => "0001111111011000000100",
			3583 => "0000000011100010010001",
			3584 => "0000000011100010010001",
			3585 => "0000000011100010010001",
			3586 => "0000000011100010010001",
			3587 => "0000010111110000000100",
			3588 => "0000000011100010010001",
			3589 => "0000000011100010010001",
			3590 => "0000100111010000001100",
			3591 => "0011010110001100000100",
			3592 => "0000000011100010010001",
			3593 => "0001010010111000000100",
			3594 => "0000000011100010010001",
			3595 => "0000000011100010010001",
			3596 => "0000101011100000010000",
			3597 => "0001010010001100001100",
			3598 => "0000111011000000001000",
			3599 => "0000000111001100000100",
			3600 => "0000000011100010010001",
			3601 => "0000000011100010010001",
			3602 => "0000000011100010010001",
			3603 => "0000000011100010010001",
			3604 => "0011000101101100000100",
			3605 => "0000000011100010010001",
			3606 => "0000110001001000000100",
			3607 => "0000000011100010010001",
			3608 => "0000000011100010010001",
			3609 => "0010000101101100001000",
			3610 => "0001100000110100000100",
			3611 => "0000000011100010010001",
			3612 => "0000000011100010010001",
			3613 => "0001111000101000000100",
			3614 => "0000000011100010010001",
			3615 => "0010101101101100000100",
			3616 => "0000000011100010010001",
			3617 => "0000011000011000000100",
			3618 => "0000000011100010010001",
			3619 => "0000000011100010010001",
			3620 => "0011011010100101000100",
			3621 => "0001011110010100110000",
			3622 => "0011011011101100011100",
			3623 => "0001111111011000001000",
			3624 => "0001011110111000000100",
			3625 => "0000000011100101110101",
			3626 => "0000000011100101110101",
			3627 => "0001111101001000001100",
			3628 => "0001011001000000001000",
			3629 => "0000111000101000000100",
			3630 => "0000000011100101110101",
			3631 => "0000000011100101110101",
			3632 => "1111111011100101110101",
			3633 => "0001100110111000000100",
			3634 => "0000000011100101110101",
			3635 => "0000000011100101110101",
			3636 => "0000100100011100001100",
			3637 => "0001110011001000001000",
			3638 => "0000000010000000000100",
			3639 => "0000000011100101110101",
			3640 => "0000000011100101110101",
			3641 => "0000000011100101110101",
			3642 => "0001001001010100000100",
			3643 => "0000000011100101110101",
			3644 => "0000001011100101110101",
			3645 => "0001000001011000001000",
			3646 => "0000000000000100000100",
			3647 => "0000000011100101110101",
			3648 => "0000001011100101110101",
			3649 => "0011100000100000001000",
			3650 => "0010110101010100000100",
			3651 => "0000000011100101110101",
			3652 => "0000000011100101110101",
			3653 => "0000000011100101110101",
			3654 => "0011001100101000010000",
			3655 => "0010110011010000001000",
			3656 => "0010100100101100000100",
			3657 => "0000000011100101110101",
			3658 => "0000000011100101110101",
			3659 => "0010010011000000000100",
			3660 => "1111111011100101110101",
			3661 => "0000000011100101110101",
			3662 => "0010001001000100010000",
			3663 => "0010100000111100001000",
			3664 => "0000010001110000000100",
			3665 => "0000000011100101110101",
			3666 => "0000000011100101110101",
			3667 => "0001001110010100000100",
			3668 => "0000001011100101110101",
			3669 => "0000000011100101110101",
			3670 => "0001000001101000000100",
			3671 => "0000000011100101110101",
			3672 => "0011111110111100000100",
			3673 => "0000000011100101110101",
			3674 => "0010101101101100000100",
			3675 => "0000000011100101110101",
			3676 => "0000000011100101110101",
			3677 => "0011011110011000101100",
			3678 => "0001011110010100100100",
			3679 => "0001111000000100010000",
			3680 => "0001011110111000001100",
			3681 => "0000010001110000000100",
			3682 => "0000000011101001000001",
			3683 => "0000010111110000000100",
			3684 => "0000000011101001000001",
			3685 => "0000000011101001000001",
			3686 => "0000000011101001000001",
			3687 => "0001101010001100000100",
			3688 => "0000000011101001000001",
			3689 => "0010110011010000001000",
			3690 => "0011011011101100000100",
			3691 => "0000000011101001000001",
			3692 => "0000000011101001000001",
			3693 => "0001100011101100000100",
			3694 => "0000000011101001000001",
			3695 => "0000000011101001000001",
			3696 => "0010010011000000000100",
			3697 => "0000000011101001000001",
			3698 => "0000000011101001000001",
			3699 => "0000000000100100011000",
			3700 => "0001111100000000001000",
			3701 => "0000000100111000000100",
			3702 => "0000000011101001000001",
			3703 => "0000000011101001000001",
			3704 => "0000111011111000001000",
			3705 => "0010011101101000000100",
			3706 => "0000000011101001000001",
			3707 => "0000000011101001000001",
			3708 => "0010100000111000000100",
			3709 => "0000000011101001000001",
			3710 => "0000000011101001000001",
			3711 => "0011101110000000001000",
			3712 => "0011110001001100000100",
			3713 => "0000000011101001000001",
			3714 => "0000000011101001000001",
			3715 => "0011001001001000001100",
			3716 => "0010101000100000001000",
			3717 => "0010101011000000000100",
			3718 => "0000000011101001000001",
			3719 => "0000000011101001000001",
			3720 => "0000000011101001000001",
			3721 => "0000100111000100001100",
			3722 => "0000111001111100001000",
			3723 => "0010101001000000000100",
			3724 => "0000000011101001000001",
			3725 => "0000000011101001000001",
			3726 => "0000000011101001000001",
			3727 => "0000000011101001000001",
			3728 => "0001010001011000000100",
			3729 => "1111111011101010101101",
			3730 => "0010001111011000101100",
			3731 => "0010101100110100011100",
			3732 => "0001111000000100000100",
			3733 => "0000001011101010101101",
			3734 => "0000000001111000001000",
			3735 => "0011000101011100000100",
			3736 => "0000000011101010101101",
			3737 => "1111111011101010101101",
			3738 => "0011100010011100001000",
			3739 => "0011110000010100000100",
			3740 => "0000000011101010101101",
			3741 => "0000001011101010101101",
			3742 => "0000100111010000000100",
			3743 => "1111111011101010101101",
			3744 => "0000000011101010101101",
			3745 => "0000111001111100001100",
			3746 => "0010001001000100000100",
			3747 => "0000001011101010101101",
			3748 => "0010011000000100000100",
			3749 => "0000000011101010101101",
			3750 => "0000001011101010101101",
			3751 => "1111111011101010101101",
			3752 => "0000011101000000000100",
			3753 => "0000000011101010101101",
			3754 => "1111111011101010101101",
			3755 => "0011011010100100111000",
			3756 => "0000101000100100101100",
			3757 => "0000001110101100011000",
			3758 => "0011100101110000010000",
			3759 => "0001010000111000001100",
			3760 => "0001111000000100001000",
			3761 => "0001010001011000000100",
			3762 => "0000000011101110000001",
			3763 => "0000000011101110000001",
			3764 => "0000000011101110000001",
			3765 => "0000000011101110000001",
			3766 => "0011010110001100000100",
			3767 => "0000000011101110000001",
			3768 => "0000000011101110000001",
			3769 => "0011100000010100001100",
			3770 => "0000011000111100000100",
			3771 => "0000000011101110000001",
			3772 => "0001001001010100000100",
			3773 => "0000000011101110000001",
			3774 => "0000000011101110000001",
			3775 => "0000010000011000000100",
			3776 => "0000000011101110000001",
			3777 => "0000000011101110000001",
			3778 => "0001110110101100000100",
			3779 => "0000000011101110000001",
			3780 => "0000111011111000000100",
			3781 => "0000000011101110000001",
			3782 => "0000000011101110000001",
			3783 => "0011001100101000001100",
			3784 => "0010110011010000001000",
			3785 => "0001101001011100000100",
			3786 => "0000000011101110000001",
			3787 => "0000000011101110000001",
			3788 => "0000000011101110000001",
			3789 => "0000011000011000011000",
			3790 => "0010100000111100001000",
			3791 => "0010001111111100000100",
			3792 => "0000000011101110000001",
			3793 => "0000000011101110000001",
			3794 => "0001011101101100000100",
			3795 => "0000000011101110000001",
			3796 => "0000110001101000000100",
			3797 => "0000000011101110000001",
			3798 => "0001011110010000000100",
			3799 => "0000000011101110000001",
			3800 => "0000000011101110000001",
			3801 => "0011010101010100001000",
			3802 => "0000000101100100000100",
			3803 => "0000000011101110000001",
			3804 => "0000000011101110000001",
			3805 => "0000001011110100000100",
			3806 => "0000000011101110000001",
			3807 => "0000000011101110000001",
			3808 => "0001010001011000000100",
			3809 => "1111111011110000001101",
			3810 => "0011011010100100100000",
			3811 => "0000111011000000001100",
			3812 => "0001111000000100000100",
			3813 => "0000001011110000001101",
			3814 => "0000001011011100000100",
			3815 => "1111111011110000001101",
			3816 => "0000000011110000001101",
			3817 => "0000010110010000001100",
			3818 => "0011111010011000000100",
			3819 => "0000000011110000001101",
			3820 => "0010110011010000000100",
			3821 => "0000000011110000001101",
			3822 => "0000001011110000001101",
			3823 => "0000000010111100000100",
			3824 => "0000000011110000001101",
			3825 => "0000001011110000001101",
			3826 => "0001000001011000001100",
			3827 => "0001111001010000000100",
			3828 => "1111111011110000001101",
			3829 => "0000000011111000000100",
			3830 => "0000000011110000001101",
			3831 => "1111111011110000001101",
			3832 => "0000111110111000000100",
			3833 => "0000001011110000001101",
			3834 => "0000100010111100000100",
			3835 => "1111111011110000001101",
			3836 => "0011101110000000001000",
			3837 => "0010001111001000000100",
			3838 => "0000001011110000001101",
			3839 => "0000000011110000001101",
			3840 => "0011110011101100000100",
			3841 => "1111111011110000001101",
			3842 => "0000000011110000001101",
			3843 => "0001001111101000001100",
			3844 => "0001010001011000000100",
			3845 => "1111111011110010000001",
			3846 => "0000001011001000000100",
			3847 => "0000001011110010000001",
			3848 => "1111111011110010000001",
			3849 => "0011011001001000101100",
			3850 => "0001000000100000101000",
			3851 => "0010101100001100011000",
			3852 => "0011011010100100001100",
			3853 => "0001111000000100000100",
			3854 => "0000011011110010000001",
			3855 => "0000000001111000000100",
			3856 => "0000000011110010000001",
			3857 => "0000010011110010000001",
			3858 => "0000000101100100001000",
			3859 => "0011101111100100000100",
			3860 => "0000000011110010000001",
			3861 => "1111111011110010000001",
			3862 => "0000001011110010000001",
			3863 => "0001110110011100001100",
			3864 => "0001111100110000000100",
			3865 => "0000011011110010000001",
			3866 => "0000001101001100000100",
			3867 => "0000010011110010000001",
			3868 => "0000010011110010000001",
			3869 => "0000011011110010000001",
			3870 => "1111111011110010000001",
			3871 => "1111111011110010000001",
			3872 => "0011101101000101000000",
			3873 => "0011110001101100111000",
			3874 => "0010010110000000010000",
			3875 => "0001011100110100001100",
			3876 => "0001001111101000001000",
			3877 => "0000111101001000000100",
			3878 => "0000000011110100110101",
			3879 => "0000000011110100110101",
			3880 => "0000000011110100110101",
			3881 => "0000001011110100110101",
			3882 => "0010100000111100001100",
			3883 => "0000001110000100000100",
			3884 => "1111111011110100110101",
			3885 => "0011011010100100000100",
			3886 => "0000000011110100110101",
			3887 => "0000000011110100110101",
			3888 => "0011101111111000010000",
			3889 => "0000000100100000001000",
			3890 => "0001010001010100000100",
			3891 => "1111111011110100110101",
			3892 => "0000000011110100110101",
			3893 => "0011000101011100000100",
			3894 => "0000000011110100110101",
			3895 => "0000000011110100110101",
			3896 => "0000000100111100000100",
			3897 => "1111111011110100110101",
			3898 => "0001110100101100000100",
			3899 => "0000000011110100110101",
			3900 => "0000000011110100110101",
			3901 => "0001001001010100000100",
			3902 => "0000000011110100110101",
			3903 => "0000001011110100110101",
			3904 => "0011001001001000001100",
			3905 => "0010000101011100001000",
			3906 => "0010001001001100000100",
			3907 => "0000000011110100110101",
			3908 => "0000000011110100110101",
			3909 => "1111111011110100110101",
			3910 => "0000101110110100001100",
			3911 => "0000110000100000001000",
			3912 => "0001000110011100000100",
			3913 => "0000000011110100110101",
			3914 => "0000000011110100110101",
			3915 => "0000000011110100110101",
			3916 => "0000000011110100110101",
			3917 => "0001011010011100001100",
			3918 => "0001010001011000000100",
			3919 => "1111111011110111000001",
			3920 => "0010110111011100000100",
			3921 => "0000001011110111000001",
			3922 => "1111111011110111000001",
			3923 => "0011011001001000110000",
			3924 => "0000111001111100101100",
			3925 => "0001010001011100011000",
			3926 => "0010110111011100001100",
			3927 => "0001011110010100001000",
			3928 => "0001111000000100000100",
			3929 => "0000010011110111000001",
			3930 => "0000000011110111000001",
			3931 => "0000010011110111000001",
			3932 => "0011111010011000000100",
			3933 => "1111111011110111000001",
			3934 => "0011100010011100000100",
			3935 => "0000001011110111000001",
			3936 => "0000000011110111000001",
			3937 => "0000001101001100001000",
			3938 => "0010010011000000000100",
			3939 => "0000010011110111000001",
			3940 => "0000000011110111000001",
			3941 => "0000111010011100000100",
			3942 => "0000010011110111000001",
			3943 => "0000111100110100000100",
			3944 => "0000001011110111000001",
			3945 => "0000001011110111000001",
			3946 => "1111111011110111000001",
			3947 => "0000010001100100001000",
			3948 => "0001011010110000000100",
			3949 => "0000001011110111000001",
			3950 => "1111111011110111000001",
			3951 => "1111111011110111000001",
			3952 => "0011101010011000110000",
			3953 => "0000000010111100100000",
			3954 => "0001101010011000011100",
			3955 => "0010001001000100010100",
			3956 => "0000000100100000010000",
			3957 => "0010010110000000001000",
			3958 => "0000000011101100000100",
			3959 => "0000000011111010010101",
			3960 => "0000001011111010010101",
			3961 => "0001010001010100000100",
			3962 => "1111111011111010010101",
			3963 => "0000000011111010010101",
			3964 => "0000000011111010010101",
			3965 => "0010011001000100000100",
			3966 => "0000000011111010010101",
			3967 => "1111111011111010010101",
			3968 => "1111111011111010010101",
			3969 => "0001111000000000000100",
			3970 => "0000000011111010010101",
			3971 => "0011010101011100001000",
			3972 => "0000001100111100000100",
			3973 => "0000000011111010010101",
			3974 => "0000001011111010010101",
			3975 => "0000000011111010010101",
			3976 => "0010100001101000101100",
			3977 => "0010001111111100011100",
			3978 => "0000000011100000001000",
			3979 => "0000000100111100000100",
			3980 => "0000000011111010010101",
			3981 => "0000001011111010010101",
			3982 => "0000011001100100001000",
			3983 => "0001110110101100000100",
			3984 => "0000000011111010010101",
			3985 => "0000000011111010010101",
			3986 => "0011011011101100000100",
			3987 => "1111111011111010010101",
			3988 => "0001111101001000000100",
			3989 => "0000000011111010010101",
			3990 => "0000000011111010010101",
			3991 => "0011001001001000001000",
			3992 => "0010110101011100000100",
			3993 => "1111111011111010010101",
			3994 => "0000000011111010010101",
			3995 => "0000001010101000000100",
			3996 => "0000000011111010010101",
			3997 => "0000000011111010010101",
			3998 => "0010101101101100001000",
			3999 => "0000001110110100000100",
			4000 => "0000000011111010010101",
			4001 => "0000000011111010010101",
			4002 => "0011011001001000000100",
			4003 => "0000000011111010010101",
			4004 => "0000000011111010010101",
			4005 => "0001011110010100110100",
			4006 => "0011011011101100010100",
			4007 => "0001111000000100001000",
			4008 => "0001011110111000000100",
			4009 => "0000000011111101100001",
			4010 => "0000000011111101100001",
			4011 => "0001011001000000001000",
			4012 => "0001010110011100000100",
			4013 => "0000000011111101100001",
			4014 => "0000000011111101100001",
			4015 => "0000000011111101100001",
			4016 => "0010100000111100011000",
			4017 => "0001111100000000001100",
			4018 => "0010010110000000001000",
			4019 => "0000001101100100000100",
			4020 => "0000000011111101100001",
			4021 => "0000000011111101100001",
			4022 => "0000000011111101100001",
			4023 => "0000010000011000001000",
			4024 => "0000001001111000000100",
			4025 => "0000000011111101100001",
			4026 => "0000000011111101100001",
			4027 => "0000000011111101100001",
			4028 => "0000000000011100000100",
			4029 => "0000000011111101100001",
			4030 => "0000000011111101100001",
			4031 => "0011011110011000001100",
			4032 => "0001001100011100001000",
			4033 => "0000010001110000000100",
			4034 => "0000000011111101100001",
			4035 => "0000000011111101100001",
			4036 => "0000000011111101100001",
			4037 => "0000111000100000000100",
			4038 => "0000000011111101100001",
			4039 => "0000100111000000001000",
			4040 => "0000110011110100000100",
			4041 => "0000000011111101100001",
			4042 => "0000000011111101100001",
			4043 => "0011100010010100010000",
			4044 => "0010001111001000001000",
			4045 => "0001001110010100000100",
			4046 => "0000000011111101100001",
			4047 => "0000000011111101100001",
			4048 => "0000011000011000000100",
			4049 => "0000000011111101100001",
			4050 => "0000000011111101100001",
			4051 => "0011101111000100000100",
			4052 => "0000000011111101100001",
			4053 => "0000011101000000000100",
			4054 => "0000000011111101100001",
			4055 => "0000000011111101100001",
			4056 => "0010110111011100100000",
			4057 => "0001011110010100011000",
			4058 => "0001111000000100001000",
			4059 => "0001010001011000000100",
			4060 => "0000000100000000000101",
			4061 => "0000000100000000000101",
			4062 => "0000001110101100000100",
			4063 => "0000000100000000000101",
			4064 => "0000100011100000001000",
			4065 => "0000111100010000000100",
			4066 => "0000000100000000000101",
			4067 => "0000000100000000000101",
			4068 => "0000000100000000000101",
			4069 => "0001011111100000000100",
			4070 => "0000000100000000000101",
			4071 => "0000000100000000000101",
			4072 => "0000100100011100000100",
			4073 => "0000000100000000000101",
			4074 => "0000001010111100001000",
			4075 => "0011010011010000000100",
			4076 => "0000000100000000000101",
			4077 => "0000000100000000000101",
			4078 => "0011000101011100001100",
			4079 => "0001110110101100000100",
			4080 => "0000000100000000000101",
			4081 => "0010110101010100000100",
			4082 => "0000000100000000000101",
			4083 => "0000000100000000000101",
			4084 => "0000010110010000001100",
			4085 => "0011100000010100001000",
			4086 => "0001001001011000000100",
			4087 => "0000000100000000000101",
			4088 => "0000000100000000000101",
			4089 => "0000000100000000000101",
			4090 => "0000100010111100001000",
			4091 => "0000010011110000000100",
			4092 => "0000000100000000000101",
			4093 => "0000000100000000000101",
			4094 => "0011011001001000000100",
			4095 => "0000000100000000000101",
			4096 => "0000000100000000000101",
			4097 => "0001010001011000000100",
			4098 => "1111111100000001111001",
			4099 => "0000100111000100110000",
			4100 => "0010110111011100010000",
			4101 => "0001011110010100001000",
			4102 => "0001111111011000000100",
			4103 => "0000001100000001111001",
			4104 => "0000000100000001111001",
			4105 => "0001010001011100000100",
			4106 => "0000001100000001111001",
			4107 => "0000000100000001111001",
			4108 => "0000100111100000000100",
			4109 => "1111111100000001111001",
			4110 => "0011001100101000001100",
			4111 => "0011011010100100001000",
			4112 => "0011101001111100000100",
			4113 => "0000001100000001111001",
			4114 => "0000000100000001111001",
			4115 => "1111111100000001111001",
			4116 => "0011010011010000001000",
			4117 => "0010110101011100000100",
			4118 => "0000000100000001111001",
			4119 => "0000001100000001111001",
			4120 => "0001111000101000000100",
			4121 => "0000000100000001111001",
			4122 => "0000000100000001111001",
			4123 => "0001011010100000000100",
			4124 => "1111111100000001111001",
			4125 => "0000000100000001111001",
			4126 => "0010001111001001001100",
			4127 => "0010101011000000010100",
			4128 => "0001111000000100001000",
			4129 => "0001010000111100000100",
			4130 => "0000000100000100100101",
			4131 => "0000000100000100100101",
			4132 => "0010011010000100000100",
			4133 => "0000000100000100100101",
			4134 => "0010010011000000000100",
			4135 => "0000000100000100100101",
			4136 => "0000000100000100100101",
			4137 => "0001000010111000101100",
			4138 => "0001011110010100010100",
			4139 => "0011011011101100001000",
			4140 => "0001111100110000000100",
			4141 => "0000000100000100100101",
			4142 => "0000000100000100100101",
			4143 => "0000000000001100000100",
			4144 => "0000000100000100100101",
			4145 => "0001101111110100000100",
			4146 => "0000000100000100100101",
			4147 => "0000000100000100100101",
			4148 => "0001111100010000001000",
			4149 => "0000010111110000000100",
			4150 => "0000000100000100100101",
			4151 => "0000001100000100100101",
			4152 => "0000001101001100001000",
			4153 => "0000010110010000000100",
			4154 => "0000000100000100100101",
			4155 => "0000000100000100100101",
			4156 => "0001001100001100000100",
			4157 => "0000001100000100100101",
			4158 => "0000000100000100100101",
			4159 => "0001110001010000000100",
			4160 => "0000000100000100100101",
			4161 => "0010111001000100000100",
			4162 => "0000000100000100100101",
			4163 => "0000000100000100100101",
			4164 => "0001001110010100000100",
			4165 => "0000000100000100100101",
			4166 => "0001010011101100000100",
			4167 => "0000000100000100100101",
			4168 => "0000000100000100100101",
			4169 => "0010110111011100010000",
			4170 => "0001010001011000000100",
			4171 => "0000000100000111001001",
			4172 => "0001011110010100001000",
			4173 => "0001011100110100000100",
			4174 => "0000000100000111001001",
			4175 => "0000000100000111001001",
			4176 => "0000000100000111001001",
			4177 => "0001010001011100100100",
			4178 => "0010011001000100000100",
			4179 => "0000000100000111001001",
			4180 => "0000000000001100001000",
			4181 => "0000011001100100000100",
			4182 => "0000000100000111001001",
			4183 => "0000000100000111001001",
			4184 => "0001101010011000001000",
			4185 => "0000101110000100000100",
			4186 => "0000000100000111001001",
			4187 => "0000000100000111001001",
			4188 => "0000011001100000001000",
			4189 => "0001111101001000000100",
			4190 => "0000000100000111001001",
			4191 => "0000000100000111001001",
			4192 => "0000011101000000000100",
			4193 => "0000000100000111001001",
			4194 => "0000000100000111001001",
			4195 => "0010010011000000000100",
			4196 => "0000000100000111001001",
			4197 => "0000000100111100001000",
			4198 => "0010100000111000000100",
			4199 => "0000000100000111001001",
			4200 => "0000000100000111001001",
			4201 => "0010101101101100001000",
			4202 => "0000001101110100000100",
			4203 => "0000000100000111001001",
			4204 => "0000000100000111001001",
			4205 => "0000011000011000000100",
			4206 => "0000000100000111001001",
			4207 => "0000100101100100000100",
			4208 => "0000000100000111001001",
			4209 => "0000000100000111001001",
			4210 => "0001000110101100000100",
			4211 => "1111111100001001010101",
			4212 => "0010110111011100010100",
			4213 => "0000001011001000010000",
			4214 => "0011110100100100001000",
			4215 => "0001111000000100000100",
			4216 => "0000001100001001010101",
			4217 => "0000000100001001010101",
			4218 => "0010101010011100000100",
			4219 => "0000001100001001010101",
			4220 => "0000000100001001010101",
			4221 => "1111111100001001010101",
			4222 => "0001010001011100011000",
			4223 => "0000000000001100000100",
			4224 => "1111111100001001010101",
			4225 => "0010101010011100010000",
			4226 => "0000000000011100001000",
			4227 => "0000110001001000000100",
			4228 => "0000001100001001010101",
			4229 => "0000000100001001010101",
			4230 => "0000110001001000000100",
			4231 => "1111111100001001010101",
			4232 => "0000001100001001010101",
			4233 => "1111111100001001010101",
			4234 => "0011011110011000001000",
			4235 => "0011101111000000000100",
			4236 => "0000001100001001010101",
			4237 => "0000000100001001010101",
			4238 => "0010110101011100000100",
			4239 => "0000000100001001010101",
			4240 => "0000111110111000000100",
			4241 => "0000001100001001010101",
			4242 => "0000100010111100000100",
			4243 => "1111111100001001010101",
			4244 => "0000000100001001010101",
			4245 => "0001010001011000000100",
			4246 => "1111111100001011011001",
			4247 => "0010001001000100100100",
			4248 => "0000100111101100100000",
			4249 => "0000000100111100010100",
			4250 => "0011100000100000010000",
			4251 => "0000001110101100001000",
			4252 => "0011101111100100000100",
			4253 => "0000000100001011011001",
			4254 => "1111111100001011011001",
			4255 => "0001111100010000000100",
			4256 => "0000000100001011011001",
			4257 => "0000001100001011011001",
			4258 => "1111111100001011011001",
			4259 => "0000010001110000000100",
			4260 => "0000001100001011011001",
			4261 => "0000000000011100000100",
			4262 => "0000001100001011011001",
			4263 => "0000000100001011011001",
			4264 => "0000000100001011011001",
			4265 => "0011111110111100001000",
			4266 => "0011111111000000000100",
			4267 => "0000000100001011011001",
			4268 => "1111111100001011011001",
			4269 => "0011100101001000000100",
			4270 => "0000001100001011011001",
			4271 => "0011000101101100000100",
			4272 => "1111111100001011011001",
			4273 => "0011010101101100001000",
			4274 => "0000110000100000000100",
			4275 => "0000001100001011011001",
			4276 => "0000000100001011011001",
			4277 => "1111111100001011011001",
			4278 => "0011011010100100110000",
			4279 => "0000111110111000101000",
			4280 => "0000000111001100100100",
			4281 => "0010110101010100010100",
			4282 => "0000001110101100001100",
			4283 => "0011100111010100001000",
			4284 => "0001010000111000000100",
			4285 => "0000000100001110000101",
			4286 => "0000000100001110000101",
			4287 => "0000000100001110000101",
			4288 => "0001001001010100000100",
			4289 => "0000000100001110000101",
			4290 => "0000000100001110000101",
			4291 => "0011001001001000001000",
			4292 => "0000111011111000000100",
			4293 => "0000000100001110000101",
			4294 => "0000000100001110000101",
			4295 => "0001111100010000000100",
			4296 => "0000000100001110000101",
			4297 => "0000000100001110000101",
			4298 => "0000000100001110000101",
			4299 => "0000011000111100000100",
			4300 => "0000000100001110000101",
			4301 => "0000000100001110000101",
			4302 => "0001101111111000001000",
			4303 => "0010110011010000000100",
			4304 => "0000000100001110000101",
			4305 => "1111111100001110000101",
			4306 => "0010110101011100000100",
			4307 => "0000000100001110000101",
			4308 => "0000010110010000000100",
			4309 => "0000001100001110000101",
			4310 => "0010100000111000001100",
			4311 => "0011001001001000000100",
			4312 => "0000000100001110000101",
			4313 => "0001011110001100000100",
			4314 => "0000000100001110000101",
			4315 => "0000000100001110000101",
			4316 => "0010101101101100001000",
			4317 => "0001001100001100000100",
			4318 => "0000000100001110000101",
			4319 => "0000000100001110000101",
			4320 => "0000000100001110000101",
			4321 => "0000001011100001010100",
			4322 => "0000001101001100101100",
			4323 => "0001100010010100100100",
			4324 => "0010011001000100001000",
			4325 => "0001010001011000000100",
			4326 => "0000000100010001001001",
			4327 => "0000001100010001001001",
			4328 => "0000001110101100010000",
			4329 => "0010100000111100001000",
			4330 => "0001111000000100000100",
			4331 => "0000000100010001001001",
			4332 => "1111111100010001001001",
			4333 => "0001111100010000000100",
			4334 => "0000000100010001001001",
			4335 => "0000000100010001001001",
			4336 => "0001101010001100000100",
			4337 => "0000000100010001001001",
			4338 => "0001101010011000000100",
			4339 => "0000001100010001001001",
			4340 => "0000000100010001001001",
			4341 => "0011011011101100000100",
			4342 => "0000000100010001001001",
			4343 => "1111111100010001001001",
			4344 => "0000000000011100010100",
			4345 => "0011010101010100001000",
			4346 => "0001001001010100000100",
			4347 => "0000000100010001001001",
			4348 => "0000001100010001001001",
			4349 => "0000011000011000000100",
			4350 => "0000000100010001001001",
			4351 => "0001110100101100000100",
			4352 => "0000000100010001001001",
			4353 => "0000000100010001001001",
			4354 => "0011100000010100000100",
			4355 => "1111111100010001001001",
			4356 => "0011011010100100000100",
			4357 => "0000001100010001001001",
			4358 => "0000101011011000000100",
			4359 => "0000000100010001001001",
			4360 => "0000111010011000000100",
			4361 => "0000000100010001001001",
			4362 => "0000000100010001001001",
			4363 => "0000111001000000000100",
			4364 => "1111111100010001001001",
			4365 => "0000011101000000001000",
			4366 => "0011110100101000000100",
			4367 => "0000000100010001001001",
			4368 => "0000001100010001001001",
			4369 => "0000000100010001001001",
			4370 => "0011011010100100111000",
			4371 => "0000111000100000101000",
			4372 => "0001111000000100001000",
			4373 => "0001011110111000000100",
			4374 => "0000000100010100101101",
			4375 => "0000000100010100101101",
			4376 => "0001111000111000001100",
			4377 => "0010011001000100001000",
			4378 => "0011010110001100000100",
			4379 => "0000000100010100101101",
			4380 => "0000000100010100101101",
			4381 => "0000000100010100101101",
			4382 => "0000000111001100010000",
			4383 => "0000010110010000001000",
			4384 => "0010110101011100000100",
			4385 => "0000000100010100101101",
			4386 => "0000000100010100101101",
			4387 => "0000001011011100000100",
			4388 => "0000000100010100101101",
			4389 => "0000000100010100101101",
			4390 => "0000000100010100101101",
			4391 => "0001000001011000000100",
			4392 => "0000000100010100101101",
			4393 => "0010001111111100001000",
			4394 => "0010011010000100000100",
			4395 => "0000000100010100101101",
			4396 => "0000000100010100101101",
			4397 => "0000000100010100101101",
			4398 => "0010110101011100010100",
			4399 => "0010110011010000001000",
			4400 => "0001101001011100000100",
			4401 => "0000000100010100101101",
			4402 => "0000000100010100101101",
			4403 => "0001001000101000001000",
			4404 => "0010101011000000000100",
			4405 => "0000000100010100101101",
			4406 => "0000000100010100101101",
			4407 => "0000000100010100101101",
			4408 => "0010100000111100000100",
			4409 => "0000000100010100101101",
			4410 => "0001000000111000010100",
			4411 => "0000010011110000001000",
			4412 => "0001011010100000000100",
			4413 => "0000000100010100101101",
			4414 => "0000000100010100101101",
			4415 => "0001101111000100000100",
			4416 => "0000000100010100101101",
			4417 => "0001101000110100000100",
			4418 => "0000000100010100101101",
			4419 => "0000000100010100101101",
			4420 => "0011111110111100000100",
			4421 => "0000000100010100101101",
			4422 => "0011100000010100000100",
			4423 => "0000000100010100101101",
			4424 => "0011101100100000000100",
			4425 => "0000000100010100101101",
			4426 => "0000000100010100101101",
			4427 => "0011101010011000110000",
			4428 => "0000100010111100100100",
			4429 => "0011101001111100100000",
			4430 => "0010001001000100010100",
			4431 => "0011001100101000001100",
			4432 => "0000111000100000001000",
			4433 => "0010011001000100000100",
			4434 => "0000001100011000000001",
			4435 => "0000000100011000000001",
			4436 => "0000000100011000000001",
			4437 => "0000000111101000000100",
			4438 => "0000000100011000000001",
			4439 => "0000001100011000000001",
			4440 => "0010010110000000001000",
			4441 => "0011000111011100000100",
			4442 => "0000000100011000000001",
			4443 => "0000000100011000000001",
			4444 => "1111111100011000000001",
			4445 => "1111111100011000000001",
			4446 => "0011111001110000000100",
			4447 => "0000000100011000000001",
			4448 => "0000100100111100000100",
			4449 => "0000001100011000000001",
			4450 => "0000000100011000000001",
			4451 => "0000011000111100001100",
			4452 => "0000000110001000000100",
			4453 => "1111111100011000000001",
			4454 => "0000001100100100000100",
			4455 => "0000000100011000000001",
			4456 => "0000000100011000000001",
			4457 => "0000111110111000011000",
			4458 => "0010001111111100010100",
			4459 => "0000000011100000001000",
			4460 => "0001011000000100000100",
			4461 => "0000000100011000000001",
			4462 => "0000001100011000000001",
			4463 => "0001110110101100000100",
			4464 => "1111111100011000000001",
			4465 => "0001111101001000000100",
			4466 => "0000000100011000000001",
			4467 => "0000000100011000000001",
			4468 => "1111111100011000000001",
			4469 => "0001101111000100000100",
			4470 => "0000000100011000000001",
			4471 => "0000011000011000000100",
			4472 => "0000001100011000000001",
			4473 => "0011111100011000001000",
			4474 => "0001101110111100000100",
			4475 => "0000000100011000000001",
			4476 => "0000000100011000000001",
			4477 => "0000011101000000000100",
			4478 => "0000000100011000000001",
			4479 => "0000000100011000000001",
			4480 => "0001010001011000000100",
			4481 => "1111111100011001111101",
			4482 => "0010001111011000110100",
			4483 => "0001111000000100001000",
			4484 => "0000111011111000000100",
			4485 => "0000001100011001111101",
			4486 => "0000001100011001111101",
			4487 => "0001011110010100010000",
			4488 => "0011011011101100000100",
			4489 => "1111111100011001111101",
			4490 => "0010101001011000000100",
			4491 => "1111111100011001111101",
			4492 => "0011011010100100000100",
			4493 => "0000001100011001111101",
			4494 => "0000000100011001111101",
			4495 => "0011011110011000001100",
			4496 => "0010011101101000000100",
			4497 => "0000001100011001111101",
			4498 => "0010001111111100000100",
			4499 => "0000001100011001111101",
			4500 => "0000000100011001111101",
			4501 => "0010110101011100001000",
			4502 => "0010001111111100000100",
			4503 => "0000000100011001111101",
			4504 => "1111111100011001111101",
			4505 => "0000111001111100000100",
			4506 => "0000001100011001111101",
			4507 => "1111111100011001111101",
			4508 => "0000011101000000000100",
			4509 => "0000000100011001111101",
			4510 => "1111111100011001111101",
			4511 => "0001010001011000000100",
			4512 => "1111111100011100001001",
			4513 => "0000100111101100110100",
			4514 => "0010011001000100000100",
			4515 => "0000001100011100001001",
			4516 => "0000001110101100010100",
			4517 => "0001000000111100001100",
			4518 => "0011100100000000001000",
			4519 => "0001100101110000000100",
			4520 => "1111111100011100001001",
			4521 => "0000000100011100001001",
			4522 => "1111111100011100001001",
			4523 => "0010010011000000000100",
			4524 => "0000001100011100001001",
			4525 => "1111111100011100001001",
			4526 => "0001000001011000001100",
			4527 => "0011011010100100001000",
			4528 => "0001111100010000000100",
			4529 => "0000001100011100001001",
			4530 => "0000001100011100001001",
			4531 => "0000000100011100001001",
			4532 => "0001101101000100001000",
			4533 => "0010011100000000000100",
			4534 => "0000001100011100001001",
			4535 => "1111111100011100001001",
			4536 => "0000000100111100000100",
			4537 => "1111111100011100001001",
			4538 => "0000000100011100001001",
			4539 => "0001011111100000001000",
			4540 => "0000111001000000000100",
			4541 => "1111111100011100001001",
			4542 => "0000000100011100001001",
			4543 => "0011011001001000000100",
			4544 => "0000001100011100001001",
			4545 => "1111111100011100001001",
			4546 => "0000001011100001101000",
			4547 => "0000010110010000111000",
			4548 => "0000010111110000110000",
			4549 => "0010001111111100011100",
			4550 => "0001111000000000001100",
			4551 => "0001111000000100001000",
			4552 => "0001011001011000000100",
			4553 => "0000000100011111110111",
			4554 => "0000000100011111110111",
			4555 => "0000000100011111110111",
			4556 => "0011010110001100001000",
			4557 => "0011111110100100000100",
			4558 => "0000000100011111110111",
			4559 => "0000000100011111110111",
			4560 => "0001101101101100000100",
			4561 => "0000000100011111110111",
			4562 => "0000000100011111110111",
			4563 => "0011011110011000001100",
			4564 => "0000000001111000001000",
			4565 => "0011000101010100000100",
			4566 => "0000000100011111110111",
			4567 => "0000000100011111110111",
			4568 => "0000000100011111110111",
			4569 => "0011001001001000000100",
			4570 => "0000000100011111110111",
			4571 => "0000000100011111110111",
			4572 => "0010100000111100000100",
			4573 => "0000000100011111110111",
			4574 => "0000000100011111110111",
			4575 => "0000100010111100011000",
			4576 => "0011101111100100010100",
			4577 => "0010000101101100001000",
			4578 => "0001011100011100000100",
			4579 => "0000000100011111110111",
			4580 => "0000000100011111110111",
			4581 => "0000101010111100001000",
			4582 => "0010010110000000000100",
			4583 => "0000000100011111110111",
			4584 => "0000000100011111110111",
			4585 => "0000000100011111110111",
			4586 => "0000000100011111110111",
			4587 => "0001000001111100010000",
			4588 => "0010001111001000001000",
			4589 => "0001001100101100000100",
			4590 => "0000000100011111110111",
			4591 => "0000000100011111110111",
			4592 => "0001110001010000000100",
			4593 => "0000000100011111110111",
			4594 => "0000000100011111110111",
			4595 => "0011100110100000000100",
			4596 => "0000000100011111110111",
			4597 => "0000000100011111110111",
			4598 => "0001011111100000001000",
			4599 => "0000111001000000000100",
			4600 => "0000000100011111110111",
			4601 => "0000000100011111110111",
			4602 => "0000111010100000000100",
			4603 => "0000000100011111110111",
			4604 => "0000000100011111110111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1473, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2995, initial_addr_3'length));
	end generate gen_rom_8;

	gen_rom_9: if SELECT_ROM = 9 generate
		bank <= (
			0 => "0011111101101100010100",
			1 => "0000101101000100001100",
			2 => "0000111100101000001000",
			3 => "0000100000111000000100",
			4 => "0000000000000001001101",
			5 => "0000000000000001001101",
			6 => "0000000000000001001101",
			7 => "0000111001010100000100",
			8 => "0000000000000001001101",
			9 => "0000000000000001001101",
			10 => "0000100111010000001000",
			11 => "0000100010111100000100",
			12 => "0000000000000001001101",
			13 => "0000000000000001001101",
			14 => "0000101011001000001000",
			15 => "0001001111100000000100",
			16 => "0000000000000001001101",
			17 => "0000000000000001001101",
			18 => "0000000000000001001101",
			19 => "0001010011000000011000",
			20 => "0011110101110000010000",
			21 => "0000100000111000000100",
			22 => "0000000000000010101001",
			23 => "0010001010000100001000",
			24 => "0000111101101000000100",
			25 => "0000000000000010101001",
			26 => "0000000000000010101001",
			27 => "0000000000000010101001",
			28 => "0000000101100000000100",
			29 => "0000000000000010101001",
			30 => "0000000000000010101001",
			31 => "0000001010101100001100",
			32 => "0001000101010100000100",
			33 => "0000000000000010101001",
			34 => "0011000110000000000100",
			35 => "0000000000000010101001",
			36 => "0000000000000010101001",
			37 => "0011111001110000000100",
			38 => "0000000000000010101001",
			39 => "0001111000000000000100",
			40 => "0000000000000010101001",
			41 => "0000000000000010101001",
			42 => "0011111111100000011100",
			43 => "0000101101000100010100",
			44 => "0000111100101000010000",
			45 => "0000010001110000001000",
			46 => "0000100001001000000100",
			47 => "0000000000000100000101",
			48 => "0000000000000100000101",
			49 => "0001000001110000000100",
			50 => "0000000000000100000101",
			51 => "0000000000000100000101",
			52 => "0000000000000100000101",
			53 => "0000111111011000000100",
			54 => "0000000000000100000101",
			55 => "0000000000000100000101",
			56 => "0000100010111100001000",
			57 => "0010100101101100000100",
			58 => "0000000000000100000101",
			59 => "0000000000000100000101",
			60 => "0011110001001100001000",
			61 => "0001000000100000000100",
			62 => "0000000000000100000101",
			63 => "0000000000000100000101",
			64 => "0000000000000100000101",
			65 => "0011110100100100100100",
			66 => "0000101101000100010000",
			67 => "0000111100101000001100",
			68 => "0010011010100100000100",
			69 => "0000000000000101101001",
			70 => "0000000001101000000100",
			71 => "0000000000000101101001",
			72 => "0000000000000101101001",
			73 => "0000000000000101101001",
			74 => "0011111111100000001000",
			75 => "0000111111011000000100",
			76 => "0000000000000101101001",
			77 => "0000000000000101101001",
			78 => "0000101000110100001000",
			79 => "0010110101010100000100",
			80 => "0000000000000101101001",
			81 => "0000000000000101101001",
			82 => "0000000000000101101001",
			83 => "0010111111011000001000",
			84 => "0010001010100100000100",
			85 => "0000000000000101101001",
			86 => "0000000000000101101001",
			87 => "0010010001010000000100",
			88 => "0000000000000101101001",
			89 => "0000000000000101101001",
			90 => "0001100000010100100000",
			91 => "0000100000111000000100",
			92 => "0000000000000110110101",
			93 => "0001011100011100001000",
			94 => "0011011010000100000100",
			95 => "0000000000000110110101",
			96 => "0000000000000110110101",
			97 => "0001000110011100001000",
			98 => "0000111000100000000100",
			99 => "0000000000000110110101",
			100 => "0000000000000110110101",
			101 => "0010100000111100000100",
			102 => "0000000000000110110101",
			103 => "0001001101111100000100",
			104 => "0000000000000110110101",
			105 => "0000000000000110110101",
			106 => "0011011000000100000100",
			107 => "0000000000000110110101",
			108 => "0000000000000110110101",
			109 => "0011110100100100101100",
			110 => "0000100010110000011000",
			111 => "0001101110111000010000",
			112 => "0000101101101100001000",
			113 => "0010110110110100000100",
			114 => "0000000000001000110001",
			115 => "0000000000001000110001",
			116 => "0000110011000000000100",
			117 => "0000000000001000110001",
			118 => "0000000000001000110001",
			119 => "0000011101000000000100",
			120 => "0000000000001000110001",
			121 => "0000000000001000110001",
			122 => "0001010001101000001100",
			123 => "0010111001001000000100",
			124 => "0000000000001000110001",
			125 => "0000111001010100000100",
			126 => "0000000000001000110001",
			127 => "0000000000001000110001",
			128 => "0010010011000000000100",
			129 => "0000000000001000110001",
			130 => "0000000000001000110001",
			131 => "0011001010000100001000",
			132 => "0000011000111100000100",
			133 => "0000000000001000110001",
			134 => "0000000000001000110001",
			135 => "0001111000100000001000",
			136 => "0000101011011000000100",
			137 => "0000000000001000110001",
			138 => "0000000000001000110001",
			139 => "0000000000001000110001",
			140 => "0001100000010100101100",
			141 => "0000101110010000011100",
			142 => "0011111010011100001100",
			143 => "0000100000111000000100",
			144 => "0000000000001010010101",
			145 => "0000110011000000000100",
			146 => "0000000000001010010101",
			147 => "0000000000001010010101",
			148 => "0010110101010100001000",
			149 => "0000011101000000000100",
			150 => "0000000000001010010101",
			151 => "0000000000001010010101",
			152 => "0010101000101000000100",
			153 => "0000000000001010010101",
			154 => "0000000000001010010101",
			155 => "0001010001101000000100",
			156 => "0000000000001010010101",
			157 => "0001011010100000000100",
			158 => "0000000000001010010101",
			159 => "0001001101111100000100",
			160 => "0000000000001010010101",
			161 => "0000000000001010010101",
			162 => "0011011000000100000100",
			163 => "0000000000001010010101",
			164 => "0000000000001010010101",
			165 => "0011110001001100101000",
			166 => "0000100001100000011100",
			167 => "0011110001010100010100",
			168 => "0000111111011000001100",
			169 => "0000100000111000000100",
			170 => "0000000000001011101001",
			171 => "0000111101101000000100",
			172 => "0000000000001011101001",
			173 => "0000000000001011101001",
			174 => "0001110011001000000100",
			175 => "0000000000001011101001",
			176 => "0000000000001011101001",
			177 => "0001011001001000000100",
			178 => "0000000000001011101001",
			179 => "0000000000001011101001",
			180 => "0001010001101000000100",
			181 => "0000000000001011101001",
			182 => "0000100100111100000100",
			183 => "0000000000001011101001",
			184 => "0000000000001011101001",
			185 => "0000000000001011101001",
			186 => "0011110100100100101000",
			187 => "0000000111001000010100",
			188 => "0011110011110100010000",
			189 => "0001101000111000000100",
			190 => "0000000000001101010101",
			191 => "0010011001001000000100",
			192 => "0000000000001101010101",
			193 => "0000110111011100000100",
			194 => "0000000000001101010101",
			195 => "0000000000001101010101",
			196 => "0000000000001101010101",
			197 => "0011010110000000010000",
			198 => "0011110000100000001000",
			199 => "0001010001101000000100",
			200 => "0000000000001101010101",
			201 => "0000000000001101010101",
			202 => "0011111010011000000100",
			203 => "0000000000001101010101",
			204 => "0000000000001101010101",
			205 => "0000000000001101010101",
			206 => "0011011101000000000100",
			207 => "0000000000001101010101",
			208 => "0011001010000100000100",
			209 => "0000000000001101010101",
			210 => "0001111000100000000100",
			211 => "0000000000001101010101",
			212 => "0000000000001101010101",
			213 => "0011110001001100101100",
			214 => "0000101110010000011100",
			215 => "0011111010011100001100",
			216 => "0000110011000000001000",
			217 => "0000100000111000000100",
			218 => "0000000000001110110001",
			219 => "0000000000001110110001",
			220 => "0000000000001110110001",
			221 => "0010110101010100001000",
			222 => "0000011101000000000100",
			223 => "0000000000001110110001",
			224 => "0000000000001110110001",
			225 => "0010101000101000000100",
			226 => "0000000000001110110001",
			227 => "0000000000001110110001",
			228 => "0001010001101000000100",
			229 => "0000000000001110110001",
			230 => "0010100000111000000100",
			231 => "0000000000001110110001",
			232 => "0001001101111100000100",
			233 => "0000000000001110110001",
			234 => "0000000000001110110001",
			235 => "0000000000001110110001",
			236 => "0010001010100100001000",
			237 => "0011011101000000000100",
			238 => "0000000000010000100101",
			239 => "0000000000010000100101",
			240 => "0010110101010100011100",
			241 => "0011110011110100001100",
			242 => "0011110110011100001000",
			243 => "0001011001100000000100",
			244 => "0000000000010000100101",
			245 => "0000000000010000100101",
			246 => "0000000000010000100101",
			247 => "0000011000111100000100",
			248 => "0000000000010000100101",
			249 => "0001000001011000000100",
			250 => "0000000000010000100101",
			251 => "0001001110111000000100",
			252 => "0000000000010000100101",
			253 => "0000000000010000100101",
			254 => "0000101101100100001000",
			255 => "0001111101101000000100",
			256 => "0000000000010000100101",
			257 => "0000000000010000100101",
			258 => "0011111001110000001000",
			259 => "0010101010011000000100",
			260 => "0000000000010000100101",
			261 => "0000000000010000100101",
			262 => "0011011000000100000100",
			263 => "0000000000010000100101",
			264 => "0000000000010000100101",
			265 => "0001100101001000110000",
			266 => "0000101101000100010000",
			267 => "0001101001011000001100",
			268 => "0000100000111000000100",
			269 => "0000000000010010010001",
			270 => "0010100110000000000100",
			271 => "0000000000010010010001",
			272 => "0000000000010010010001",
			273 => "0000000000010010010001",
			274 => "0011111111100000001000",
			275 => "0001011001010100000100",
			276 => "0000000000010010010001",
			277 => "0000000000010010010001",
			278 => "0000101000110100001100",
			279 => "0011011110011000000100",
			280 => "0000000000010010010001",
			281 => "0001001101101000000100",
			282 => "0000000000010010010001",
			283 => "0000000000010010010001",
			284 => "0001010001101000000100",
			285 => "0000000000010010010001",
			286 => "0000000010101000000100",
			287 => "0000000000010010010001",
			288 => "0000000000010010010001",
			289 => "0011011000000100000100",
			290 => "0000000000010010010001",
			291 => "0000000000010010010001",
			292 => "0001100101001000110100",
			293 => "0000101101100000100000",
			294 => "0011111010011100011000",
			295 => "0011000101010100001100",
			296 => "0000100000111000000100",
			297 => "0000000000010100000101",
			298 => "0011011011101100000100",
			299 => "0000000000010100000101",
			300 => "0000000000010100000101",
			301 => "0001000001100100001000",
			302 => "0001111111011000000100",
			303 => "0000000000010100000101",
			304 => "0000000000010100000101",
			305 => "0000000000010100000101",
			306 => "0000011101000000000100",
			307 => "0000000000010100000101",
			308 => "0000000000010100000101",
			309 => "0001011100110100001000",
			310 => "0011110100100100000100",
			311 => "0000000000010100000101",
			312 => "0000000000010100000101",
			313 => "0010111001000100001000",
			314 => "0011111001111100000100",
			315 => "0000000000010100000101",
			316 => "0000000000010100000101",
			317 => "0000000000010100000101",
			318 => "0011011000000100000100",
			319 => "0000000000010100000101",
			320 => "0000000000010100000101",
			321 => "0010001010100100001000",
			322 => "0011011101000000000100",
			323 => "0000000000010110000001",
			324 => "0000000000010110000001",
			325 => "0010110101010100011100",
			326 => "0011110011110100001100",
			327 => "0011110110011100001000",
			328 => "0001011001100000000100",
			329 => "0000000000010110000001",
			330 => "0000000000010110000001",
			331 => "0000000000010110000001",
			332 => "0000011000111100000100",
			333 => "0000000000010110000001",
			334 => "0001000001011000000100",
			335 => "0000000000010110000001",
			336 => "0001001110111000000100",
			337 => "0000000000010110000001",
			338 => "0000000000010110000001",
			339 => "0000101101100100001100",
			340 => "0001111111011000001000",
			341 => "0001111101101000000100",
			342 => "0000000000010110000001",
			343 => "0000000000010110000001",
			344 => "0000000000010110000001",
			345 => "0011111001110000001000",
			346 => "0010101010011000000100",
			347 => "0000000000010110000001",
			348 => "0000000000010110000001",
			349 => "0011011000000100000100",
			350 => "0000000000010110000001",
			351 => "0000000000010110000001",
			352 => "0011110110100000110000",
			353 => "0000101000110100100100",
			354 => "0001011001010100011100",
			355 => "0000101101000100010000",
			356 => "0001101001011000001100",
			357 => "0000100000111000000100",
			358 => "0000000000010111110101",
			359 => "0010100101101100000100",
			360 => "0000000000010111110101",
			361 => "0000000000010111110101",
			362 => "0000000000010111110101",
			363 => "0011110111010100001000",
			364 => "0000010110010000000100",
			365 => "0000001000010111110101",
			366 => "0000000000010111110101",
			367 => "0000000000010111110101",
			368 => "0001000101111000000100",
			369 => "0000000000010111110101",
			370 => "1111111000010111110101",
			371 => "0011110100100100000100",
			372 => "0000001000010111110101",
			373 => "0000100100110100000100",
			374 => "0000000000010111110101",
			375 => "0000000000010111110101",
			376 => "0011011000000100000100",
			377 => "1111111000010111110101",
			378 => "0001001001010000000100",
			379 => "0000000000010111110101",
			380 => "0000000000010111110101",
			381 => "0011110001001100110000",
			382 => "0000000000110100010100",
			383 => "0011110011110100010000",
			384 => "0000100000111000000100",
			385 => "0000000000011001011001",
			386 => "0010011001001000000100",
			387 => "0000000000011001011001",
			388 => "0001110101111000000100",
			389 => "0000000000011001011001",
			390 => "0000000000011001011001",
			391 => "0000000000011001011001",
			392 => "0001100001111100001000",
			393 => "0001011001010000000100",
			394 => "0000001000011001011001",
			395 => "0000000000011001011001",
			396 => "0000100101001100001000",
			397 => "0001000101010100000100",
			398 => "0000000000011001011001",
			399 => "0000000000011001011001",
			400 => "0001010001101000000100",
			401 => "0000000000011001011001",
			402 => "0000100100111100000100",
			403 => "0000000000011001011001",
			404 => "0000000000011001011001",
			405 => "0000000000011001011001",
			406 => "0001100000010100110100",
			407 => "0000101101100000100000",
			408 => "0001101100011100011000",
			409 => "0011000101010100001100",
			410 => "0000100000111000000100",
			411 => "0000000000011011001101",
			412 => "0011011011101100000100",
			413 => "0000000000011011001101",
			414 => "0000000000011011001101",
			415 => "0001010110001100001000",
			416 => "0001110101111000000100",
			417 => "0000000000011011001101",
			418 => "0000000000011011001101",
			419 => "0000000000011011001101",
			420 => "0000011101000000000100",
			421 => "0000000000011011001101",
			422 => "0000000000011011001101",
			423 => "0001011100110100000100",
			424 => "0000000000011011001101",
			425 => "0000100101111100001100",
			426 => "0001111000000000001000",
			427 => "0001111100000000000100",
			428 => "0000000000011011001101",
			429 => "0000000000011011001101",
			430 => "0000000000011011001101",
			431 => "0000000000011011001101",
			432 => "0011011000000100000100",
			433 => "0000000000011011001101",
			434 => "0000000000011011001101",
			435 => "0011110001001100110100",
			436 => "0000101101000100001100",
			437 => "0010000011010000000100",
			438 => "0000000000011100111001",
			439 => "0001000001110000000100",
			440 => "0000000000011100111001",
			441 => "1111111000011100111001",
			442 => "0001010100101100010100",
			443 => "0001101101111100001100",
			444 => "0000100010110000001000",
			445 => "0001111101101000000100",
			446 => "0000001000011100111001",
			447 => "0000000000011100111001",
			448 => "0000001000011100111001",
			449 => "0000001101010000000100",
			450 => "0000000000011100111001",
			451 => "0000001000011100111001",
			452 => "0000100000100100001100",
			453 => "0011111101101100001000",
			454 => "0000001101100100000100",
			455 => "0000000000011100111001",
			456 => "0000000000011100111001",
			457 => "1111111000011100111001",
			458 => "0001000000100000000100",
			459 => "0000001000011100111001",
			460 => "0000000000011100111001",
			461 => "1111111000011100111001",
			462 => "0011110001001100110100",
			463 => "0000101100100000010100",
			464 => "0011110011110100010000",
			465 => "0000100000111000000100",
			466 => "0000000000011110100101",
			467 => "0010011001001000000100",
			468 => "0000000000011110100101",
			469 => "0001110101111000000100",
			470 => "0000000000011110100101",
			471 => "0000000000011110100101",
			472 => "0000000000011110100101",
			473 => "0001100001111100001100",
			474 => "0001011001010000001000",
			475 => "0010001010000100000100",
			476 => "0000001000011110100101",
			477 => "0000000000011110100101",
			478 => "0000000000011110100101",
			479 => "0000101000110100001000",
			480 => "0001000101010100000100",
			481 => "0000000000011110100101",
			482 => "0000000000011110100101",
			483 => "0011110100100100000100",
			484 => "0000000000011110100101",
			485 => "0000101011011000000100",
			486 => "0000000000011110100101",
			487 => "0000000000011110100101",
			488 => "0000000000011110100101",
			489 => "0001100000010100101100",
			490 => "0000100010111100101000",
			491 => "0001101111100000011100",
			492 => "0000101101000100010000",
			493 => "0001101001011000001100",
			494 => "0000100000111000000100",
			495 => "0000000000100000001001",
			496 => "0010100110000000000100",
			497 => "0000000000100000001001",
			498 => "0000000000100000001001",
			499 => "0000000000100000001001",
			500 => "0001000101111000001000",
			501 => "0010001010000100000100",
			502 => "0000000000100000001001",
			503 => "0000000000100000001001",
			504 => "0000000000100000001001",
			505 => "0000101000010100000100",
			506 => "0000000000100000001001",
			507 => "0011011011101100000100",
			508 => "0000000000100000001001",
			509 => "0000000000100000001001",
			510 => "0000000000100000001001",
			511 => "0011011000000100000100",
			512 => "0000000000100000001001",
			513 => "0000000000100000001001",
			514 => "0011110001001100100100",
			515 => "0000101111100000000100",
			516 => "1111111000100001010101",
			517 => "0001111000100000011100",
			518 => "0000001000001000010100",
			519 => "0001101111100100001100",
			520 => "0010101111111100000100",
			521 => "0000001000100001010101",
			522 => "0000000111001000000100",
			523 => "1111111000100001010101",
			524 => "0000001000100001010101",
			525 => "0000100010111100000100",
			526 => "1111111000100001010101",
			527 => "0000000000100001010101",
			528 => "0001000000100000000100",
			529 => "0000001000100001010101",
			530 => "1111111000100001010101",
			531 => "1111111000100001010101",
			532 => "1111111000100001010101",
			533 => "0011110001001100110000",
			534 => "0000100111010000101000",
			535 => "0011110100000000011100",
			536 => "0000000000110100010000",
			537 => "0011110001011000001100",
			538 => "0000100000111000000100",
			539 => "0000000000100010111001",
			540 => "0010011001001000000100",
			541 => "0000000000100010111001",
			542 => "0000000000100010111001",
			543 => "0000000000100010111001",
			544 => "0000111001010100001000",
			545 => "0010001010000100000100",
			546 => "0000000000100010111001",
			547 => "0000000000100010111001",
			548 => "0000000000100010111001",
			549 => "0000101000010100000100",
			550 => "0000000000100010111001",
			551 => "0000000010111100000100",
			552 => "0000000000100010111001",
			553 => "0000000000100010111001",
			554 => "0001000000100000000100",
			555 => "0000000000100010111001",
			556 => "0000000000100010111001",
			557 => "0000000000100010111001",
			558 => "0000011001100100011000",
			559 => "0001001110011000001100",
			560 => "0010101010100100001000",
			561 => "0011110110000000000100",
			562 => "0000000000100101001101",
			563 => "0000000000100101001101",
			564 => "0000000000100101001101",
			565 => "0011011011101100001000",
			566 => "0001111000000000000100",
			567 => "0000000000100101001101",
			568 => "0000000000100101001101",
			569 => "0000000000100101001101",
			570 => "0010001010100100000100",
			571 => "0000000000100101001101",
			572 => "0010110101010100010100",
			573 => "0001011111011100001000",
			574 => "0011110011001000000100",
			575 => "0000000000100101001101",
			576 => "0000000000100101001101",
			577 => "0001000001011000000100",
			578 => "0000000000100101001101",
			579 => "0001001100011100000100",
			580 => "0000000000100101001101",
			581 => "0000000000100101001101",
			582 => "0010101000101000001100",
			583 => "0000000010000000000100",
			584 => "0000000000100101001101",
			585 => "0001110001010000000100",
			586 => "0000000000100101001101",
			587 => "0000000000100101001101",
			588 => "0000101011110100000100",
			589 => "0000000000100101001101",
			590 => "0001101001110000001000",
			591 => "0000111001111100000100",
			592 => "0000000000100101001101",
			593 => "0000000000100101001101",
			594 => "0000000000100101001101",
			595 => "0011110001001100111000",
			596 => "0000100001100000100100",
			597 => "0011110001010100011000",
			598 => "0000100000111000000100",
			599 => "1111111000100111000001",
			600 => "0000110101111000001100",
			601 => "0000111100101000000100",
			602 => "0000001000100111000001",
			603 => "0010101010000100000100",
			604 => "0000000000100111000001",
			605 => "0000001000100111000001",
			606 => "0001110011001000000100",
			607 => "1111111000100111000001",
			608 => "0000000000100111000001",
			609 => "0000000111001000000100",
			610 => "1111111000100111000001",
			611 => "0011110111010100000100",
			612 => "0000000000100111000001",
			613 => "1111111000100111000001",
			614 => "0011110000100000000100",
			615 => "0000001000100111000001",
			616 => "0000000101000100001000",
			617 => "0000100111000000000100",
			618 => "1111111000100111000001",
			619 => "0000000000100111000001",
			620 => "0001000000100000000100",
			621 => "0000001000100111000001",
			622 => "0000000000100111000001",
			623 => "1111111000100111000001",
			624 => "0001100000010100110100",
			625 => "0000101111100000001000",
			626 => "0011011101000000000100",
			627 => "0000000000101000111101",
			628 => "1111111000101000111101",
			629 => "0001010001101000100100",
			630 => "0000100101001100011000",
			631 => "0001101001101100010000",
			632 => "0001011001010100001000",
			633 => "0000101101000100000100",
			634 => "0000001000101000111101",
			635 => "0000001000101000111101",
			636 => "0001001000000100000100",
			637 => "0000000000101000111101",
			638 => "1111111000101000111101",
			639 => "0001011101101000000100",
			640 => "0000000000101000111101",
			641 => "1111111000101000111101",
			642 => "0011011011101100000100",
			643 => "0000001000101000111101",
			644 => "0010011010000100000100",
			645 => "0000001000101000111101",
			646 => "0000001000101000111101",
			647 => "0000011101000000000100",
			648 => "1111111000101000111101",
			649 => "0000001000101000111101",
			650 => "0011110001001100001000",
			651 => "0001011111111000000100",
			652 => "0000001000101000111101",
			653 => "1111111000101000111101",
			654 => "1111111000101000111101",
			655 => "0011110001001100110100",
			656 => "0000101101000100001100",
			657 => "0010000011010000000100",
			658 => "0000000000101010101001",
			659 => "0001000001110000000100",
			660 => "0000000000101010101001",
			661 => "1111111000101010101001",
			662 => "0001010001101000100000",
			663 => "0000001010101100011000",
			664 => "0001100001111100001100",
			665 => "0001011001010100001000",
			666 => "0000010110010000000100",
			667 => "0000001000101010101001",
			668 => "0000001000101010101001",
			669 => "0000000000101010101001",
			670 => "0000100100101000000100",
			671 => "1111111000101010101001",
			672 => "0011101001101100000100",
			673 => "0000001000101010101001",
			674 => "1111111000101010101001",
			675 => "0011110100100100000100",
			676 => "0000001000101010101001",
			677 => "0000000000101010101001",
			678 => "0000000111001100000100",
			679 => "1111111000101010101001",
			680 => "0000001000101010101001",
			681 => "1111111000101010101001",
			682 => "0001100101001000111100",
			683 => "0000101111100000001000",
			684 => "0011011101000000000100",
			685 => "0000000000101100110101",
			686 => "1111111000101100110101",
			687 => "0001010011110100100100",
			688 => "0000101101100100010000",
			689 => "0001011001001000001000",
			690 => "0001101110111000000100",
			691 => "0000001000101100110101",
			692 => "0000001000101100110101",
			693 => "0000010001110000000100",
			694 => "0000001000101100110101",
			695 => "1111111000101100110101",
			696 => "0001101101101100001100",
			697 => "0011111111100100001000",
			698 => "0000011001100000000100",
			699 => "0000010000101100110101",
			700 => "0000001000101100110101",
			701 => "0000001000101100110101",
			702 => "0000000111000000000100",
			703 => "1111111000101100110101",
			704 => "0000010000101100110101",
			705 => "0000001000001000001100",
			706 => "0000010000011000001000",
			707 => "0001101010110100000100",
			708 => "0000000000101100110101",
			709 => "1111111000101100110101",
			710 => "1111111000101100110101",
			711 => "0000010000101100110101",
			712 => "0011011000000100000100",
			713 => "1111111000101100110101",
			714 => "0001100010010000000100",
			715 => "0000000000101100110101",
			716 => "1111111000101100110101",
			717 => "0011110001001100101000",
			718 => "0000101111100000000100",
			719 => "1111111000101110001001",
			720 => "0010101010100100000100",
			721 => "0000001000101110001001",
			722 => "0000100111010000010100",
			723 => "0011110000100000010000",
			724 => "0000101000101100001000",
			725 => "0011111111100000000100",
			726 => "0000000000101110001001",
			727 => "1111111000101110001001",
			728 => "0011111101101100000100",
			729 => "0000001000101110001001",
			730 => "0000000000101110001001",
			731 => "1111111000101110001001",
			732 => "0000111001111100001000",
			733 => "0000000101000100000100",
			734 => "0000000000101110001001",
			735 => "0000001000101110001001",
			736 => "1111111000101110001001",
			737 => "1111111000101110001001",
			738 => "0011110001001100111100",
			739 => "0000101101000100010000",
			740 => "0010110110001100001000",
			741 => "0011000110110100000100",
			742 => "0000000000110000000101",
			743 => "0000001000110000000101",
			744 => "0001001001100100000100",
			745 => "0000000000110000000101",
			746 => "1111111000110000000101",
			747 => "0000011001100100001000",
			748 => "0011110000100000000100",
			749 => "0000001000110000000101",
			750 => "0000000000110000000101",
			751 => "0010110101010100010000",
			752 => "0001011001001000000100",
			753 => "0000000000110000000101",
			754 => "0000100001100000000100",
			755 => "1111111000110000000101",
			756 => "0001101011110000000100",
			757 => "0000000000110000000101",
			758 => "0000000000110000000101",
			759 => "0010101000101000001000",
			760 => "0011100001011100000100",
			761 => "0000001000110000000101",
			762 => "0000000000110000000101",
			763 => "0000101011110100000100",
			764 => "1111111000110000000101",
			765 => "0001000000100000000100",
			766 => "0000001000110000000101",
			767 => "0000000000110000000101",
			768 => "1111111000110000000101",
			769 => "0011110110100000111100",
			770 => "0000100000111000000100",
			771 => "1111111000110010010001",
			772 => "0001011000101000100000",
			773 => "0000000000110100001100",
			774 => "0000111100101000000100",
			775 => "0000001000110010010001",
			776 => "0001001101101000000100",
			777 => "1111111000110010010001",
			778 => "0000000000110010010001",
			779 => "0011111101101100001100",
			780 => "0010001111111100000100",
			781 => "0000001000110010010001",
			782 => "0010110101010100000100",
			783 => "0000001000110010010001",
			784 => "0000001000110010010001",
			785 => "0000001101010000000100",
			786 => "1111111000110010010001",
			787 => "0000001000110010010001",
			788 => "0000100101111100001100",
			789 => "0000001010101100000100",
			790 => "1111111000110010010001",
			791 => "0011110101001000000100",
			792 => "0000001000110010010001",
			793 => "1111111000110010010001",
			794 => "0000110000100000001000",
			795 => "0001001111101000000100",
			796 => "0000001000110010010001",
			797 => "0000001000110010010001",
			798 => "1111111000110010010001",
			799 => "0011011000000100000100",
			800 => "1111111000110010010001",
			801 => "0011011000000000000100",
			802 => "0000001000110010010001",
			803 => "1111111000110010010001",
			804 => "0011110001001101001000",
			805 => "0000101101100000100100",
			806 => "0001101110111000011100",
			807 => "0011000101010100001100",
			808 => "0000100000111000000100",
			809 => "0000000000110100100101",
			810 => "0001011111011000000100",
			811 => "0000001000110100100101",
			812 => "0000000000110100100101",
			813 => "0001000001100100001100",
			814 => "0001110101111000001000",
			815 => "0001111001000100000100",
			816 => "0000000000110100100101",
			817 => "0000000000110100100101",
			818 => "0000000000110100100101",
			819 => "0000000000110100100101",
			820 => "0000011101000000000100",
			821 => "1111111000110100100101",
			822 => "0000000000110100100101",
			823 => "0011110000100000010100",
			824 => "0001010001101000010000",
			825 => "0010111010100100001000",
			826 => "0000100100111000000100",
			827 => "0000000000110100100101",
			828 => "0000000000110100100101",
			829 => "0000011101000000000100",
			830 => "0000001000110100100101",
			831 => "0000000000110100100101",
			832 => "0000000000110100100101",
			833 => "0000000101000100001000",
			834 => "0000010011110000000100",
			835 => "1111111000110100100101",
			836 => "0000000000110100100101",
			837 => "0001000000100000000100",
			838 => "0000001000110100100101",
			839 => "0000000000110100100101",
			840 => "1111111000110100100101",
			841 => "0011110001001100110000",
			842 => "0000101111100000000100",
			843 => "1111111000110110001001",
			844 => "0001010001101000100100",
			845 => "0000100101001100011000",
			846 => "0011110100000000010000",
			847 => "0001011101001000001000",
			848 => "0000000000110100000100",
			849 => "0000000000110110001001",
			850 => "0000001000110110001001",
			851 => "0001000101111000000100",
			852 => "0000000000110110001001",
			853 => "1111111000110110001001",
			854 => "0010001001000100000100",
			855 => "1111111000110110001001",
			856 => "0000000000110110001001",
			857 => "0011110100100100001000",
			858 => "0000010000011000000100",
			859 => "0000001000110110001001",
			860 => "0000001000110110001001",
			861 => "0000001000110110001001",
			862 => "0000010110110100000100",
			863 => "1111111000110110001001",
			864 => "0000001000110110001001",
			865 => "1111111000110110001001",
			866 => "0011110001001100101100",
			867 => "0000101111100000000100",
			868 => "1111111000110111100101",
			869 => "0000100011111100100100",
			870 => "0001101010001100011000",
			871 => "0000101000101100010000",
			872 => "0010101111111100001000",
			873 => "0010000101101100000100",
			874 => "0000001000110111100101",
			875 => "0000001000110111100101",
			876 => "0000000111001000000100",
			877 => "1111111000110111100101",
			878 => "0000000000110111100101",
			879 => "0001010001101000000100",
			880 => "0000001000110111100101",
			881 => "0000000000110111100101",
			882 => "0000000101000100000100",
			883 => "1111111000110111100101",
			884 => "0001000001000000000100",
			885 => "0000000000110111100101",
			886 => "1111111000110111100101",
			887 => "0000001000110111100101",
			888 => "1111111000110111100101",
			889 => "0011110001001100110100",
			890 => "0000100000111000000100",
			891 => "1111111000111001010001",
			892 => "0000100111010000100100",
			893 => "0011111101101100011000",
			894 => "0000001101100100001100",
			895 => "0000110011000000001000",
			896 => "0011111100001100000100",
			897 => "0000001000111001010001",
			898 => "0000000000111001010001",
			899 => "1111111000111001010001",
			900 => "0010111001001000001000",
			901 => "0011000101010100000100",
			902 => "0000001000111001010001",
			903 => "0000001000111001010001",
			904 => "0000001000111001010001",
			905 => "0000101110001000000100",
			906 => "1111111000111001010001",
			907 => "0000110001001000000100",
			908 => "0000001000111001010001",
			909 => "1111111000111001010001",
			910 => "0001000000100000001000",
			911 => "0000100011111100000100",
			912 => "0000001000111001010001",
			913 => "0000001000111001010001",
			914 => "1111111000111001010001",
			915 => "1111111000111001010001",
			916 => "0011110001001100111100",
			917 => "0000001000001000110100",
			918 => "0011111101101100101000",
			919 => "0000101100100000011000",
			920 => "0000010001110000001100",
			921 => "0000111100101000001000",
			922 => "0000001100001100000100",
			923 => "0000000000111011001101",
			924 => "0000001000111011001101",
			925 => "0000000000111011001101",
			926 => "0001000001110000000100",
			927 => "0000000000111011001101",
			928 => "0010101000011000000100",
			929 => "0000000000111011001101",
			930 => "1111111000111011001101",
			931 => "0001010110011100001100",
			932 => "0010001010000100001000",
			933 => "0010111010100100000100",
			934 => "0000000000111011001101",
			935 => "0000001000111011001101",
			936 => "0000000000111011001101",
			937 => "0000000000111011001101",
			938 => "0000101110101100000100",
			939 => "1111111000111011001101",
			940 => "0000001001111000000100",
			941 => "0000000000111011001101",
			942 => "0000000000111011001101",
			943 => "0001000000100000000100",
			944 => "0000001000111011001101",
			945 => "0000000000111011001101",
			946 => "1111111000111011001101",
			947 => "0011110001001100110000",
			948 => "0000100000111000000100",
			949 => "1111111000111100110001",
			950 => "0010101010011000101000",
			951 => "0000001011110100011100",
			952 => "0001010100101100010000",
			953 => "0011110111010100001000",
			954 => "0000101101000100000100",
			955 => "0000000000111100110001",
			956 => "0000001000111100110001",
			957 => "0000100001000000000100",
			958 => "1111111000111100110001",
			959 => "0000001000111100110001",
			960 => "0000100101001100000100",
			961 => "1111111000111100110001",
			962 => "0001011110010100000100",
			963 => "0000001000111100110001",
			964 => "1111111000111100110001",
			965 => "0000000111101100001000",
			966 => "0011101111100100000100",
			967 => "0000001000111100110001",
			968 => "0000001000111100110001",
			969 => "0000001000111100110001",
			970 => "1111111000111100110001",
			971 => "1111111000111100110001",
			972 => "0011110001001100111100",
			973 => "0010001010100100000100",
			974 => "0000001000111110101101",
			975 => "0000001101100100010000",
			976 => "0001101001000000001100",
			977 => "0000101001111100001000",
			978 => "0001010111100100000100",
			979 => "0000000000111110101101",
			980 => "1111111000111110101101",
			981 => "0000001000111110101101",
			982 => "1111111000111110101101",
			983 => "0001101111100100010100",
			984 => "0001010001101000010000",
			985 => "0010110011010000001000",
			986 => "0000001110010000000100",
			987 => "0000000000111110101101",
			988 => "0000000000111110101101",
			989 => "0000010110110100000100",
			990 => "0000001000111110101101",
			991 => "0000000000111110101101",
			992 => "0000000000111110101101",
			993 => "0000100000101100001100",
			994 => "0000100111000000000100",
			995 => "1111111000111110101101",
			996 => "0001001100001100000100",
			997 => "0000000000111110101101",
			998 => "0000000000111110101101",
			999 => "0001000000100000000100",
			1000 => "0000001000111110101101",
			1001 => "0000000000111110101101",
			1002 => "1111111000111110101101",
			1003 => "0011110001001101000000",
			1004 => "0011010011110000000100",
			1005 => "0000001001000000110001",
			1006 => "0000101101000100010000",
			1007 => "0000111001100000001000",
			1008 => "0000001101001000000100",
			1009 => "0000000001000000110001",
			1010 => "0000001001000000110001",
			1011 => "0010001001001100000100",
			1012 => "0000000001000000110001",
			1013 => "1111111001000000110001",
			1014 => "0011110100000000010100",
			1015 => "0000001101100100001100",
			1016 => "0001100000111000001000",
			1017 => "0000010110010000000100",
			1018 => "0000001001000000110001",
			1019 => "0000000001000000110001",
			1020 => "1111111001000000110001",
			1021 => "0010111001001000000100",
			1022 => "0000001001000000110001",
			1023 => "0000000001000000110001",
			1024 => "0000100100011000010000",
			1025 => "0010001001000100001000",
			1026 => "0000101011011100000100",
			1027 => "1111111001000000110001",
			1028 => "0000000001000000110001",
			1029 => "0000111001010100000100",
			1030 => "0000000001000000110001",
			1031 => "1111111001000000110001",
			1032 => "0001000000100000000100",
			1033 => "0000001001000000110001",
			1034 => "1111111001000000110001",
			1035 => "1111111001000000110001",
			1036 => "0011110001001100110100",
			1037 => "0000100000111000000100",
			1038 => "1111111001000010011111",
			1039 => "0010101010100100000100",
			1040 => "0000001001000010011111",
			1041 => "0000001101100100010000",
			1042 => "0001101100011100001100",
			1043 => "0000110011000000001000",
			1044 => "0000010110010000000100",
			1045 => "0000001001000010011111",
			1046 => "0000000001000010011111",
			1047 => "1111111001000010011111",
			1048 => "1111111001000010011111",
			1049 => "0011111011110000001100",
			1050 => "0001010001101000001000",
			1051 => "0001001000111000000100",
			1052 => "0000001001000010011111",
			1053 => "0000001001000010011111",
			1054 => "1111111001000010011111",
			1055 => "0000001101001100001000",
			1056 => "0011110000100000000100",
			1057 => "0000000001000010011111",
			1058 => "1111111001000010011111",
			1059 => "0001000000100000000100",
			1060 => "0000001001000010011111",
			1061 => "1111111001000010011111",
			1062 => "1111111001000010011111",
			1063 => "0011111101101100011000",
			1064 => "0000101101000100001100",
			1065 => "0000111100101000001000",
			1066 => "0000100000111000000100",
			1067 => "0000000001000011110001",
			1068 => "0000000001000011110001",
			1069 => "0000000001000011110001",
			1070 => "0001010110011100001000",
			1071 => "0010001010000100000100",
			1072 => "0000000001000011110001",
			1073 => "0000000001000011110001",
			1074 => "0000000001000011110001",
			1075 => "0000100111010000001000",
			1076 => "0000100010111100000100",
			1077 => "0000000001000011110001",
			1078 => "0000000001000011110001",
			1079 => "0000101011001000001000",
			1080 => "0001001111100000000100",
			1081 => "0000000001000011110001",
			1082 => "0000000001000011110001",
			1083 => "0000000001000011110001",
			1084 => "0011110100000000011100",
			1085 => "0000000000110100010000",
			1086 => "0011100110011100001100",
			1087 => "0010011001001000001000",
			1088 => "0000001110010100000100",
			1089 => "0000000001000101001101",
			1090 => "0000000001000101001101",
			1091 => "0000000001000101001101",
			1092 => "0000000001000101001101",
			1093 => "0010101111101000001000",
			1094 => "0010001010000100000100",
			1095 => "0000000001000101001101",
			1096 => "0000000001000101001101",
			1097 => "0000000001000101001101",
			1098 => "0000101001111000001000",
			1099 => "0011010110110100000100",
			1100 => "0000000001000101001101",
			1101 => "0000000001000101001101",
			1102 => "0001101001110000001000",
			1103 => "0000111001111100000100",
			1104 => "0000000001000101001101",
			1105 => "0000000001000101001101",
			1106 => "0000000001000101001101",
			1107 => "0011111111100000011100",
			1108 => "0000101101000100010100",
			1109 => "0000111100101000010000",
			1110 => "0000010001110000001000",
			1111 => "0000100001001000000100",
			1112 => "0000000001000110101001",
			1113 => "0000000001000110101001",
			1114 => "0001000001110000000100",
			1115 => "0000000001000110101001",
			1116 => "0000000001000110101001",
			1117 => "0000000001000110101001",
			1118 => "0000111111011000000100",
			1119 => "0000000001000110101001",
			1120 => "0000000001000110101001",
			1121 => "0000100010111100001000",
			1122 => "0010100101101100000100",
			1123 => "0000000001000110101001",
			1124 => "0000000001000110101001",
			1125 => "0011110001001100001000",
			1126 => "0001000000100000000100",
			1127 => "0000000001000110101001",
			1128 => "0000000001000110101001",
			1129 => "0000000001000110101001",
			1130 => "0011110000100000100000",
			1131 => "0000101101000100001100",
			1132 => "0000011000111100000100",
			1133 => "0000000001001000010101",
			1134 => "0001000001110000000100",
			1135 => "0000000001001000010101",
			1136 => "0000000001001000010101",
			1137 => "0011111111100000001000",
			1138 => "0001011001010100000100",
			1139 => "0000000001001000010101",
			1140 => "0000000001001000010101",
			1141 => "0000001100000100001000",
			1142 => "0000100100111000000100",
			1143 => "0000000001001000010101",
			1144 => "0000000001001000010101",
			1145 => "0000000001001000010101",
			1146 => "0011001010000100001100",
			1147 => "0010000011010000001000",
			1148 => "0001111000111000000100",
			1149 => "0000000001001000010101",
			1150 => "0000000001001000010101",
			1151 => "0000000001001000010101",
			1152 => "0001111000100000001000",
			1153 => "0001001101111100000100",
			1154 => "0000000001001000010101",
			1155 => "0000000001001000010101",
			1156 => "0000000001001000010101",
			1157 => "0001101111100100100100",
			1158 => "0000101101000100001100",
			1159 => "0000011000111100000100",
			1160 => "0000000001001010001001",
			1161 => "0001000001110000000100",
			1162 => "0000000001001010001001",
			1163 => "0000000001001010001001",
			1164 => "0011111111100000001000",
			1165 => "0001011001010100000100",
			1166 => "0000000001001010001001",
			1167 => "0000000001001010001001",
			1168 => "0000100100111000000100",
			1169 => "0000000001001010001001",
			1170 => "0000101000110100001000",
			1171 => "0001011110001100000100",
			1172 => "0000000001001010001001",
			1173 => "0000000001001010001001",
			1174 => "0000000001001010001001",
			1175 => "0011001010000100001100",
			1176 => "0010000011010000001000",
			1177 => "0001111000111000000100",
			1178 => "0000000001001010001001",
			1179 => "0000000001001010001001",
			1180 => "0000000001001010001001",
			1181 => "0001111000100000001000",
			1182 => "0001001101111100000100",
			1183 => "0000000001001010001001",
			1184 => "0000000001001010001001",
			1185 => "0000000001001010001001",
			1186 => "0011111101000100101100",
			1187 => "0000100111100000011100",
			1188 => "0001101001000000010000",
			1189 => "0000100000111000000100",
			1190 => "0000000001001011111101",
			1191 => "0000110011000000001000",
			1192 => "0010000101011100000100",
			1193 => "0000000001001011111101",
			1194 => "0000000001001011111101",
			1195 => "0000000001001011111101",
			1196 => "0000000111001000000100",
			1197 => "1111111001001011111101",
			1198 => "0011111010100000000100",
			1199 => "0000000001001011111101",
			1200 => "0000000001001011111101",
			1201 => "0011110000100000001000",
			1202 => "0001010001101000000100",
			1203 => "0000001001001011111101",
			1204 => "0000000001001011111101",
			1205 => "0000100111000000000100",
			1206 => "0000000001001011111101",
			1207 => "0000000001001011111101",
			1208 => "0010111000000100001000",
			1209 => "0011000110001100000100",
			1210 => "0000000001001011111101",
			1211 => "1111111001001011111101",
			1212 => "0010011111101000000100",
			1213 => "0000000001001011111101",
			1214 => "0000000001001011111101",
			1215 => "0000101101000100010000",
			1216 => "0001110101011100001000",
			1217 => "0011111000000100000100",
			1218 => "0000000001001101100001",
			1219 => "0000000001001101100001",
			1220 => "0001001001100100000100",
			1221 => "0000000001001101100001",
			1222 => "0000000001001101100001",
			1223 => "0011110110100000011100",
			1224 => "0001010001101000010100",
			1225 => "0001000111110000000100",
			1226 => "0000000001001101100001",
			1227 => "0000101101100000001100",
			1228 => "0000101111110000000100",
			1229 => "0000000001001101100001",
			1230 => "0000000111001000000100",
			1231 => "0000000001001101100001",
			1232 => "0000000001001101100001",
			1233 => "0000000001001101100001",
			1234 => "0011011001001000000100",
			1235 => "0000000001001101100001",
			1236 => "0000000001001101100001",
			1237 => "0011011000000100000100",
			1238 => "0000000001001101100001",
			1239 => "0000000001001101100001",
			1240 => "0001101001110000101000",
			1241 => "0000001101100100010100",
			1242 => "0011111010011100010000",
			1243 => "0001010011000000001100",
			1244 => "0000100000111000000100",
			1245 => "0000000001001110110101",
			1246 => "0010111100101000000100",
			1247 => "0000000001001110110101",
			1248 => "0000000001001110110101",
			1249 => "0000000001001110110101",
			1250 => "0000000001001110110101",
			1251 => "0001010001101000001100",
			1252 => "0011110100100100000100",
			1253 => "0000000001001110110101",
			1254 => "0001101010011000000100",
			1255 => "0000000001001110110101",
			1256 => "0000000001001110110101",
			1257 => "0000100100111100000100",
			1258 => "0000000001001110110101",
			1259 => "0000000001001110110101",
			1260 => "0000000001001110110101",
			1261 => "0000001101100100010100",
			1262 => "0011111010011100010000",
			1263 => "0001010011000000001100",
			1264 => "0000100000111000000100",
			1265 => "0000000001010000110001",
			1266 => "0010111100101000000100",
			1267 => "0000000001010000110001",
			1268 => "0000000001010000110001",
			1269 => "0000000001010000110001",
			1270 => "0000000001010000110001",
			1271 => "0011110100100100010100",
			1272 => "0001010001101000001100",
			1273 => "0010111001001000000100",
			1274 => "0000000001010000110001",
			1275 => "0010110101101100000100",
			1276 => "0000000001010000110001",
			1277 => "0000000001010000110001",
			1278 => "0001011101111100000100",
			1279 => "0000000001010000110001",
			1280 => "0000000001010000110001",
			1281 => "0011001010000100001100",
			1282 => "0010000011010000001000",
			1283 => "0001111000111000000100",
			1284 => "0000000001010000110001",
			1285 => "0000000001010000110001",
			1286 => "0000000001010000110001",
			1287 => "0001111000100000001000",
			1288 => "0000101011011000000100",
			1289 => "0000000001010000110001",
			1290 => "0000000001010000110001",
			1291 => "0000000001010000110001",
			1292 => "0011110100100100110000",
			1293 => "0000100010110000011000",
			1294 => "0011111010011100010100",
			1295 => "0000010001110000001000",
			1296 => "0000001110010100000100",
			1297 => "0000000001010010110101",
			1298 => "0000000001010010110101",
			1299 => "0001010110001100001000",
			1300 => "0000001010011100000100",
			1301 => "0000000001010010110101",
			1302 => "0000000001010010110101",
			1303 => "0000000001010010110101",
			1304 => "0000000001010010110101",
			1305 => "0001010001101000010000",
			1306 => "0010111010100100001000",
			1307 => "0010111110011000000100",
			1308 => "0000000001010010110101",
			1309 => "0000000001010010110101",
			1310 => "0011011001000100000100",
			1311 => "0000000001010010110101",
			1312 => "0000000001010010110101",
			1313 => "0010010011000000000100",
			1314 => "0000000001010010110101",
			1315 => "0000000001010010110101",
			1316 => "0010000011010000001000",
			1317 => "0001111000111000000100",
			1318 => "0000000001010010110101",
			1319 => "0000000001010010110101",
			1320 => "0010111010000100000100",
			1321 => "0000000001010010110101",
			1322 => "0001111000100000000100",
			1323 => "0000000001010010110101",
			1324 => "0000000001010010110101",
			1325 => "0001100000010100101000",
			1326 => "0000100000111000000100",
			1327 => "0000000001010100010001",
			1328 => "0001011100011100010000",
			1329 => "0011011010000100001100",
			1330 => "0001101001101100000100",
			1331 => "0000000001010100010001",
			1332 => "0001101111100000000100",
			1333 => "0000000001010100010001",
			1334 => "0000000001010100010001",
			1335 => "0000000001010100010001",
			1336 => "0001000110011100001000",
			1337 => "0000111000100000000100",
			1338 => "0000000001010100010001",
			1339 => "0000000001010100010001",
			1340 => "0010100000111100000100",
			1341 => "0000000001010100010001",
			1342 => "0001001101111100000100",
			1343 => "0000000001010100010001",
			1344 => "0000000001010100010001",
			1345 => "0011011000000100000100",
			1346 => "0000000001010100010001",
			1347 => "0000000001010100010001",
			1348 => "0011110110100000110000",
			1349 => "0000000110100000010000",
			1350 => "0011011101000000000100",
			1351 => "0000000001010101111101",
			1352 => "0001110101011100001000",
			1353 => "0001100011000000000100",
			1354 => "0000000001010101111101",
			1355 => "0000000001010101111101",
			1356 => "0000000001010101111101",
			1357 => "0011111111100000001000",
			1358 => "0001011001010100000100",
			1359 => "0000000001010101111101",
			1360 => "0000000001010101111101",
			1361 => "0010110101010100010000",
			1362 => "0011010110110100001000",
			1363 => "0010101000111000000100",
			1364 => "0000000001010101111101",
			1365 => "0000000001010101111101",
			1366 => "0001000001011000000100",
			1367 => "0000000001010101111101",
			1368 => "0000000001010101111101",
			1369 => "0001111000100000000100",
			1370 => "0000000001010101111101",
			1371 => "0000000001010101111101",
			1372 => "0011011000000100000100",
			1373 => "0000000001010101111101",
			1374 => "0000000001010101111101",
			1375 => "0001101001110000110000",
			1376 => "0000101101000100010000",
			1377 => "0001101001011000001100",
			1378 => "0000100000111000000100",
			1379 => "0000000001010111100001",
			1380 => "0010100101101100000100",
			1381 => "0000000001010111100001",
			1382 => "0000000001010111100001",
			1383 => "0000000001010111100001",
			1384 => "0001011100011100001100",
			1385 => "0001101001101100000100",
			1386 => "0000000001010111100001",
			1387 => "0000100001000000000100",
			1388 => "0000000001010111100001",
			1389 => "0000000001010111100001",
			1390 => "0000001000001000001100",
			1391 => "0010000101011100001000",
			1392 => "0011011011101100000100",
			1393 => "0000000001010111100001",
			1394 => "0000000001010111100001",
			1395 => "0000000001010111100001",
			1396 => "0001000000100000000100",
			1397 => "0000000001010111100001",
			1398 => "0000000001010111100001",
			1399 => "0000000001010111100001",
			1400 => "0001111000000000101000",
			1401 => "0000101101101100001000",
			1402 => "0011011101000000000100",
			1403 => "1101101001011001110101",
			1404 => "1101011001011001110101",
			1405 => "0010101111111100001000",
			1406 => "0010010101011100000100",
			1407 => "1110011001011001110101",
			1408 => "1110110001011001110101",
			1409 => "0000101000110100001100",
			1410 => "0001100001101000001000",
			1411 => "0000101101000100000100",
			1412 => "1101011001011001110101",
			1413 => "1110010001011001110101",
			1414 => "1101011001011001110101",
			1415 => "0001101111100100000100",
			1416 => "1110110001011001110101",
			1417 => "0001100010010100000100",
			1418 => "1101111001011001110101",
			1419 => "1101011001011001110101",
			1420 => "0011111001110000011000",
			1421 => "0000101011011100010000",
			1422 => "0000100001100000001000",
			1423 => "0000100001000000000100",
			1424 => "1101011001011001110101",
			1425 => "1101100001011001110101",
			1426 => "0000111111101000000100",
			1427 => "1110101001011001110101",
			1428 => "1101011001011001110101",
			1429 => "0001000000111100000100",
			1430 => "1110110001011001110101",
			1431 => "1101101001011001110101",
			1432 => "0001101001110000001000",
			1433 => "0000100100111100000100",
			1434 => "1101011001011001110101",
			1435 => "1101100001011001110101",
			1436 => "1101011001011001110101",
			1437 => "0011111001110000110000",
			1438 => "0000100001100000100000",
			1439 => "0011010011110000000100",
			1440 => "0000000001011011101001",
			1441 => "0011111010011100001100",
			1442 => "0000101101101100000100",
			1443 => "0000000001011011101001",
			1444 => "0000110011000000000100",
			1445 => "0000000001011011101001",
			1446 => "0000000001011011101001",
			1447 => "0000001101100100000100",
			1448 => "0000000001011011101001",
			1449 => "0011011011101100000100",
			1450 => "0000000001011011101001",
			1451 => "0010110101010100000100",
			1452 => "0000000001011011101001",
			1453 => "0000000001011011101001",
			1454 => "0011110100100100001000",
			1455 => "0001011110010100000100",
			1456 => "0000000001011011101001",
			1457 => "0000000001011011101001",
			1458 => "0011110010010100000100",
			1459 => "0000000001011011101001",
			1460 => "0000000001011011101001",
			1461 => "0000011000111100000100",
			1462 => "0000000001011011101001",
			1463 => "0011011000000100000100",
			1464 => "0000000001011011101001",
			1465 => "0000000001011011101001",
			1466 => "0001100000010100101100",
			1467 => "0000101000010100100000",
			1468 => "0001101111100000011100",
			1469 => "0000101101000100010000",
			1470 => "0001101001011000001100",
			1471 => "0000100000111000000100",
			1472 => "0000000001011101001101",
			1473 => "0010100110000000000100",
			1474 => "0000000001011101001101",
			1475 => "0000000001011101001101",
			1476 => "0000000001011101001101",
			1477 => "0001000101111000001000",
			1478 => "0010001111001000000100",
			1479 => "0000000001011101001101",
			1480 => "0000000001011101001101",
			1481 => "0000000001011101001101",
			1482 => "0000000001011101001101",
			1483 => "0000111001000000000100",
			1484 => "0000000001011101001101",
			1485 => "0000111110001100000100",
			1486 => "0000000001011101001101",
			1487 => "0000000001011101001101",
			1488 => "0011011000000100000100",
			1489 => "0000000001011101001101",
			1490 => "0000000001011101001101",
			1491 => "0001100000010100101100",
			1492 => "0000100010111100101000",
			1493 => "0011110001010100010100",
			1494 => "0000111111011000001100",
			1495 => "0000100000111000000100",
			1496 => "0000000001011110110001",
			1497 => "0011010101010100000100",
			1498 => "0000000001011110110001",
			1499 => "0000000001011110110001",
			1500 => "0010101001010100000100",
			1501 => "0000000001011110110001",
			1502 => "0000000001011110110001",
			1503 => "0000101101100100000100",
			1504 => "0000000001011110110001",
			1505 => "0011111101101100001000",
			1506 => "0010110101011100000100",
			1507 => "0000000001011110110001",
			1508 => "0000000001011110110001",
			1509 => "0011010110001100000100",
			1510 => "0000000001011110110001",
			1511 => "0000000001011110110001",
			1512 => "0000000001011110110001",
			1513 => "0011011000000100000100",
			1514 => "0000000001011110110001",
			1515 => "0000000001011110110001",
			1516 => "0001101001110000110100",
			1517 => "0000100101001100100100",
			1518 => "0011110001010100011000",
			1519 => "0000111111011000010000",
			1520 => "0000100000111000000100",
			1521 => "0000000001100000011101",
			1522 => "0000101101000100001000",
			1523 => "0001101111101000000100",
			1524 => "0000000001100000011101",
			1525 => "0000000001100000011101",
			1526 => "0000001001100000011101",
			1527 => "0001110011001000000100",
			1528 => "0000000001100000011101",
			1529 => "0000000001100000011101",
			1530 => "0000101101100100000100",
			1531 => "1111111001100000011101",
			1532 => "0011111101101100000100",
			1533 => "0000000001100000011101",
			1534 => "0000000001100000011101",
			1535 => "0001010001101000001000",
			1536 => "0011110100100100000100",
			1537 => "0000001001100000011101",
			1538 => "0000000001100000011101",
			1539 => "0000100100111100000100",
			1540 => "0000000001100000011101",
			1541 => "0000000001100000011101",
			1542 => "1111111001100000011101",
			1543 => "0001101001110000111000",
			1544 => "0000101101000100010100",
			1545 => "0011101001010000001100",
			1546 => "0000100000111000000100",
			1547 => "0000000001100010010001",
			1548 => "0011011011101100000100",
			1549 => "0000000001100010010001",
			1550 => "0000000001100010010001",
			1551 => "0001111010000100000100",
			1552 => "0000000001100010010001",
			1553 => "0000000001100010010001",
			1554 => "0011111111100000001100",
			1555 => "0001011001010100001000",
			1556 => "0010001010000100000100",
			1557 => "0000001001100010010001",
			1558 => "0000000001100010010001",
			1559 => "0000000001100010010001",
			1560 => "0000100101001100001000",
			1561 => "0001000101010100000100",
			1562 => "0000000001100010010001",
			1563 => "0000000001100010010001",
			1564 => "0001010001101000001000",
			1565 => "0011110100100100000100",
			1566 => "0000001001100010010001",
			1567 => "0000000001100010010001",
			1568 => "0000100100111100000100",
			1569 => "0000000001100010010001",
			1570 => "0000000001100010010001",
			1571 => "0000000001100010010001",
			1572 => "0011110001001100110000",
			1573 => "0000101101100000011000",
			1574 => "0010101110011000001000",
			1575 => "0000001010100000000100",
			1576 => "0000000001100011110101",
			1577 => "0000000001100011110101",
			1578 => "0010110110001100000100",
			1579 => "0000000001100011110101",
			1580 => "0001101110111000001000",
			1581 => "0001100011000100000100",
			1582 => "0000000001100011110101",
			1583 => "0000000001100011110101",
			1584 => "0000000001100011110101",
			1585 => "0001001101111100010100",
			1586 => "0010011100101000000100",
			1587 => "0000000001100011110101",
			1588 => "0001011100110100000100",
			1589 => "0000000001100011110101",
			1590 => "0001011010100000001000",
			1591 => "0001010001101000000100",
			1592 => "0000000001100011110101",
			1593 => "0000000001100011110101",
			1594 => "0000000001100011110101",
			1595 => "0000000001100011110101",
			1596 => "0000000001100011110101",
			1597 => "0011110001001100111100",
			1598 => "0000100101001100101000",
			1599 => "0011110001010100010100",
			1600 => "0000111111011000001100",
			1601 => "0000100000111000000100",
			1602 => "0000000001100101110001",
			1603 => "0011111100001100000100",
			1604 => "0000001001100101110001",
			1605 => "0000000001100101110001",
			1606 => "0001110011001000000100",
			1607 => "0000000001100101110001",
			1608 => "0000000001100101110001",
			1609 => "0010110101010100001100",
			1610 => "0000101110010000001000",
			1611 => "0000010011110000000100",
			1612 => "1111111001100101110001",
			1613 => "0000000001100101110001",
			1614 => "0000000001100101110001",
			1615 => "0000110110101100000100",
			1616 => "0000000001100101110001",
			1617 => "0000000001100101110001",
			1618 => "0001010001101000001000",
			1619 => "0011110100100100000100",
			1620 => "0000001001100101110001",
			1621 => "0000000001100101110001",
			1622 => "0000100100111100000100",
			1623 => "0000000001100101110001",
			1624 => "0000110001000100000100",
			1625 => "0000000001100101110001",
			1626 => "0000000001100101110001",
			1627 => "1111111001100101110001",
			1628 => "0011110001001100110100",
			1629 => "0000101000010100100100",
			1630 => "0011111101101100011100",
			1631 => "0000101100100000010000",
			1632 => "0001100001011000001100",
			1633 => "0000100000111000000100",
			1634 => "0000000001100111011101",
			1635 => "0010011001001000000100",
			1636 => "0000001001100111011101",
			1637 => "0000000001100111011101",
			1638 => "1111111001100111011101",
			1639 => "0001001000000100001000",
			1640 => "0010110011010000000100",
			1641 => "0000000001100111011101",
			1642 => "0000001001100111011101",
			1643 => "0000000001100111011101",
			1644 => "0010111100101000000100",
			1645 => "1111111001100111011101",
			1646 => "0000000001100111011101",
			1647 => "0001010001101000000100",
			1648 => "0000001001100111011101",
			1649 => "0000100100111100000100",
			1650 => "0000000001100111011101",
			1651 => "0001010000001000000100",
			1652 => "0000000001100111011101",
			1653 => "0000000001100111011101",
			1654 => "1111111001100111011101",
			1655 => "0011110001001100101000",
			1656 => "0000101111100000000100",
			1657 => "1111111001101000110001",
			1658 => "0001010001101000011100",
			1659 => "0000101100111000010100",
			1660 => "0011111101101100010000",
			1661 => "0000100010110000001000",
			1662 => "0000110011000000000100",
			1663 => "0000000001101000110001",
			1664 => "1111111001101000110001",
			1665 => "0001001000111000000100",
			1666 => "0000001001101000110001",
			1667 => "0000000001101000110001",
			1668 => "1111111001101000110001",
			1669 => "0000100111000000000100",
			1670 => "0000000001101000110001",
			1671 => "0000001001101000110001",
			1672 => "0000100100111100000100",
			1673 => "1111111001101000110001",
			1674 => "0000001001101000110001",
			1675 => "1111111001101000110001",
			1676 => "0011110001001100111000",
			1677 => "0000101100100000010000",
			1678 => "0011110001011000001100",
			1679 => "0000100000111000000100",
			1680 => "0000000001101010100101",
			1681 => "0010011001001000000100",
			1682 => "0000000001101010100101",
			1683 => "0000000001101010100101",
			1684 => "0000000001101010100101",
			1685 => "0001100001111100001100",
			1686 => "0001011001010100001000",
			1687 => "0010001010000100000100",
			1688 => "0000001001101010100101",
			1689 => "0000000001101010100101",
			1690 => "0000000001101010100101",
			1691 => "0000101000010100001100",
			1692 => "0011111101101100001000",
			1693 => "0000100100010000000100",
			1694 => "0000000001101010100101",
			1695 => "0000000001101010100101",
			1696 => "0000000001101010100101",
			1697 => "0001000000100000001100",
			1698 => "0000100101111100001000",
			1699 => "0011110100100100000100",
			1700 => "0000000001101010100101",
			1701 => "0000000001101010100101",
			1702 => "0000000001101010100101",
			1703 => "0000000001101010100101",
			1704 => "0000000001101010100101",
			1705 => "0011111001110000110100",
			1706 => "0000101000110100101000",
			1707 => "0001011001010100100000",
			1708 => "0011010011110000000100",
			1709 => "0000000001101100100001",
			1710 => "0000101101000100001100",
			1711 => "0000111001100000001000",
			1712 => "0011000101010100000100",
			1713 => "0000000001101100100001",
			1714 => "0000000001101100100001",
			1715 => "0000000001101100100001",
			1716 => "0010011001000100001000",
			1717 => "0001100010111000000100",
			1718 => "0000000001101100100001",
			1719 => "0000000001101100100001",
			1720 => "0000010001100100000100",
			1721 => "0000000001101100100001",
			1722 => "0000000001101100100001",
			1723 => "0001000101111000000100",
			1724 => "0000000001101100100001",
			1725 => "0000000001101100100001",
			1726 => "0011110100100100000100",
			1727 => "0000000001101100100001",
			1728 => "0011110010010100000100",
			1729 => "0000000001101100100001",
			1730 => "0000000001101100100001",
			1731 => "0000011000111100000100",
			1732 => "0000000001101100100001",
			1733 => "0011011000000100000100",
			1734 => "0000000001101100100001",
			1735 => "0000000001101100100001",
			1736 => "0011110001001100111100",
			1737 => "0000101101000100010000",
			1738 => "0010000011010000000100",
			1739 => "0000000001101110011101",
			1740 => "0001000001110000000100",
			1741 => "0000000001101110011101",
			1742 => "0010010011010000000100",
			1743 => "1111111001101110011101",
			1744 => "1111111001101110011101",
			1745 => "0011110100000000010000",
			1746 => "0000100010110000001000",
			1747 => "0001101110001100000100",
			1748 => "0000001001101110011101",
			1749 => "1111111001101110011101",
			1750 => "0001000011000000000100",
			1751 => "0000001001101110011101",
			1752 => "0000001001101110011101",
			1753 => "0000100010111100001100",
			1754 => "0001101111100100001000",
			1755 => "0000101000101100000100",
			1756 => "1111111001101110011101",
			1757 => "0000001001101110011101",
			1758 => "1111111001101110011101",
			1759 => "0001000000100000001100",
			1760 => "0000101001111000001000",
			1761 => "0011111001110000000100",
			1762 => "0000001001101110011101",
			1763 => "1111111001101110011101",
			1764 => "0000001001101110011101",
			1765 => "1111111001101110011101",
			1766 => "1111111001101110011101",
			1767 => "0011110001001100111000",
			1768 => "0000100001100000100100",
			1769 => "0011010011110000000100",
			1770 => "0000001001110000010001",
			1771 => "0011110001010100010100",
			1772 => "0000101101000100001100",
			1773 => "0000110110001100001000",
			1774 => "0000000000111100000100",
			1775 => "0000000001110000010001",
			1776 => "0000001001110000010001",
			1777 => "1111111001110000010001",
			1778 => "0000010110010000000100",
			1779 => "0000001001110000010001",
			1780 => "0000000001110000010001",
			1781 => "0000100111100000000100",
			1782 => "1111111001110000010001",
			1783 => "0001001001010100000100",
			1784 => "0000000001110000010001",
			1785 => "0000000001110000010001",
			1786 => "0011110000100000000100",
			1787 => "0000001001110000010001",
			1788 => "0000000101000100001000",
			1789 => "0010001001000100000100",
			1790 => "1111111001110000010001",
			1791 => "0000000001110000010001",
			1792 => "0001000000100000000100",
			1793 => "0000001001110000010001",
			1794 => "0000000001110000010001",
			1795 => "1111111001110000010001",
			1796 => "0001100000010100111100",
			1797 => "0000101111100000001000",
			1798 => "0011011101000000000100",
			1799 => "0000000001110010011101",
			1800 => "1111111001110010011101",
			1801 => "0001011110111000100100",
			1802 => "0000101101100100010100",
			1803 => "0001011001001000001100",
			1804 => "0011110011110100001000",
			1805 => "0010011001001000000100",
			1806 => "0000011001110010011101",
			1807 => "0000010001110010011101",
			1808 => "0000001001110010011101",
			1809 => "0000010001110000000100",
			1810 => "0000001001110010011101",
			1811 => "1111111001110010011101",
			1812 => "0001101010001100001100",
			1813 => "0001101101111100001000",
			1814 => "0010011010000100000100",
			1815 => "0000010001110010011101",
			1816 => "0000011001110010011101",
			1817 => "0000010001110010011101",
			1818 => "0000010001110010011101",
			1819 => "0000100000100100001100",
			1820 => "0000010000011000001000",
			1821 => "0001011110010100000100",
			1822 => "0000001001110010011101",
			1823 => "1111111001110010011101",
			1824 => "1111111001110010011101",
			1825 => "0000010001110010011101",
			1826 => "0011011000000100000100",
			1827 => "1111111001110010011101",
			1828 => "0011100001100000000100",
			1829 => "0000000001110010011101",
			1830 => "1111111001110010011101",
			1831 => "0011110001001100110100",
			1832 => "0000100000111000000100",
			1833 => "1111111001110100001001",
			1834 => "0001010100101100011100",
			1835 => "0011110111010100010000",
			1836 => "0000101100100000001100",
			1837 => "0000111100101000000100",
			1838 => "0000001001110100001001",
			1839 => "0001011101001000000100",
			1840 => "1111111001110100001001",
			1841 => "0000000001110100001001",
			1842 => "0000001001110100001001",
			1843 => "0000100001000000000100",
			1844 => "1111111001110100001001",
			1845 => "0010001111111100000100",
			1846 => "0000000001110100001001",
			1847 => "0000001001110100001001",
			1848 => "0000001000001000001100",
			1849 => "0011101010100000001000",
			1850 => "0000001100000100000100",
			1851 => "1111111001110100001001",
			1852 => "0000001001110100001001",
			1853 => "1111111001110100001001",
			1854 => "0001000000100000000100",
			1855 => "0000001001110100001001",
			1856 => "1111111001110100001001",
			1857 => "1111111001110100001001",
			1858 => "0001100000010101000000",
			1859 => "0000101111100000001000",
			1860 => "0000011000111100000100",
			1861 => "0000000001110110011101",
			1862 => "1111111001110110011101",
			1863 => "0001010011110100101000",
			1864 => "0000000010110100010100",
			1865 => "0010100101011100001000",
			1866 => "0001101011000000000100",
			1867 => "0000100001110110011101",
			1868 => "0000011001110110011101",
			1869 => "0000010001110000000100",
			1870 => "0000001001110110011101",
			1871 => "0000111101101000000100",
			1872 => "0000000001110110011101",
			1873 => "1111111001110110011101",
			1874 => "0000100101001100001100",
			1875 => "0011111101101100001000",
			1876 => "0001001011101100000100",
			1877 => "0000011001110110011101",
			1878 => "0000100001110110011101",
			1879 => "1111111001110110011101",
			1880 => "0011111111111000000100",
			1881 => "0000011001110110011101",
			1882 => "0000100001110110011101",
			1883 => "0000001011011000001100",
			1884 => "0011101010100000001000",
			1885 => "0010000101011100000100",
			1886 => "0000000001110110011101",
			1887 => "1111111001110110011101",
			1888 => "1111111001110110011101",
			1889 => "0000011001110110011101",
			1890 => "0011011000000100000100",
			1891 => "1111111001110110011101",
			1892 => "0000110011000100000100",
			1893 => "1111111001110110011101",
			1894 => "0000000001110110011101",
			1895 => "0011110110100000111100",
			1896 => "0000100000111000000100",
			1897 => "1111111001111000101001",
			1898 => "0001011000101000100000",
			1899 => "0000101101000100001000",
			1900 => "0000111100101000000100",
			1901 => "0000001001111000101001",
			1902 => "1111111001111000101001",
			1903 => "0001101101111100001100",
			1904 => "0000010111110000000100",
			1905 => "0000001001111000101001",
			1906 => "0000000011101100000100",
			1907 => "0000001001111000101001",
			1908 => "0000001001111000101001",
			1909 => "0000101110010000000100",
			1910 => "1111111001111000101001",
			1911 => "0000010111100100000100",
			1912 => "0000001001111000101001",
			1913 => "0000001001111000101001",
			1914 => "0000100101111100001100",
			1915 => "0000001010101100000100",
			1916 => "1111111001111000101001",
			1917 => "0011110101001000000100",
			1918 => "0000001001111000101001",
			1919 => "1111111001111000101001",
			1920 => "0000110000100000001000",
			1921 => "0001001111101000000100",
			1922 => "0000001001111000101001",
			1923 => "0000010001111000101001",
			1924 => "1111111001111000101001",
			1925 => "0011011000000100000100",
			1926 => "1111111001111000101001",
			1927 => "0001101010110000000100",
			1928 => "0000000001111000101001",
			1929 => "1111111001111000101001",
			1930 => "0011110001001101000000",
			1931 => "0000011001100100010000",
			1932 => "0000110001001000001100",
			1933 => "0001001110011000001000",
			1934 => "0001110011000000000100",
			1935 => "0000000001111010101101",
			1936 => "0000000001111010101101",
			1937 => "0000001001111010101101",
			1938 => "0000000001111010101101",
			1939 => "0000001101100100010100",
			1940 => "0001011001001000010000",
			1941 => "0010001001001100000100",
			1942 => "0000000001111010101101",
			1943 => "0011001110011000000100",
			1944 => "0000000001111010101101",
			1945 => "0010011010000100000100",
			1946 => "0000000001111010101101",
			1947 => "0000000001111010101101",
			1948 => "1111111001111010101101",
			1949 => "0001010100101100001000",
			1950 => "0010111010100100000100",
			1951 => "0000000001111010101101",
			1952 => "0000001001111010101101",
			1953 => "0000000101000100001100",
			1954 => "0010001001001100000100",
			1955 => "0000000001111010101101",
			1956 => "0011011100101000000100",
			1957 => "1111111001111010101101",
			1958 => "0000000001111010101101",
			1959 => "0001000000100000000100",
			1960 => "0000001001111010101101",
			1961 => "0000000001111010101101",
			1962 => "1111111001111010101101",
			1963 => "0011110001001100111100",
			1964 => "0000101000010100101100",
			1965 => "0011110100000000100100",
			1966 => "0000101100100000010100",
			1967 => "0011110011110100010000",
			1968 => "0010011001001000001000",
			1969 => "0000001110010100000100",
			1970 => "0000000001111100101001",
			1971 => "0000001001111100101001",
			1972 => "0010000101011100000100",
			1973 => "0000000001111100101001",
			1974 => "0000000001111100101001",
			1975 => "1111111001111100101001",
			1976 => "0010001010000100001100",
			1977 => "0001001000000100001000",
			1978 => "0011111111100000000100",
			1979 => "0000001001111100101001",
			1980 => "0000000001111100101001",
			1981 => "0000000001111100101001",
			1982 => "0000000001111100101001",
			1983 => "0011010101011100000100",
			1984 => "1111111001111100101001",
			1985 => "0000000001111100101001",
			1986 => "0001000000100000001100",
			1987 => "0011111001110000000100",
			1988 => "0000001001111100101001",
			1989 => "0011111111000100000100",
			1990 => "0000000001111100101001",
			1991 => "0000000001111100101001",
			1992 => "0000000001111100101001",
			1993 => "1111111001111100101001",
			1994 => "0011110001001100111000",
			1995 => "0000101111100000000100",
			1996 => "1111111001111110011101",
			1997 => "0001011110111000100100",
			1998 => "0000001101100100010000",
			1999 => "0010100101011100001000",
			2000 => "0001110110000000000100",
			2001 => "0000001001111110011101",
			2002 => "0000001001111110011101",
			2003 => "0011010110001100000100",
			2004 => "0000000001111110011101",
			2005 => "1111111001111110011101",
			2006 => "0011111111100100001000",
			2007 => "0000001000110100000100",
			2008 => "0000001001111110011101",
			2009 => "0000001001111110011101",
			2010 => "0000000101111100000100",
			2011 => "1111111001111110011101",
			2012 => "0001101010110100000100",
			2013 => "0000001001111110011101",
			2014 => "0000001001111110011101",
			2015 => "0000000011100000001100",
			2016 => "0011110100100100001000",
			2017 => "0000100101001100000100",
			2018 => "1111111001111110011101",
			2019 => "0000001001111110011101",
			2020 => "1111111001111110011101",
			2021 => "0000001001111110011101",
			2022 => "1111111001111110011101",
			2023 => "0011110001001100111100",
			2024 => "0000001000001000110100",
			2025 => "0011111101101100101000",
			2026 => "0000101100100000011000",
			2027 => "0000010001110000001100",
			2028 => "0000111100101000001000",
			2029 => "0000001100001100000100",
			2030 => "0000000010000000011001",
			2031 => "0000001010000000011001",
			2032 => "0000000010000000011001",
			2033 => "0001000001110000000100",
			2034 => "0000000010000000011001",
			2035 => "0010101000011000000100",
			2036 => "0000000010000000011001",
			2037 => "1111111010000000011001",
			2038 => "0001010110011100001100",
			2039 => "0010111010100100000100",
			2040 => "0000000010000000011001",
			2041 => "0010001010000100000100",
			2042 => "0000001010000000011001",
			2043 => "0000000010000000011001",
			2044 => "0000000010000000011001",
			2045 => "0000101011011100000100",
			2046 => "1111111010000000011001",
			2047 => "0000001001111000000100",
			2048 => "0000000010000000011001",
			2049 => "0000000010000000011001",
			2050 => "0001000000100000000100",
			2051 => "0000001010000000011001",
			2052 => "0000000010000000011001",
			2053 => "1111111010000000011001",
			2054 => "0011110001001100110000",
			2055 => "0000100000111000000100",
			2056 => "1111111010000001111101",
			2057 => "0011010011110000000100",
			2058 => "0000001010000001111101",
			2059 => "0000101101000100001100",
			2060 => "0001101011111000001000",
			2061 => "0001010101101100000100",
			2062 => "0000000010000001111101",
			2063 => "1111111010000001111101",
			2064 => "1111111010000001111101",
			2065 => "0001100001111100001100",
			2066 => "0000000111001000001000",
			2067 => "0000110011000000000100",
			2068 => "0000001010000001111101",
			2069 => "1111111010000001111101",
			2070 => "0000001010000001111101",
			2071 => "0000100101001100001000",
			2072 => "0001000101010100000100",
			2073 => "0000000010000001111101",
			2074 => "1111111010000001111101",
			2075 => "0011110100100100000100",
			2076 => "0000001010000001111101",
			2077 => "0000000010000001111101",
			2078 => "1111111010000001111101",
			2079 => "0011110001001100111100",
			2080 => "0010001011101100000100",
			2081 => "0000001010000011111001",
			2082 => "0000101101100000010100",
			2083 => "0011111100011100010000",
			2084 => "0000101111100000000100",
			2085 => "1111111010000011111001",
			2086 => "0000110011000000001000",
			2087 => "0010000101011100000100",
			2088 => "0000001010000011111001",
			2089 => "0000000010000011111001",
			2090 => "0000000010000011111001",
			2091 => "1111111010000011111001",
			2092 => "0001101111100100010100",
			2093 => "0001010001101000010000",
			2094 => "0010111010100100001000",
			2095 => "0000100100111000000100",
			2096 => "0000000010000011111001",
			2097 => "0000000010000011111001",
			2098 => "0000010110110100000100",
			2099 => "0000001010000011111001",
			2100 => "0000000010000011111001",
			2101 => "0000000010000011111001",
			2102 => "0000000101000100001000",
			2103 => "0000100111000000000100",
			2104 => "1111111010000011111001",
			2105 => "0000000010000011111001",
			2106 => "0001000000100000000100",
			2107 => "0000001010000011111001",
			2108 => "0000000010000011111001",
			2109 => "1111111010000011111001",
			2110 => "0011110001001101000000",
			2111 => "0010001010100100000100",
			2112 => "0000001010000101111111",
			2113 => "0000000110100000010000",
			2114 => "0001000001110000001000",
			2115 => "0011101010000100000100",
			2116 => "0000000010000101111111",
			2117 => "0000000010000101111111",
			2118 => "0010001001001100000100",
			2119 => "0000000010000101111111",
			2120 => "1111111010000101111111",
			2121 => "0011110100000000010100",
			2122 => "0000001101100100001100",
			2123 => "0001101100011100001000",
			2124 => "0011000111011100000100",
			2125 => "0000001010000101111111",
			2126 => "0000000010000101111111",
			2127 => "1111111010000101111111",
			2128 => "0010111001001000000100",
			2129 => "0000001010000101111111",
			2130 => "0000000010000101111111",
			2131 => "0000101100111100010000",
			2132 => "0010001001000100001000",
			2133 => "0000101011011100000100",
			2134 => "1111111010000101111111",
			2135 => "0000000010000101111111",
			2136 => "0001011011111000000100",
			2137 => "0000000010000101111111",
			2138 => "1111111010000101111111",
			2139 => "0001000000100000000100",
			2140 => "0000001010000101111111",
			2141 => "0000000010000101111111",
			2142 => "1111111010000101111111",
			2143 => "0001010011000000011000",
			2144 => "0011110101110000010000",
			2145 => "0000100000111000000100",
			2146 => "0000000010000111011001",
			2147 => "0010001010000100001000",
			2148 => "0000111101101000000100",
			2149 => "0000000010000111011001",
			2150 => "0000000010000111011001",
			2151 => "0000000010000111011001",
			2152 => "0000000101100000000100",
			2153 => "0000000010000111011001",
			2154 => "0000000010000111011001",
			2155 => "0000001010101100001100",
			2156 => "0010011010000100000100",
			2157 => "0000000010000111011001",
			2158 => "0001000101111000000100",
			2159 => "0000000010000111011001",
			2160 => "0000000010000111011001",
			2161 => "0011111001110000000100",
			2162 => "0000000010000111011001",
			2163 => "0001111000000000000100",
			2164 => "0000000010000111011001",
			2165 => "0000000010000111011001",
			2166 => "0000101101000100010000",
			2167 => "0001110101011100001000",
			2168 => "0001100011001000000100",
			2169 => "0000000010001000101101",
			2170 => "0000000010001000101101",
			2171 => "0001001001100100000100",
			2172 => "0000000010001000101101",
			2173 => "0000000010001000101101",
			2174 => "0011111111100000001000",
			2175 => "0000111111011000000100",
			2176 => "0000000010001000101101",
			2177 => "0000000010001000101101",
			2178 => "0000100101001100000100",
			2179 => "0000000010001000101101",
			2180 => "0011111001110000000100",
			2181 => "0000000010001000101101",
			2182 => "0011011000000100001000",
			2183 => "0001111100000000000100",
			2184 => "0000000010001000101101",
			2185 => "0000000010001000101101",
			2186 => "0000000010001000101101",
			2187 => "0011110100100100100100",
			2188 => "0000101101000100010000",
			2189 => "0000111100101000001100",
			2190 => "0010011010100100000100",
			2191 => "0000000010001010010001",
			2192 => "0000000001101000000100",
			2193 => "0000000010001010010001",
			2194 => "0000000010001010010001",
			2195 => "0000000010001010010001",
			2196 => "0011111111100000001000",
			2197 => "0000111111011000000100",
			2198 => "0000000010001010010001",
			2199 => "0000000010001010010001",
			2200 => "0000101000110100001000",
			2201 => "0010110101010100000100",
			2202 => "0000000010001010010001",
			2203 => "0000000010001010010001",
			2204 => "0000000010001010010001",
			2205 => "0010111111011000001000",
			2206 => "0010001010100100000100",
			2207 => "0000000010001010010001",
			2208 => "0000000010001010010001",
			2209 => "0010010001010000000100",
			2210 => "0000000010001010010001",
			2211 => "0000000010001010010001",
			2212 => "0011110001010100011100",
			2213 => "0000111111011000010000",
			2214 => "0000100000111000000100",
			2215 => "0000000010001011110101",
			2216 => "0010001001000100000100",
			2217 => "0000000010001011110101",
			2218 => "0010001111001000000100",
			2219 => "0000000010001011110101",
			2220 => "0000000010001011110101",
			2221 => "0010001001000100000100",
			2222 => "0000000010001011110101",
			2223 => "0010001010000100000100",
			2224 => "0000000010001011110101",
			2225 => "0000000010001011110101",
			2226 => "0000101101100100000100",
			2227 => "0000000010001011110101",
			2228 => "0001101001110000010000",
			2229 => "0001011100110100001000",
			2230 => "0001001010100100000100",
			2231 => "0000000010001011110101",
			2232 => "0000000010001011110101",
			2233 => "0000100100111100000100",
			2234 => "0000000010001011110101",
			2235 => "0000000010001011110101",
			2236 => "0000000010001011110101",
			2237 => "0000011001100100010100",
			2238 => "0001001110011000001000",
			2239 => "0010101110011000000100",
			2240 => "0000000010001101101001",
			2241 => "0000000010001101101001",
			2242 => "0011011011101100001000",
			2243 => "0001111000000000000100",
			2244 => "0000000010001101101001",
			2245 => "0000000010001101101001",
			2246 => "0000000010001101101001",
			2247 => "0001011001001000010000",
			2248 => "0000001101000100001000",
			2249 => "0000011001100000000100",
			2250 => "0000000010001101101001",
			2251 => "0000000010001101101001",
			2252 => "0001100001010100000100",
			2253 => "0000000010001101101001",
			2254 => "0000000010001101101001",
			2255 => "0011000101101100001000",
			2256 => "0010001010100100000100",
			2257 => "0000000010001101101001",
			2258 => "0000000010001101101001",
			2259 => "0001111000100000001100",
			2260 => "0001001111100000001000",
			2261 => "0000000100011100000100",
			2262 => "0000000010001101101001",
			2263 => "0000000010001101101001",
			2264 => "0000000010001101101001",
			2265 => "0000000010001101101001",
			2266 => "0001101001110000100000",
			2267 => "0000100000111000000100",
			2268 => "0000000010001110101101",
			2269 => "0001011100011100001000",
			2270 => "0011011101101000000100",
			2271 => "0000000010001110101101",
			2272 => "0000000010001110101101",
			2273 => "0011011100101000001100",
			2274 => "0000011001100100000100",
			2275 => "0000000010001110101101",
			2276 => "0010001001001100000100",
			2277 => "0000000010001110101101",
			2278 => "0000000010001110101101",
			2279 => "0001001101111100000100",
			2280 => "0000000010001110101101",
			2281 => "0000000010001110101101",
			2282 => "0000000010001110101101",
			2283 => "0000101101000100010000",
			2284 => "0001110101011100001000",
			2285 => "0011111000000100000100",
			2286 => "0000000010010000010001",
			2287 => "0000000010010000010001",
			2288 => "0001001001100100000100",
			2289 => "0000000010010000010001",
			2290 => "0000000010010000010001",
			2291 => "0011110110100000011100",
			2292 => "0001010001101000010100",
			2293 => "0001000111110000000100",
			2294 => "0000000010010000010001",
			2295 => "0000101101100000001100",
			2296 => "0000101111110000000100",
			2297 => "0000000010010000010001",
			2298 => "0000101111110100000100",
			2299 => "0000000010010000010001",
			2300 => "0000000010010000010001",
			2301 => "0000000010010000010001",
			2302 => "0011011001001000000100",
			2303 => "0000000010010000010001",
			2304 => "0000000010010000010001",
			2305 => "0011011000000100000100",
			2306 => "0000000010010000010001",
			2307 => "0000000010010000010001",
			2308 => "0001100100100100101100",
			2309 => "0000101101000100010000",
			2310 => "0001101001011000001100",
			2311 => "0000100000111000000100",
			2312 => "1111111010010001111101",
			2313 => "0010100101101100000100",
			2314 => "0000001010010001111101",
			2315 => "0000000010010001111101",
			2316 => "1111111010010001111101",
			2317 => "0011111111100000001000",
			2318 => "0001011001010100000100",
			2319 => "0000001010010001111101",
			2320 => "0000000010010001111101",
			2321 => "0000100101001100001000",
			2322 => "0011110100000000000100",
			2323 => "0000000010010001111101",
			2324 => "1111111010010001111101",
			2325 => "0001010001101000000100",
			2326 => "0000001010010001111101",
			2327 => "0000100010111100000100",
			2328 => "0000000010010001111101",
			2329 => "0000000010010001111101",
			2330 => "0011011000000100000100",
			2331 => "1111111010010001111101",
			2332 => "0011001100010000000100",
			2333 => "0000000010010001111101",
			2334 => "0000000010010001111101",
			2335 => "0001100000010100101100",
			2336 => "0000101101000100010000",
			2337 => "0001110101011100001000",
			2338 => "0011111100000000000100",
			2339 => "0000000010010011011001",
			2340 => "0000000010010011011001",
			2341 => "0001001001100100000100",
			2342 => "0000000010010011011001",
			2343 => "0000000010010011011001",
			2344 => "0001010000111100001100",
			2345 => "0001101001101100000100",
			2346 => "0000000010010011011001",
			2347 => "0000100001000000000100",
			2348 => "0000000010010011011001",
			2349 => "0000000010010011011001",
			2350 => "0000001000001000001100",
			2351 => "0011000111011100001000",
			2352 => "0001001100101100000100",
			2353 => "0000000010010011011001",
			2354 => "0000000010010011011001",
			2355 => "0000000010010011011001",
			2356 => "0000000010010011011001",
			2357 => "0000000010010011011001",
			2358 => "0011110001001100101100",
			2359 => "0000101101000100001100",
			2360 => "0001111100101000001000",
			2361 => "0000011001100100000100",
			2362 => "0000000010010100110101",
			2363 => "0000000010010100110101",
			2364 => "1111111010010100110101",
			2365 => "0011110000100000010100",
			2366 => "0000100001000000001100",
			2367 => "0011111111100000001000",
			2368 => "0000111111011000000100",
			2369 => "0000001010010100110101",
			2370 => "0000000010010100110101",
			2371 => "1111111010010100110101",
			2372 => "0001010001101000000100",
			2373 => "0000001010010100110101",
			2374 => "0000000010010100110101",
			2375 => "0000000101000100000100",
			2376 => "1111111010010100110101",
			2377 => "0001000000100000000100",
			2378 => "0000001010010100110101",
			2379 => "0000000010010100110101",
			2380 => "1111111010010100110101",
			2381 => "0011110001001100101100",
			2382 => "0000101101100000011000",
			2383 => "0010101110011000001000",
			2384 => "0000001010100000000100",
			2385 => "0000000010010110010001",
			2386 => "0000000010010110010001",
			2387 => "0010110110001100000100",
			2388 => "0000000010010110010001",
			2389 => "0001101110111000001000",
			2390 => "0001100011000100000100",
			2391 => "0000000010010110010001",
			2392 => "0000000010010110010001",
			2393 => "0000000010010110010001",
			2394 => "0001001101111100010000",
			2395 => "0000100101001100001100",
			2396 => "0001011011000000001000",
			2397 => "0010111010100100000100",
			2398 => "0000000010010110010001",
			2399 => "0000000010010110010001",
			2400 => "0000000010010110010001",
			2401 => "0000000010010110010001",
			2402 => "0000000010010110010001",
			2403 => "0000000010010110010001",
			2404 => "0001100100100100110100",
			2405 => "0000101101000100010100",
			2406 => "0001111100101000001000",
			2407 => "0000001100110100000100",
			2408 => "0000000010011000001101",
			2409 => "0000001010011000001101",
			2410 => "0001101001011000001000",
			2411 => "0011111011111000000100",
			2412 => "0000000010011000001101",
			2413 => "0000000010011000001101",
			2414 => "1111111010011000001101",
			2415 => "0011111111100000001000",
			2416 => "0001011001010100000100",
			2417 => "0000001010011000001101",
			2418 => "0000000010011000001101",
			2419 => "0000100101001100001000",
			2420 => "0001000101010100000100",
			2421 => "0000000010011000001101",
			2422 => "1111111010011000001101",
			2423 => "0001010001101000001000",
			2424 => "0001101011110000000100",
			2425 => "0000001010011000001101",
			2426 => "0000000010011000001101",
			2427 => "0000100010111100000100",
			2428 => "0000000010011000001101",
			2429 => "0000000010011000001101",
			2430 => "0011011000000100000100",
			2431 => "1111111010011000001101",
			2432 => "0011001100010000000100",
			2433 => "0000000010011000001101",
			2434 => "0000000010011000001101",
			2435 => "0001101001110000110000",
			2436 => "0000101101000100010000",
			2437 => "0001101001011000001100",
			2438 => "0000100000111000000100",
			2439 => "0000000010011001110001",
			2440 => "0010100101101100000100",
			2441 => "0000000010011001110001",
			2442 => "0000000010011001110001",
			2443 => "0000000010011001110001",
			2444 => "0001011100011100001100",
			2445 => "0001101001101100000100",
			2446 => "0000000010011001110001",
			2447 => "0000100001000000000100",
			2448 => "0000000010011001110001",
			2449 => "0000000010011001110001",
			2450 => "0000001000001000001100",
			2451 => "0010000101011100001000",
			2452 => "0011011011101100000100",
			2453 => "0000000010011001110001",
			2454 => "0000000010011001110001",
			2455 => "0000000010011001110001",
			2456 => "0001000000100000000100",
			2457 => "0000000010011001110001",
			2458 => "0000000010011001110001",
			2459 => "0000000010011001110001",
			2460 => "0011110100100100100100",
			2461 => "0000101110010000011100",
			2462 => "0001101001000000010000",
			2463 => "0000100000111000000100",
			2464 => "0000000010011011110101",
			2465 => "0010000101011100000100",
			2466 => "0000001010011011110101",
			2467 => "0000110111011100000100",
			2468 => "0000000010011011110101",
			2469 => "0000000010011011110101",
			2470 => "0000000111001000000100",
			2471 => "1111111010011011110101",
			2472 => "0011111010100000000100",
			2473 => "0000000010011011110101",
			2474 => "0000000010011011110101",
			2475 => "0001010001101000000100",
			2476 => "0000001010011011110101",
			2477 => "0000000010011011110101",
			2478 => "0010001010100100000100",
			2479 => "0000000010011011110101",
			2480 => "0010111111011000010100",
			2481 => "0011001111011000001100",
			2482 => "0010000011010000001000",
			2483 => "0011001110011000000100",
			2484 => "0000000010011011110101",
			2485 => "0000000010011011110101",
			2486 => "1111111010011011110101",
			2487 => "0010011101001000000100",
			2488 => "0000000010011011110101",
			2489 => "0000000010011011110101",
			2490 => "0001110000111100000100",
			2491 => "0000000010011011110101",
			2492 => "0000000010011011110101",
			2493 => "0011110001001100110000",
			2494 => "0000101101000100010000",
			2495 => "0001101001011000001100",
			2496 => "0000100000111000000100",
			2497 => "0000000010011101011001",
			2498 => "0010100101101100000100",
			2499 => "0000000010011101011001",
			2500 => "0000000010011101011001",
			2501 => "0000000010011101011001",
			2502 => "0011111111100000001000",
			2503 => "0001011001010100000100",
			2504 => "0000001010011101011001",
			2505 => "0000000010011101011001",
			2506 => "0000100101001100001000",
			2507 => "0001000101010100000100",
			2508 => "0000000010011101011001",
			2509 => "0000000010011101011001",
			2510 => "0001010001101000001000",
			2511 => "0011110100100100000100",
			2512 => "0000001010011101011001",
			2513 => "0000000010011101011001",
			2514 => "0000100100111100000100",
			2515 => "0000000010011101011001",
			2516 => "0000000010011101011001",
			2517 => "0000000010011101011001",
			2518 => "0011110001001100110100",
			2519 => "0000101101000100010000",
			2520 => "0001101001011000001100",
			2521 => "0010000011010000000100",
			2522 => "0000000010011111000101",
			2523 => "0001000001110000000100",
			2524 => "0000000010011111000101",
			2525 => "0000000010011111000101",
			2526 => "0000000010011111000101",
			2527 => "0001011110111000010000",
			2528 => "0000101101100000001000",
			2529 => "0001100001101000000100",
			2530 => "0000000010011111000101",
			2531 => "0000000010011111000101",
			2532 => "0001000001100100000100",
			2533 => "0000000010011111000101",
			2534 => "0000000010011111000101",
			2535 => "0000001000001000001100",
			2536 => "0011000111011100001000",
			2537 => "0001001100101100000100",
			2538 => "0000000010011111000101",
			2539 => "0000000010011111000101",
			2540 => "0000000010011111000101",
			2541 => "0001000000100000000100",
			2542 => "0000000010011111000101",
			2543 => "0000000010011111000101",
			2544 => "0000000010011111000101",
			2545 => "0011110001001100110100",
			2546 => "0000101101000100001100",
			2547 => "0010000011010000000100",
			2548 => "0000000010100000110001",
			2549 => "0001000001110000000100",
			2550 => "0000000010100000110001",
			2551 => "1111111010100000110001",
			2552 => "0001010100101100010100",
			2553 => "0001101101111100001100",
			2554 => "0000010110010000000100",
			2555 => "0000001010100000110001",
			2556 => "0000001111010100000100",
			2557 => "0000000010100000110001",
			2558 => "0000001010100000110001",
			2559 => "0000000101100000000100",
			2560 => "1111111010100000110001",
			2561 => "0000001010100000110001",
			2562 => "0000100000100100001100",
			2563 => "0011111101101100001000",
			2564 => "0000001101100100000100",
			2565 => "0000000010100000110001",
			2566 => "0000000010100000110001",
			2567 => "1111111010100000110001",
			2568 => "0001000000100000000100",
			2569 => "0000001010100000110001",
			2570 => "0000000010100000110001",
			2571 => "1111111010100000110001",
			2572 => "0011110110100000101100",
			2573 => "0000101000010100100100",
			2574 => "0011110100000000100000",
			2575 => "0000101101000100010000",
			2576 => "0001101001011000001100",
			2577 => "0010011001001000001000",
			2578 => "0000001110010100000100",
			2579 => "0000000010100010011101",
			2580 => "0000000010100010011101",
			2581 => "0000000010100010011101",
			2582 => "1111111010100010011101",
			2583 => "0001011001010100001000",
			2584 => "0001011111011000000100",
			2585 => "0000001010100010011101",
			2586 => "0000000010100010011101",
			2587 => "0000001110100100000100",
			2588 => "0000000010100010011101",
			2589 => "0000000010100010011101",
			2590 => "0000000010100010011101",
			2591 => "0001000100100100000100",
			2592 => "0000001010100010011101",
			2593 => "0000000010100010011101",
			2594 => "0011011000000100000100",
			2595 => "1111111010100010011101",
			2596 => "0001001001010000000100",
			2597 => "0000000010100010011101",
			2598 => "0000000010100010011101",
			2599 => "0011110110100000110100",
			2600 => "0000000110100000010000",
			2601 => "0011011101000000000100",
			2602 => "0000000010100100010001",
			2603 => "0001110101011100001000",
			2604 => "0001100011000000000100",
			2605 => "0000000010100100010001",
			2606 => "0000000010100100010001",
			2607 => "0000000010100100010001",
			2608 => "0011111111100000001000",
			2609 => "0001011001010100000100",
			2610 => "0000000010100100010001",
			2611 => "0000000010100100010001",
			2612 => "0000101000010100001100",
			2613 => "0011110100000000001000",
			2614 => "0000000010110100000100",
			2615 => "0000000010100100010001",
			2616 => "0000000010100100010001",
			2617 => "0000000010100100010001",
			2618 => "0001000100100100001100",
			2619 => "0000100010111100001000",
			2620 => "0000000000000100000100",
			2621 => "0000000010100100010001",
			2622 => "0000000010100100010001",
			2623 => "0000000010100100010001",
			2624 => "0000000010100100010001",
			2625 => "0011011000000100000100",
			2626 => "0000000010100100010001",
			2627 => "0000000010100100010001",
			2628 => "0011110001001100110100",
			2629 => "0000000110100000001100",
			2630 => "0010000011010000000100",
			2631 => "0000000010100101111101",
			2632 => "0001000001110000000100",
			2633 => "0000000010100101111101",
			2634 => "0000000010100101111101",
			2635 => "0001011100110100011000",
			2636 => "0011110100100100010000",
			2637 => "0000010110010000000100",
			2638 => "0000000010100101111101",
			2639 => "0000000010110100001000",
			2640 => "0001010101010100000100",
			2641 => "0000000010100101111101",
			2642 => "0000000010100101111101",
			2643 => "0000000010100101111101",
			2644 => "0001101111111000000100",
			2645 => "0000000010100101111101",
			2646 => "0000000010100101111101",
			2647 => "0000100100111100001000",
			2648 => "0010001001001100000100",
			2649 => "0000000010100101111101",
			2650 => "0000000010100101111101",
			2651 => "0000011101000000000100",
			2652 => "0000000010100101111101",
			2653 => "0000000010100101111101",
			2654 => "0000000010100101111101",
			2655 => "0001101001110000110000",
			2656 => "0000100111010000101000",
			2657 => "0011110100000000011100",
			2658 => "0000000000110100010000",
			2659 => "0011110001011000001100",
			2660 => "0000100000111000000100",
			2661 => "0000000010100111100001",
			2662 => "0010011001001000000100",
			2663 => "0000000010100111100001",
			2664 => "0000000010100111100001",
			2665 => "0000000010100111100001",
			2666 => "0000111001010100001000",
			2667 => "0010001010000100000100",
			2668 => "0000000010100111100001",
			2669 => "0000000010100111100001",
			2670 => "0000000010100111100001",
			2671 => "0000101000010100000100",
			2672 => "0000000010100111100001",
			2673 => "0011011011101100000100",
			2674 => "0000000010100111100001",
			2675 => "0000000010100111100001",
			2676 => "0001000000100000000100",
			2677 => "0000000010100111100001",
			2678 => "0000000010100111100001",
			2679 => "0000000010100111100001",
			2680 => "0011110001001100110100",
			2681 => "0000101101000100001100",
			2682 => "0010000011010000000100",
			2683 => "0000000010101001001101",
			2684 => "0001001001100100000100",
			2685 => "0000000010101001001101",
			2686 => "0000000010101001001101",
			2687 => "0001000101111000001100",
			2688 => "0001101010100000000100",
			2689 => "0000000010101001001101",
			2690 => "0000101011011100000100",
			2691 => "0000000010101001001101",
			2692 => "0000000010101001001101",
			2693 => "0000101000010100001100",
			2694 => "0001000001011000000100",
			2695 => "0000000010101001001101",
			2696 => "0000100101100000000100",
			2697 => "0000000010101001001101",
			2698 => "0000000010101001001101",
			2699 => "0001000000100000001100",
			2700 => "0000001000001000001000",
			2701 => "0011110010010100000100",
			2702 => "0000000010101001001101",
			2703 => "0000000010101001001101",
			2704 => "0000000010101001001101",
			2705 => "0000000010101001001101",
			2706 => "0000000010101001001101",
			2707 => "0001101001110000110100",
			2708 => "0000101101000100010000",
			2709 => "0000111100101000001100",
			2710 => "0010011010100100000100",
			2711 => "0000000010101010111001",
			2712 => "0000101100110100000100",
			2713 => "0000000010101010111001",
			2714 => "0000000010101010111001",
			2715 => "0000000010101010111001",
			2716 => "0011111111100000001000",
			2717 => "0000111111011000000100",
			2718 => "0000000010101010111001",
			2719 => "0000000010101010111001",
			2720 => "0000100101100000001000",
			2721 => "0001000101010100000100",
			2722 => "0000000010101010111001",
			2723 => "0000000010101010111001",
			2724 => "0001001101111100010000",
			2725 => "0000101000010100001000",
			2726 => "0001101011110000000100",
			2727 => "0000000010101010111001",
			2728 => "0000000010101010111001",
			2729 => "0001100000010100000100",
			2730 => "0000000010101010111001",
			2731 => "0000000010101010111001",
			2732 => "0000000010101010111001",
			2733 => "0000000010101010111001",
			2734 => "0011110001001100111000",
			2735 => "0000000000110100010000",
			2736 => "0011110001011000001100",
			2737 => "0000100000111000000100",
			2738 => "0000000010101100101101",
			2739 => "0010011001001000000100",
			2740 => "0000000010101100101101",
			2741 => "0000000010101100101101",
			2742 => "0000000010101100101101",
			2743 => "0001100001111100001100",
			2744 => "0001011001010100001000",
			2745 => "0010001010000100000100",
			2746 => "0000001010101100101101",
			2747 => "0000000010101100101101",
			2748 => "0000000010101100101101",
			2749 => "0000101000010100001100",
			2750 => "0011111101101100001000",
			2751 => "0000100100010000000100",
			2752 => "0000000010101100101101",
			2753 => "0000000010101100101101",
			2754 => "0000000010101100101101",
			2755 => "0001000000100000001100",
			2756 => "0000100101111100001000",
			2757 => "0011110100100100000100",
			2758 => "0000000010101100101101",
			2759 => "0000000010101100101101",
			2760 => "0000000010101100101101",
			2761 => "0000000010101100101101",
			2762 => "0000000010101100101101",
			2763 => "0001101001110000110000",
			2764 => "0000100000111000000100",
			2765 => "0000000010101110010001",
			2766 => "0001011000101000010100",
			2767 => "0001101001101100001100",
			2768 => "0000000110100000001000",
			2769 => "0010111010100100000100",
			2770 => "0000000010101110010001",
			2771 => "0000000010101110010001",
			2772 => "0000000010101110010001",
			2773 => "0000001010001000000100",
			2774 => "0000000010101110010001",
			2775 => "0000000010101110010001",
			2776 => "0000001000001000010000",
			2777 => "0010000101011100001100",
			2778 => "0000000000010000000100",
			2779 => "0000000010101110010001",
			2780 => "0000010000011000000100",
			2781 => "0000000010101110010001",
			2782 => "0000000010101110010001",
			2783 => "0000000010101110010001",
			2784 => "0001000000100000000100",
			2785 => "0000000010101110010001",
			2786 => "0000000010101110010001",
			2787 => "0000000010101110010001",
			2788 => "0001100101001000111100",
			2789 => "0000101111100000001000",
			2790 => "0000011000111100000100",
			2791 => "0000000010110000011101",
			2792 => "1111111010110000011101",
			2793 => "0001010011110100100100",
			2794 => "0000101101100100010000",
			2795 => "0001011001001000001000",
			2796 => "0001101110111000000100",
			2797 => "0000010010110000011101",
			2798 => "0000001010110000011101",
			2799 => "0000010001110000000100",
			2800 => "0000001010110000011101",
			2801 => "1111111010110000011101",
			2802 => "0011111111100100001000",
			2803 => "0000100100000100000100",
			2804 => "0000010010110000011101",
			2805 => "0000010010110000011101",
			2806 => "0000000111000000000100",
			2807 => "1111111010110000011101",
			2808 => "0011111111111000000100",
			2809 => "0000010010110000011101",
			2810 => "0000010010110000011101",
			2811 => "0000001000001000001100",
			2812 => "0000010000011000001000",
			2813 => "0001101010110100000100",
			2814 => "0000000010110000011101",
			2815 => "1111111010110000011101",
			2816 => "1111111010110000011101",
			2817 => "0000010010110000011101",
			2818 => "0011011000000100000100",
			2819 => "1111111010110000011101",
			2820 => "0010011011111000000100",
			2821 => "0000000010110000011101",
			2822 => "1111111010110000011101",
			2823 => "0011110001001100111000",
			2824 => "0000100111010000110000",
			2825 => "0001010011000000011100",
			2826 => "0000100110100000010100",
			2827 => "0001110101011100001000",
			2828 => "0000100011000100000100",
			2829 => "0000000010110010010001",
			2830 => "0000000010110010010001",
			2831 => "0010101110011000001000",
			2832 => "0001011110011000000100",
			2833 => "0000000010110010010001",
			2834 => "0000000010110010010001",
			2835 => "0000000010110010010001",
			2836 => "0001101001101100000100",
			2837 => "0000000010110010010001",
			2838 => "0000000010110010010001",
			2839 => "0000010111110000001100",
			2840 => "0011110000100000001000",
			2841 => "0000001101100100000100",
			2842 => "0000000010110010010001",
			2843 => "0000000010110010010001",
			2844 => "0000000010110010010001",
			2845 => "0000101110000100000100",
			2846 => "0000000010110010010001",
			2847 => "0000000010110010010001",
			2848 => "0001000000100000000100",
			2849 => "0000000010110010010001",
			2850 => "0000000010110010010001",
			2851 => "0000000010110010010001",
			2852 => "0001101001110001000000",
			2853 => "0000101100100000010100",
			2854 => "0011110011110100010000",
			2855 => "0010000101011100001000",
			2856 => "0000100000111000000100",
			2857 => "0000000010110100010101",
			2858 => "0000000010110100010101",
			2859 => "0000101101101100000100",
			2860 => "0000000010110100010101",
			2861 => "0000000010110100010101",
			2862 => "0000000010110100010101",
			2863 => "0001001111011000010000",
			2864 => "0011110111010100000100",
			2865 => "0000000010110100010101",
			2866 => "0010110101010100001000",
			2867 => "0010111110011000000100",
			2868 => "0000000010110100010101",
			2869 => "0000000010110100010101",
			2870 => "0000000010110100010101",
			2871 => "0000101000010100001100",
			2872 => "0001000001011000000100",
			2873 => "0000000010110100010101",
			2874 => "0000100101100000000100",
			2875 => "0000000010110100010101",
			2876 => "0000000010110100010101",
			2877 => "0001000000100000001100",
			2878 => "0000001000001000001000",
			2879 => "0011110010010100000100",
			2880 => "0000000010110100010101",
			2881 => "0000000010110100010101",
			2882 => "0000000010110100010101",
			2883 => "0000000010110100010101",
			2884 => "0000000010110100010101",
			2885 => "0011110001001100110100",
			2886 => "0000100000111000000100",
			2887 => "1111111010110110000001",
			2888 => "0001010100101100011100",
			2889 => "0001101001101100010000",
			2890 => "0000101100100000001100",
			2891 => "0000111100101000000100",
			2892 => "0000001010110110000001",
			2893 => "0001011101001000000100",
			2894 => "1111111010110110000001",
			2895 => "0000000010110110000001",
			2896 => "0000001010110110000001",
			2897 => "0000100001000000000100",
			2898 => "1111111010110110000001",
			2899 => "0000010000011000000100",
			2900 => "0000000010110110000001",
			2901 => "0000001010110110000001",
			2902 => "0000001000001000001100",
			2903 => "0011101010100000001000",
			2904 => "0000001100000100000100",
			2905 => "1111111010110110000001",
			2906 => "0000001010110110000001",
			2907 => "1111111010110110000001",
			2908 => "0001000000100000000100",
			2909 => "0000001010110110000001",
			2910 => "1111111010110110000001",
			2911 => "1111111010110110000001",
			2912 => "0001100000010101000000",
			2913 => "0000101111100000001000",
			2914 => "0000011000111100000100",
			2915 => "0000000010111000010101",
			2916 => "1111111010111000010101",
			2917 => "0001011110111000101000",
			2918 => "0000101101100000010000",
			2919 => "0000110111011100001000",
			2920 => "0000010001110000000100",
			2921 => "0000010010111000010101",
			2922 => "0000010010111000010101",
			2923 => "0010001111111100000100",
			2924 => "0000000010111000010101",
			2925 => "1111111010111000010101",
			2926 => "0011110101110000001100",
			2927 => "0000001000110100001000",
			2928 => "0001000110001100000100",
			2929 => "0000010010111000010101",
			2930 => "0000011010111000010101",
			2931 => "0000010010111000010101",
			2932 => "0000000000000100000100",
			2933 => "1111111010111000010101",
			2934 => "0010111010100100000100",
			2935 => "0000010010111000010101",
			2936 => "0000010010111000010101",
			2937 => "0000100000100100001100",
			2938 => "0000011000111100000100",
			2939 => "0000000010111000010101",
			2940 => "0011110101110000000100",
			2941 => "0000000010111000010101",
			2942 => "1111111010111000010101",
			2943 => "0000010010111000010101",
			2944 => "0011011000000100000100",
			2945 => "1111111010111000010101",
			2946 => "0011011000000000000100",
			2947 => "0000000010111000010101",
			2948 => "1111111010111000010101",
			2949 => "0011110001001100110000",
			2950 => "0000101111100000000100",
			2951 => "1111111010111001111001",
			2952 => "0001010001101000100100",
			2953 => "0000101101100000001100",
			2954 => "0001010011000000001000",
			2955 => "0010101010100100000100",
			2956 => "0000001010111001111001",
			2957 => "0000000010111001111001",
			2958 => "1111111010111001111001",
			2959 => "0011110100000000001000",
			2960 => "0001111100000000000100",
			2961 => "0000001010111001111001",
			2962 => "0000001010111001111001",
			2963 => "0000001101010000001000",
			2964 => "0001101010100000000100",
			2965 => "0000000010111001111001",
			2966 => "1111111010111001111001",
			2967 => "0000100111010000000100",
			2968 => "0000001010111001111001",
			2969 => "0000001010111001111001",
			2970 => "0000010110110100000100",
			2971 => "1111111010111001111001",
			2972 => "0000001010111001111001",
			2973 => "1111111010111001111001",
			2974 => "0011110001001101000000",
			2975 => "0000011001100100010000",
			2976 => "0000110001001000001100",
			2977 => "0001001110011000001000",
			2978 => "0001110011000000000100",
			2979 => "0000000010111011111101",
			2980 => "0000000010111011111101",
			2981 => "0000001010111011111101",
			2982 => "0000000010111011111101",
			2983 => "0000001101100100010100",
			2984 => "0001011001001000010000",
			2985 => "0010001001001100000100",
			2986 => "0000000010111011111101",
			2987 => "0011001110011000000100",
			2988 => "0000000010111011111101",
			2989 => "0010011010000100000100",
			2990 => "0000000010111011111101",
			2991 => "0000000010111011111101",
			2992 => "1111111010111011111101",
			2993 => "0001010100101100001000",
			2994 => "0010111010100100000100",
			2995 => "0000000010111011111101",
			2996 => "0000001010111011111101",
			2997 => "0000000101000100001100",
			2998 => "0010001001001100000100",
			2999 => "0000000010111011111101",
			3000 => "0011011100101000000100",
			3001 => "1111111010111011111101",
			3002 => "0000000010111011111101",
			3003 => "0001000000100000000100",
			3004 => "0000000010111011111101",
			3005 => "0000000010111011111101",
			3006 => "1111111010111011111101",
			3007 => "0011110001001100101000",
			3008 => "0000101111100000000100",
			3009 => "1111111010111101010001",
			3010 => "0010101010100100000100",
			3011 => "0000001010111101010001",
			3012 => "0000100110100000000100",
			3013 => "1111111010111101010001",
			3014 => "0001100001111100001100",
			3015 => "0001011001010100001000",
			3016 => "0000011001100000000100",
			3017 => "0000001010111101010001",
			3018 => "0000001010111101010001",
			3019 => "0000000010111101010001",
			3020 => "0000100101001100001000",
			3021 => "0011110101110000000100",
			3022 => "0000000010111101010001",
			3023 => "1111111010111101010001",
			3024 => "0001001101111100000100",
			3025 => "0000001010111101010001",
			3026 => "1111111010111101010001",
			3027 => "1111111010111101010001",
			3028 => "0001100000010101000000",
			3029 => "0000101111100000001000",
			3030 => "0001011010000100000100",
			3031 => "1111111010111111100101",
			3032 => "0000000010111111100101",
			3033 => "0001010001101000110000",
			3034 => "0000101110010000011100",
			3035 => "0001010011000000001100",
			3036 => "0001100010001100001000",
			3037 => "0000001110111100000100",
			3038 => "0000001010111111100101",
			3039 => "0000001010111111100101",
			3040 => "0000000010111111100101",
			3041 => "0010011010000100001000",
			3042 => "0011111100011100000100",
			3043 => "0000000010111111100101",
			3044 => "1111111010111111100101",
			3045 => "0001001000000000000100",
			3046 => "0000001010111111100101",
			3047 => "1111111010111111100101",
			3048 => "0000100101001100001000",
			3049 => "0001101111100000000100",
			3050 => "0000001010111111100101",
			3051 => "0000000010111111100101",
			3052 => "0011011011101100000100",
			3053 => "0000001010111111100101",
			3054 => "0000100100001000000100",
			3055 => "0000001010111111100101",
			3056 => "0000001010111111100101",
			3057 => "0000011101000000000100",
			3058 => "1111111010111111100101",
			3059 => "0000001010111111100101",
			3060 => "0011011000000100000100",
			3061 => "1111111010111111100101",
			3062 => "0011011000000000000100",
			3063 => "0000000010111111100101",
			3064 => "1111111010111111100101",
			3065 => "0011110001001100110000",
			3066 => "0000100111010000101000",
			3067 => "0011110000100000100100",
			3068 => "0000101000101100100000",
			3069 => "0011111010011100010000",
			3070 => "0000010001110000001000",
			3071 => "0000001110010100000100",
			3072 => "0000000011000001001001",
			3073 => "0000001011000001001001",
			3074 => "0001010011010000000100",
			3075 => "0000000011000001001001",
			3076 => "1111111011000001001001",
			3077 => "0000000111001000001000",
			3078 => "0000010011110000000100",
			3079 => "1111111011000001001001",
			3080 => "0000000011000001001001",
			3081 => "0001000101111000000100",
			3082 => "0000000011000001001001",
			3083 => "1111111011000001001001",
			3084 => "0000001011000001001001",
			3085 => "1111111011000001001001",
			3086 => "0000111001111100000100",
			3087 => "0000001011000001001001",
			3088 => "0000000011000001001001",
			3089 => "1111111011000001001001",
			3090 => "0011110001001100111100",
			3091 => "0010001010100100000100",
			3092 => "0000000011000011000101",
			3093 => "0000000110100000010000",
			3094 => "0000111001100000001000",
			3095 => "0001010001100100000100",
			3096 => "0000000011000011000101",
			3097 => "0000000011000011000101",
			3098 => "0010001001001100000100",
			3099 => "0000000011000011000101",
			3100 => "0000000011000011000101",
			3101 => "0001000101111000010100",
			3102 => "0010111110011000000100",
			3103 => "0000000011000011000101",
			3104 => "0001101010100000001000",
			3105 => "0000011111011100000100",
			3106 => "0000000011000011000101",
			3107 => "0000000011000011000101",
			3108 => "0011010011010000000100",
			3109 => "0000000011000011000101",
			3110 => "0000000011000011000101",
			3111 => "0000100101001100001000",
			3112 => "0000111001010100000100",
			3113 => "0000000011000011000101",
			3114 => "0000000011000011000101",
			3115 => "0011110100100100000100",
			3116 => "0000000011000011000101",
			3117 => "0000101011011000000100",
			3118 => "0000000011000011000101",
			3119 => "0000000011000011000101",
			3120 => "0000000011000011000101",
			3121 => "0011110001001100110100",
			3122 => "0000100000111000000100",
			3123 => "1111111011000100110001",
			3124 => "0011010011110000000100",
			3125 => "0000001011000100110001",
			3126 => "0000101101000100010000",
			3127 => "0001101011111000001000",
			3128 => "0001000110001100000100",
			3129 => "0000000011000100110001",
			3130 => "1111111011000100110001",
			3131 => "0011001010100100000100",
			3132 => "1111111011000100110001",
			3133 => "1111111011000100110001",
			3134 => "0001100001111100001100",
			3135 => "0001011001010100001000",
			3136 => "0000010110010000000100",
			3137 => "0000001011000100110001",
			3138 => "0000001011000100110001",
			3139 => "0000000011000100110001",
			3140 => "0000100101100000001000",
			3141 => "0001000101010100000100",
			3142 => "0000000011000100110001",
			3143 => "1111111011000100110001",
			3144 => "0011110100100100000100",
			3145 => "0000001011000100110001",
			3146 => "0000000011000100110001",
			3147 => "1111111011000100110001",
			3148 => "0011110001001100110100",
			3149 => "0000100000111000000100",
			3150 => "1111111011000110011111",
			3151 => "0010101010011000101100",
			3152 => "0000100111010000100000",
			3153 => "0011110100000000010000",
			3154 => "0000101100100000001000",
			3155 => "0010001001001100000100",
			3156 => "0000001011000110011111",
			3157 => "0000000011000110011111",
			3158 => "0001001000000100000100",
			3159 => "0000001011000110011111",
			3160 => "0000000011000110011111",
			3161 => "0000101000010100001000",
			3162 => "0011111101101100000100",
			3163 => "0000000011000110011111",
			3164 => "1111111011000110011111",
			3165 => "0010101001000000000100",
			3166 => "0000001011000110011111",
			3167 => "1111111011000110011111",
			3168 => "0000000111101100001000",
			3169 => "0011101001111100000100",
			3170 => "0000001011000110011111",
			3171 => "0000000011000110011111",
			3172 => "0000001011000110011111",
			3173 => "1111111011000110011111",
			3174 => "1111111011000110011111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1063, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2143, initial_addr_3'length));
	end generate gen_rom_9;

	gen_rom_10: if SELECT_ROM = 10 generate
		bank <= (
			0 => "0010111101101000000100",
			1 => "0000000000000000011101",
			2 => "0001001010000100000100",
			3 => "0000000000000000011101",
			4 => "0011110011101000000100",
			5 => "0000000000000000011101",
			6 => "0000000000000000011101",
			7 => "0010101001111100001100",
			8 => "0011001000000100000100",
			9 => "0000000000000001000001",
			10 => "0010101100001100000100",
			11 => "0000000000000001000001",
			12 => "0000000000000001000001",
			13 => "0001000000100000000100",
			14 => "0000000000000001000001",
			15 => "0000000000000001000001",
			16 => "0000110000100000010000",
			17 => "0011110001101000001000",
			18 => "0010101001010100000100",
			19 => "0000000000000001100101",
			20 => "0000000000000001100101",
			21 => "0011001100110000000100",
			22 => "1111111000000001100101",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0011001101101000000100",
			26 => "0000000000000010001001",
			27 => "0000100011111100001000",
			28 => "0001001010000100000100",
			29 => "0000000000000010001001",
			30 => "0000000000000010001001",
			31 => "0000110000100000000100",
			32 => "0000000000000010001001",
			33 => "0000000000000010001001",
			34 => "0011001101101000000100",
			35 => "0000000000000010101101",
			36 => "0000100011111100001000",
			37 => "0000111011000000000100",
			38 => "0000000000000010101101",
			39 => "0000000000000010101101",
			40 => "0000110000100000000100",
			41 => "0000000000000010101101",
			42 => "0000000000000010101101",
			43 => "0000110000100000010000",
			44 => "0011110001101000001000",
			45 => "0010101000101000000100",
			46 => "0000000000000011010001",
			47 => "0000000000000011010001",
			48 => "0011001100110000000100",
			49 => "0000000000000011010001",
			50 => "0000000000000011010001",
			51 => "0000000000000011010001",
			52 => "0010101001111100010000",
			53 => "0011111010011100001000",
			54 => "0000111101001000000100",
			55 => "0000000000000011110101",
			56 => "0000000000000011110101",
			57 => "0011001100110000000100",
			58 => "0000000000000011110101",
			59 => "0000000000000011110101",
			60 => "0000000000000011110101",
			61 => "0000110011110100000100",
			62 => "0000000000000100011001",
			63 => "0000100011111100001000",
			64 => "0010111001000100000100",
			65 => "0000000000000100011001",
			66 => "0000000000000100011001",
			67 => "0000110000100000000100",
			68 => "0000000000000100011001",
			69 => "0000000000000100011001",
			70 => "0000111011000000000100",
			71 => "0000000000000100111101",
			72 => "0000100011111100001000",
			73 => "0010111001000100000100",
			74 => "0000000000000100111101",
			75 => "0000000000000100111101",
			76 => "0000110000100000000100",
			77 => "0000000000000100111101",
			78 => "0000000000000100111101",
			79 => "0001010011101100010000",
			80 => "0011111010011100001000",
			81 => "0001001010000100000100",
			82 => "0000000000000101100001",
			83 => "0000000000000101100001",
			84 => "0011001100110000000100",
			85 => "0000000000000101100001",
			86 => "0000000000000101100001",
			87 => "0000000000000101100001",
			88 => "0010101001111100010000",
			89 => "0011110001101000001000",
			90 => "0010101000101000000100",
			91 => "0000000000000110001101",
			92 => "0000000000000110001101",
			93 => "0011001100110000000100",
			94 => "1111111000000110001101",
			95 => "0000000000000110001101",
			96 => "0011010101111000000100",
			97 => "0000001000000110001101",
			98 => "0000000000000110001101",
			99 => "0010101001111100010000",
			100 => "0000100000010100001000",
			101 => "0010101101001000000100",
			102 => "0000000000000110111001",
			103 => "0000000000000110111001",
			104 => "0011001100110000000100",
			105 => "0000000000000110111001",
			106 => "0000000000000110111001",
			107 => "0001000000100000000100",
			108 => "0000000000000110111001",
			109 => "0000000000000110111001",
			110 => "0010101001111100010000",
			111 => "0011001000000100000100",
			112 => "1111111000000111011101",
			113 => "0000000110001000001000",
			114 => "0001001100101000000100",
			115 => "0000000000000111011101",
			116 => "0000000000000111011101",
			117 => "1111111000000111011101",
			118 => "0000001000000111011101",
			119 => "0010101001111100010000",
			120 => "0010111010000100000100",
			121 => "1111111000001000000001",
			122 => "0000000100110100001000",
			123 => "0010101000101000000100",
			124 => "0000000000001000000001",
			125 => "0000000000001000000001",
			126 => "0000000000001000000001",
			127 => "0000000000001000000001",
			128 => "0000111011000000000100",
			129 => "0000000000001000100101",
			130 => "0011001101101000000100",
			131 => "0000000000001000100101",
			132 => "0000100011111100000100",
			133 => "0000000000001000100101",
			134 => "0000110000100000000100",
			135 => "0000000000001000100101",
			136 => "0000000000001000100101",
			137 => "0000111011000000000100",
			138 => "0000000000001001001001",
			139 => "0011001101101000000100",
			140 => "0000000000001001001001",
			141 => "0000101011001000000100",
			142 => "0000000000001001001001",
			143 => "0000011110011000000100",
			144 => "0000000000001001001001",
			145 => "0000000000001001001001",
			146 => "0000111011000000000100",
			147 => "0000000000001001101101",
			148 => "0011001101101000000100",
			149 => "0000000000001001101101",
			150 => "0000101011001000000100",
			151 => "0000000000001001101101",
			152 => "0000011110011000000100",
			153 => "0000000000001001101101",
			154 => "0000000000001001101101",
			155 => "0010101001111100010000",
			156 => "0010111010000100000100",
			157 => "1111111000001010011001",
			158 => "0000111011000000000100",
			159 => "1111111000001010011001",
			160 => "0000101110011100000100",
			161 => "0000001000001010011001",
			162 => "1111111000001010011001",
			163 => "0000101011001000000100",
			164 => "0000001000001010011001",
			165 => "0000000000001010011001",
			166 => "0010111101101000001000",
			167 => "0001001111100000000100",
			168 => "1111111000001011000101",
			169 => "0000000000001011000101",
			170 => "0000111011000000000100",
			171 => "0000000000001011000101",
			172 => "0000100111111100000100",
			173 => "0000001000001011000101",
			174 => "0000110000100000000100",
			175 => "0000000000001011000101",
			176 => "0000000000001011000101",
			177 => "0010111101101000001000",
			178 => "0011000101111000000100",
			179 => "0000000000001011110001",
			180 => "0000000000001011110001",
			181 => "0001001010000100000100",
			182 => "0000000000001011110001",
			183 => "0000101011001000000100",
			184 => "0000000000001011110001",
			185 => "0000110110100000000100",
			186 => "0000000000001011110001",
			187 => "0000000000001011110001",
			188 => "0010100001101000001100",
			189 => "0000110011110100000100",
			190 => "0000000000001100100101",
			191 => "0010100000111000000100",
			192 => "0000000000001100100101",
			193 => "0000000000001100100101",
			194 => "0000100011111100001000",
			195 => "0010111001000100000100",
			196 => "0000000000001100100101",
			197 => "0000000000001100100101",
			198 => "0000110000100000000100",
			199 => "0000000000001100100101",
			200 => "0000000000001100100101",
			201 => "0001010011101100010100",
			202 => "0011110001101000001000",
			203 => "0010101000101000000100",
			204 => "0000000000001101010001",
			205 => "0000000000001101010001",
			206 => "0011001100110000000100",
			207 => "0000000000001101010001",
			208 => "0010100001101000000100",
			209 => "0000000000001101010001",
			210 => "0000000000001101010001",
			211 => "0000000000001101010001",
			212 => "0000111111100000010100",
			213 => "0010110011001000001100",
			214 => "0010111010000100000100",
			215 => "1111111000001110000101",
			216 => "0010110011000000000100",
			217 => "1111111000001110000101",
			218 => "1111111000001110000101",
			219 => "0000111011000000000100",
			220 => "1111111000001110000101",
			221 => "0000001000001110000101",
			222 => "0000110000100000000100",
			223 => "0000001000001110000101",
			224 => "0000010000001110000101",
			225 => "0000111111100000010100",
			226 => "0010110011001000001100",
			227 => "0010111010000100000100",
			228 => "1111111000001110111001",
			229 => "0010011000111000000100",
			230 => "0000001000001110111001",
			231 => "1111111000001110111001",
			232 => "0000110011000100000100",
			233 => "1111111000001110111001",
			234 => "0000001000001110111001",
			235 => "0000110000100000000100",
			236 => "0000000000001110111001",
			237 => "0000001000001110111001",
			238 => "0000111111100000010100",
			239 => "0010110011001000001100",
			240 => "0010111010000100000100",
			241 => "1111111000001111110101",
			242 => "0010110011000000000100",
			243 => "1111111000001111110101",
			244 => "1111111000001111110101",
			245 => "0010101001000000000100",
			246 => "1111111000001111110101",
			247 => "0000001000001111110101",
			248 => "0000001011110100000100",
			249 => "0000011000001111110101",
			250 => "0001000000100000000100",
			251 => "0000000000001111110101",
			252 => "0000010000001111110101",
			253 => "0011001101101000000100",
			254 => "1111111000010000100001",
			255 => "0000110000100000010000",
			256 => "0000000101000100001000",
			257 => "0001001101101000000100",
			258 => "0000000000010000100001",
			259 => "0000001000010000100001",
			260 => "0010111000111000000100",
			261 => "1111111000010000100001",
			262 => "0000000000010000100001",
			263 => "0000001000010000100001",
			264 => "0001010011101100010100",
			265 => "0010111010000100000100",
			266 => "1111111000010001001101",
			267 => "0000000100110100001000",
			268 => "0000111011000000000100",
			269 => "0000000000010001001101",
			270 => "0000000000010001001101",
			271 => "0011001100110000000100",
			272 => "0000000000010001001101",
			273 => "0000000000010001001101",
			274 => "0000001000010001001101",
			275 => "0000111011000000000100",
			276 => "0000000000010001111001",
			277 => "0011001101101000000100",
			278 => "0000000000010001111001",
			279 => "0011111100011000001000",
			280 => "0000100111111100000100",
			281 => "0000000000010001111001",
			282 => "0000000000010001111001",
			283 => "0000110000100000000100",
			284 => "0000000000010001111001",
			285 => "0000000000010001111001",
			286 => "0010101010011000011000",
			287 => "0010111010000100001000",
			288 => "0001001111100000000100",
			289 => "1111111000010010101101",
			290 => "0000000000010010101101",
			291 => "0000000100110100001000",
			292 => "0001000110000000000100",
			293 => "1111111000010010101101",
			294 => "0000001000010010101101",
			295 => "0010001000111000000100",
			296 => "0000000000010010101101",
			297 => "1111111000010010101101",
			298 => "0000001000010010101101",
			299 => "0010111101101000001000",
			300 => "0001001111100000000100",
			301 => "1111111000010011100001",
			302 => "0000000000010011100001",
			303 => "0000111011000000000100",
			304 => "0000000000010011100001",
			305 => "0011110011101000001100",
			306 => "0000010110110100000100",
			307 => "0000001000010011100001",
			308 => "0000001110011100000100",
			309 => "0000000000010011100001",
			310 => "0000000000010011100001",
			311 => "0000000000010011100001",
			312 => "0000111011000000000100",
			313 => "0000000000010100010101",
			314 => "0010111101101000001100",
			315 => "0001101110000000001000",
			316 => "0000111100110100000100",
			317 => "0000000000010100010101",
			318 => "0000000000010100010101",
			319 => "0000000000010100010101",
			320 => "0000101011001000000100",
			321 => "0000000000010100010101",
			322 => "0000010011010000000100",
			323 => "0000000000010100010101",
			324 => "0000000000010100010101",
			325 => "0010101001111100010100",
			326 => "0000111111100000010000",
			327 => "0010111000111000001100",
			328 => "0010101110010100000100",
			329 => "1101011000010101000001",
			330 => "0000000000100100000100",
			331 => "1101100000010101000001",
			332 => "1101011000010101000001",
			333 => "1101100000010101000001",
			334 => "1101101000010101000001",
			335 => "1110110000010101000001",
			336 => "0000111111100000011000",
			337 => "0010111000111000010100",
			338 => "0010101110010100001100",
			339 => "0010111010000100000100",
			340 => "1111111000010101111101",
			341 => "0001111001010100000100",
			342 => "0000000000010101111101",
			343 => "1111111000010101111101",
			344 => "0000000010101000000100",
			345 => "0000000000010101111101",
			346 => "1111111000010101111101",
			347 => "0000000000010101111101",
			348 => "0010101010011000000100",
			349 => "0000001000010101111101",
			350 => "0000010000010101111101",
			351 => "0010111101101000001000",
			352 => "0001010000010100000100",
			353 => "1111111000010110111001",
			354 => "0000000000010110111001",
			355 => "0000111011000000000100",
			356 => "1111111000010110111001",
			357 => "0000101011001000001100",
			358 => "0000001011110100000100",
			359 => "0000001000010110111001",
			360 => "0001100101001000000100",
			361 => "0000000000010110111001",
			362 => "0000001000010110111001",
			363 => "0000110011010100000100",
			364 => "1111111000010110111001",
			365 => "0000001000010110111001",
			366 => "0010100001101000010100",
			367 => "0000110011110100001100",
			368 => "0000111011000000000100",
			369 => "1111111000011000001101",
			370 => "0001111100000000000100",
			371 => "0000001000011000001101",
			372 => "1111111000011000001101",
			373 => "0011101010110100000100",
			374 => "0000001000011000001101",
			375 => "1111111000011000001101",
			376 => "0010111101101000001000",
			377 => "0011111110111100000100",
			378 => "0000000000011000001101",
			379 => "1111111000011000001101",
			380 => "0000100111111100001000",
			381 => "0010100110100000000100",
			382 => "0000001000011000001101",
			383 => "0000001000011000001101",
			384 => "0000110001001100000100",
			385 => "0000000000011000001101",
			386 => "0000001000011000001101",
			387 => "0000110000100000011100",
			388 => "0010111010000100001000",
			389 => "0011000101111000000100",
			390 => "1111111000011001001001",
			391 => "0000000000011001001001",
			392 => "0000010110110100001000",
			393 => "0001001100101000000100",
			394 => "0000000000011001001001",
			395 => "0000001000011001001001",
			396 => "0011001100110000000100",
			397 => "1111111000011001001001",
			398 => "0010101000100000000100",
			399 => "0000000000011001001001",
			400 => "0000000000011001001001",
			401 => "0000001000011001001001",
			402 => "0000111011000000000100",
			403 => "0000000000011001111101",
			404 => "0011001101101000000100",
			405 => "0000000000011001111101",
			406 => "0000100011111100000100",
			407 => "0000000000011001111101",
			408 => "0001100100001100001000",
			409 => "0010000000110000000100",
			410 => "0000000000011001111101",
			411 => "0000000000011001111101",
			412 => "0011110011101000000100",
			413 => "0000000000011001111101",
			414 => "0000000000011001111101",
			415 => "0010110110000000001100",
			416 => "0010111001000100000100",
			417 => "1111111000011011001001",
			418 => "0001010001001000000100",
			419 => "0000000000011011001001",
			420 => "0000000000011011001001",
			421 => "0000111011000000000100",
			422 => "1111111000011011001001",
			423 => "0000101011001000010000",
			424 => "0000010110110100001000",
			425 => "0001100010000000000100",
			426 => "0000001000011011001001",
			427 => "0000000000011011001001",
			428 => "0011001100110000000100",
			429 => "0000000000011011001001",
			430 => "0000001000011011001001",
			431 => "0000110110100000000100",
			432 => "1111111000011011001001",
			433 => "0000001000011011001001",
			434 => "0011001101101000000100",
			435 => "1111111000011100011111",
			436 => "0000010110110100001100",
			437 => "0000111011000000000100",
			438 => "0000000000011100011111",
			439 => "0011110110110000000100",
			440 => "0000001000011100011111",
			441 => "0000000000011100011111",
			442 => "0011001100110000010100",
			443 => "0010001000000000001100",
			444 => "0010011100010000000100",
			445 => "0000000000011100011111",
			446 => "0000001001111100000100",
			447 => "0000000000011100011111",
			448 => "0000000000011100011111",
			449 => "0010011111101000000100",
			450 => "1111111000011100011111",
			451 => "0000000000011100011111",
			452 => "0000111100110100000100",
			453 => "0000000000011100011111",
			454 => "0000000000011100011111",
			455 => "0010111101101000000100",
			456 => "0000000000011100111001",
			457 => "0001001010000100000100",
			458 => "0000000000011100111001",
			459 => "0011110011101000000100",
			460 => "0000000000011100111001",
			461 => "0000000000011100111001",
			462 => "0010101001111100001100",
			463 => "0011001000000100000100",
			464 => "0000000000011101011101",
			465 => "0010101100001100000100",
			466 => "0000000000011101011101",
			467 => "0000000000011101011101",
			468 => "0001000000100000000100",
			469 => "0000000000011101011101",
			470 => "0000000000011101011101",
			471 => "0000110000100000010000",
			472 => "0000100000010100001000",
			473 => "0010101101001000000100",
			474 => "0000000000011110000001",
			475 => "0000000000011110000001",
			476 => "0011001100110000000100",
			477 => "0000000000011110000001",
			478 => "0000000000011110000001",
			479 => "0000000000011110000001",
			480 => "0011001101101000000100",
			481 => "0000000000011110100101",
			482 => "0000100011111100001000",
			483 => "0001001010000100000100",
			484 => "0000000000011110100101",
			485 => "0000000000011110100101",
			486 => "0000110000100000000100",
			487 => "0000000000011110100101",
			488 => "0000000000011110100101",
			489 => "0010101001111100010000",
			490 => "0011110001101000001000",
			491 => "0000111101001000000100",
			492 => "0000000000011111001001",
			493 => "0000000000011111001001",
			494 => "0011001100110000000100",
			495 => "0000000000011111001001",
			496 => "0000000000011111001001",
			497 => "0000000000011111001001",
			498 => "0001010011101100010000",
			499 => "0011110001101000001000",
			500 => "0010101001010100000100",
			501 => "0000000000011111101101",
			502 => "0000000000011111101101",
			503 => "0011001100110000000100",
			504 => "0000000000011111101101",
			505 => "0000000000011111101101",
			506 => "0000000000011111101101",
			507 => "0001010011101100010000",
			508 => "0011111010011100001000",
			509 => "0000111101001000000100",
			510 => "0000000000100000010001",
			511 => "0000000000100000010001",
			512 => "0011001100110000000100",
			513 => "0000000000100000010001",
			514 => "0000000000100000010001",
			515 => "0000000000100000010001",
			516 => "0000110000100000010000",
			517 => "0011110001101000001000",
			518 => "0001011001010000000100",
			519 => "0000000000100000110101",
			520 => "0000000000100000110101",
			521 => "0011001100110000000100",
			522 => "0000000000100000110101",
			523 => "0000000000100000110101",
			524 => "0000000000100000110101",
			525 => "0000111011000000000100",
			526 => "0000000000100001011001",
			527 => "0000100011111100001000",
			528 => "0010111001000100000100",
			529 => "0000000000100001011001",
			530 => "0000000000100001011001",
			531 => "0000110000100000000100",
			532 => "0000000000100001011001",
			533 => "0000000000100001011001",
			534 => "0001010011101100010000",
			535 => "0011110001101000001000",
			536 => "0001011001010000000100",
			537 => "0000000000100001111101",
			538 => "0000000000100001111101",
			539 => "0011001100110000000100",
			540 => "0000000000100001111101",
			541 => "0000000000100001111101",
			542 => "0000000000100001111101",
			543 => "0010101001111100010000",
			544 => "0000101101101100001000",
			545 => "0010101101001000000100",
			546 => "0000000000100010101001",
			547 => "0000000000100010101001",
			548 => "0011001100110000000100",
			549 => "1111111000100010101001",
			550 => "0000000000100010101001",
			551 => "0000011110011000000100",
			552 => "0000000000100010101001",
			553 => "0000000000100010101001",
			554 => "0010101001111100010000",
			555 => "0000101100100000001000",
			556 => "0000111101001000000100",
			557 => "0000000000100011010101",
			558 => "0000000000100011010101",
			559 => "0011001100110000000100",
			560 => "0000000000100011010101",
			561 => "0000000000100011010101",
			562 => "0000010011010000000100",
			563 => "0000000000100011010101",
			564 => "0000000000100011010101",
			565 => "0011001101101000000100",
			566 => "1111111000100011111001",
			567 => "0000111011000000000100",
			568 => "1111111000100011111001",
			569 => "0000100011111100000100",
			570 => "0000001000100011111001",
			571 => "0000110000100000000100",
			572 => "1111111000100011111001",
			573 => "0000001000100011111001",
			574 => "0011001101101000000100",
			575 => "0000000000100100011101",
			576 => "0000111011000000000100",
			577 => "0000000000100100011101",
			578 => "0000101011001000000100",
			579 => "0000000000100100011101",
			580 => "0000110110100000000100",
			581 => "0000000000100100011101",
			582 => "0000000000100100011101",
			583 => "0001010011101100010000",
			584 => "0010111010000100000100",
			585 => "0000000000100101000001",
			586 => "0000000111001100001000",
			587 => "0000111011000000000100",
			588 => "0000000000100101000001",
			589 => "0000000000100101000001",
			590 => "0000000000100101000001",
			591 => "0000000000100101000001",
			592 => "0000111011000000000100",
			593 => "0000000000100101100101",
			594 => "0011001101101000000100",
			595 => "0000000000100101100101",
			596 => "0000101011001000000100",
			597 => "0000000000100101100101",
			598 => "0000011110011000000100",
			599 => "0000000000100101100101",
			600 => "0000000000100101100101",
			601 => "0010101010011000010000",
			602 => "0000100111000000001100",
			603 => "0000111011000000000100",
			604 => "0000000000100110001001",
			605 => "0011001001000100000100",
			606 => "0000000000100110001001",
			607 => "0000000000100110001001",
			608 => "0000000000100110001001",
			609 => "0000000000100110001001",
			610 => "0010101001111100010000",
			611 => "0010111010000100000100",
			612 => "1111111000100110110101",
			613 => "0000111011000000000100",
			614 => "1111111000100110110101",
			615 => "0000101110011100000100",
			616 => "0000001000100110110101",
			617 => "1111111000100110110101",
			618 => "0001010011101100000100",
			619 => "0000000000100110110101",
			620 => "0000001000100110110101",
			621 => "0010111101101000001000",
			622 => "0001001111100000000100",
			623 => "0000000000100111100001",
			624 => "0000000000100111100001",
			625 => "0001001010000100000100",
			626 => "0000000000100111100001",
			627 => "0000101011001000000100",
			628 => "0000000000100111100001",
			629 => "0000110110100000000100",
			630 => "0000000000100111100001",
			631 => "0000000000100111100001",
			632 => "0010111101101000001000",
			633 => "0011000101111000000100",
			634 => "0000000000101000001101",
			635 => "0000000000101000001101",
			636 => "0001001010000100000100",
			637 => "0000000000101000001101",
			638 => "0000101011001000000100",
			639 => "0000000000101000001101",
			640 => "0000110110100000000100",
			641 => "0000000000101000001101",
			642 => "0000000000101000001101",
			643 => "0010100001101000001100",
			644 => "0001110011001000001000",
			645 => "0000111011111000000100",
			646 => "0000000000101001000001",
			647 => "0000000000101001000001",
			648 => "0000000000101001000001",
			649 => "0000100011111100001000",
			650 => "0010111001000100000100",
			651 => "0000000000101001000001",
			652 => "0000000000101001000001",
			653 => "0000110000100000000100",
			654 => "0000000000101001000001",
			655 => "0000000000101001000001",
			656 => "0001010011101100010100",
			657 => "0011110001101000001000",
			658 => "0001011001010000000100",
			659 => "0000000000101001101101",
			660 => "0000000000101001101101",
			661 => "0011001100110000000100",
			662 => "0000000000101001101101",
			663 => "0011001000101000000100",
			664 => "0000000000101001101101",
			665 => "0000000000101001101101",
			666 => "0000000000101001101101",
			667 => "0000111111100000010100",
			668 => "0010110011001000001100",
			669 => "0010111010000100000100",
			670 => "1111111000101010100001",
			671 => "0001111001010100000100",
			672 => "0000000000101010100001",
			673 => "1111111000101010100001",
			674 => "0010101110111000000100",
			675 => "1111111000101010100001",
			676 => "0000010000101010100001",
			677 => "0010101010011000000100",
			678 => "0000001000101010100001",
			679 => "0000001000101010100001",
			680 => "0000111111100000010100",
			681 => "0000110011110100001100",
			682 => "0000111011000000000100",
			683 => "1111111000101011010101",
			684 => "0000000101000000000100",
			685 => "0000001000101011010101",
			686 => "1111111000101011010101",
			687 => "0000000100011000000100",
			688 => "0000010000101011010101",
			689 => "1111111000101011010101",
			690 => "0000110000100000000100",
			691 => "0000000000101011010101",
			692 => "0000001000101011010101",
			693 => "0000111111100000010100",
			694 => "0010100001101000001100",
			695 => "0000111011000000000100",
			696 => "1111111000101100010001",
			697 => "0001111100000000000100",
			698 => "0000000000101100010001",
			699 => "1111111000101100010001",
			700 => "0011111111000100000100",
			701 => "0000010000101100010001",
			702 => "1111111000101100010001",
			703 => "0010101001111100000100",
			704 => "0000001000101100010001",
			705 => "0000010011010000000100",
			706 => "0000001000101100010001",
			707 => "0000001000101100010001",
			708 => "0011001101101000000100",
			709 => "1111111000101100111101",
			710 => "0000110000100000010000",
			711 => "0000000101000100001000",
			712 => "0001001101101000000100",
			713 => "0000000000101100111101",
			714 => "0000001000101100111101",
			715 => "0010111000111000000100",
			716 => "1111111000101100111101",
			717 => "0000000000101100111101",
			718 => "0000001000101100111101",
			719 => "0001010011101100010100",
			720 => "0010111010000100000100",
			721 => "1111111000101101101001",
			722 => "0000000100110100001000",
			723 => "0000111011000000000100",
			724 => "0000000000101101101001",
			725 => "0000000000101101101001",
			726 => "0011001100110000000100",
			727 => "0000000000101101101001",
			728 => "0000000000101101101001",
			729 => "0000001000101101101001",
			730 => "0010101001111100011000",
			731 => "0011001000000100001100",
			732 => "0010111010000100000100",
			733 => "1111111000101110100101",
			734 => "0011000011000000000100",
			735 => "0000001000101110100101",
			736 => "1111111000101110100101",
			737 => "0000000110001000001000",
			738 => "0000111001000100000100",
			739 => "1111111000101110100101",
			740 => "0000001000101110100101",
			741 => "1111111000101110100101",
			742 => "0000010011010000000100",
			743 => "0000001000101110100101",
			744 => "0000001000101110100101",
			745 => "0010101010011000011000",
			746 => "0010111010000100001000",
			747 => "0011000101111000000100",
			748 => "1111111000101111011001",
			749 => "0000000000101111011001",
			750 => "0000000100110100001000",
			751 => "0001001001000100000100",
			752 => "1111111000101111011001",
			753 => "0000001000101111011001",
			754 => "0011011010000100000100",
			755 => "0000000000101111011001",
			756 => "1111111000101111011001",
			757 => "0000001000101111011001",
			758 => "0010101001111100010100",
			759 => "0010111010000100000100",
			760 => "1111111000110000001101",
			761 => "0001111001010100000100",
			762 => "0000000000110000001101",
			763 => "0011001100110000001000",
			764 => "0011010101101100000100",
			765 => "0000000000110000001101",
			766 => "0000000000110000001101",
			767 => "0000000000110000001101",
			768 => "0000011110011000000100",
			769 => "0000000000110000001101",
			770 => "0000000000110000001101",
			771 => "0000111011000000000100",
			772 => "0000000000110001000001",
			773 => "0010111101101000001100",
			774 => "0001101110000000001000",
			775 => "0000100000000100000100",
			776 => "0000000000110001000001",
			777 => "0000000000110001000001",
			778 => "0000000000110001000001",
			779 => "0000101011001000000100",
			780 => "0000000000110001000001",
			781 => "0000010111011100000100",
			782 => "0000000000110001000001",
			783 => "0000000000110001000001",
			784 => "0010100001101000001100",
			785 => "0010111010000100000100",
			786 => "1111111000110010000101",
			787 => "0001111001010100000100",
			788 => "0000001000110010000101",
			789 => "1111111000110010000101",
			790 => "0010111101101000001000",
			791 => "0001101110000000000100",
			792 => "0000000000110010000101",
			793 => "1111111000110010000101",
			794 => "0000100111111100001000",
			795 => "0010100110100000000100",
			796 => "0000001000110010000101",
			797 => "0000001000110010000101",
			798 => "0001000010001000000100",
			799 => "0000000000110010000101",
			800 => "0000001000110010000101",
			801 => "0010111101101000001000",
			802 => "0001001111100000000100",
			803 => "1111111000110011000001",
			804 => "0000000000110011000001",
			805 => "0000111011000000000100",
			806 => "1111111000110011000001",
			807 => "0000101011001000001100",
			808 => "0011001111011000000100",
			809 => "0000001000110011000001",
			810 => "0000100111111100000100",
			811 => "0000001000110011000001",
			812 => "0000000000110011000001",
			813 => "0000110110100000000100",
			814 => "1111111000110011000001",
			815 => "0000001000110011000001",
			816 => "0010111101101000001000",
			817 => "0001010000010100000100",
			818 => "1111111000110011111101",
			819 => "0000000000110011111101",
			820 => "0000111011000000000100",
			821 => "1111111000110011111101",
			822 => "0000011011101100001000",
			823 => "0000101011100000000100",
			824 => "0000001000110011111101",
			825 => "0000000000110011111101",
			826 => "0011001100110000001000",
			827 => "0010001000111000000100",
			828 => "0000000000110011111101",
			829 => "1111111000110011111101",
			830 => "0000001000110011111101",
			831 => "0010100001101000010100",
			832 => "0010101100110100001100",
			833 => "0000111011000000000100",
			834 => "1111111000110101010001",
			835 => "0000000101000000000100",
			836 => "0000001000110101010001",
			837 => "1111111000110101010001",
			838 => "0001000000111100000100",
			839 => "0000001000110101010001",
			840 => "1111111000110101010001",
			841 => "0010111101101000001000",
			842 => "0001101110000000000100",
			843 => "0000000000110101010001",
			844 => "1111111000110101010001",
			845 => "0000100111111100001000",
			846 => "0010100110100000000100",
			847 => "0000001000110101010001",
			848 => "0000001000110101010001",
			849 => "0000110001001100000100",
			850 => "0000000000110101010001",
			851 => "0000001000110101010001",
			852 => "0000110000100000011100",
			853 => "0010111010000100001000",
			854 => "0011000101111000000100",
			855 => "1111111000110110001101",
			856 => "0000000000110110001101",
			857 => "0000010110110100001000",
			858 => "0001001100101000000100",
			859 => "0000000000110110001101",
			860 => "0000001000110110001101",
			861 => "0011001100110000000100",
			862 => "1111111000110110001101",
			863 => "0010101000100000000100",
			864 => "0000000000110110001101",
			865 => "0000000000110110001101",
			866 => "0000001000110110001101",
			867 => "0000111011000000000100",
			868 => "0000000000110111000001",
			869 => "0011001101101000000100",
			870 => "0000000000110111000001",
			871 => "0000100011111100000100",
			872 => "0000000000110111000001",
			873 => "0001100100001100001000",
			874 => "0010000000110000000100",
			875 => "0000000000110111000001",
			876 => "0000000000110111000001",
			877 => "0011110011101000000100",
			878 => "0000000000110111000001",
			879 => "0000000000110111000001",
			880 => "0010111101101000001000",
			881 => "0001010000010100000100",
			882 => "1111111000111000001111",
			883 => "0000000000111000001111",
			884 => "0000010110110100001000",
			885 => "0000111011000000000100",
			886 => "0000000000111000001111",
			887 => "0000001000111000001111",
			888 => "0011001100110000010000",
			889 => "0010001000000000001000",
			890 => "0000111110001100000100",
			891 => "0000000000111000001111",
			892 => "0000000000111000001111",
			893 => "0010011111101000000100",
			894 => "1111111000111000001111",
			895 => "0000000000111000001111",
			896 => "0000111100110100000100",
			897 => "0000000000111000001111",
			898 => "0000001000111000001111",
			899 => "0000111011000000000100",
			900 => "0000000000111000101001",
			901 => "0011001101101000000100",
			902 => "0000000000111000101001",
			903 => "0011110011101000000100",
			904 => "0000000000111000101001",
			905 => "0000000000111000101001",
			906 => "0000110000100000010000",
			907 => "0011110001101000001000",
			908 => "0010101000101000000100",
			909 => "0000000000111001001101",
			910 => "0000000000111001001101",
			911 => "0011001100110000000100",
			912 => "1111111000111001001101",
			913 => "0000000000111001001101",
			914 => "0000001000111001001101",
			915 => "0010101001111100010000",
			916 => "0011110001101000001000",
			917 => "0010101000101000000100",
			918 => "0000000000111001110001",
			919 => "0000000000111001110001",
			920 => "0011001100110000000100",
			921 => "0000000000111001110001",
			922 => "0000000000111001110001",
			923 => "0000000000111001110001",
			924 => "0011001101101000000100",
			925 => "0000000000111010010101",
			926 => "0000100011111100001000",
			927 => "0000111011000000000100",
			928 => "0000000000111010010101",
			929 => "0000000000111010010101",
			930 => "0000110000100000000100",
			931 => "0000000000111010010101",
			932 => "0000000000111010010101",
			933 => "0010101001111100010000",
			934 => "0011110001101000001000",
			935 => "0000111101001000000100",
			936 => "0000000000111010111001",
			937 => "0000000000111010111001",
			938 => "0011001100110000000100",
			939 => "0000000000111010111001",
			940 => "0000000000111010111001",
			941 => "0000000000111010111001",
			942 => "0001010011101100010000",
			943 => "0011110001101000001000",
			944 => "0010101001010100000100",
			945 => "0000000000111011011101",
			946 => "0000000000111011011101",
			947 => "0011001100110000000100",
			948 => "0000000000111011011101",
			949 => "0000000000111011011101",
			950 => "0000000000111011011101",
			951 => "0010101100110100000100",
			952 => "0000000000111100000001",
			953 => "0000100011111100001000",
			954 => "0010111001000100000100",
			955 => "0000000000111100000001",
			956 => "0000000000111100000001",
			957 => "0000110000100000000100",
			958 => "0000000000111100000001",
			959 => "0000000000111100000001",
			960 => "0010101010011000010000",
			961 => "0011110001101000001000",
			962 => "0001011001010000000100",
			963 => "0000000000111100100101",
			964 => "0000000000111100100101",
			965 => "0011001100110000000100",
			966 => "0000000000111100100101",
			967 => "0000000000111100100101",
			968 => "0000000000111100100101",
			969 => "0001010011101100010000",
			970 => "0011111010011100001000",
			971 => "0000111101001000000100",
			972 => "0000000000111101001001",
			973 => "0000000000111101001001",
			974 => "0011001100110000000100",
			975 => "0000000000111101001001",
			976 => "0000000000111101001001",
			977 => "0000000000111101001001",
			978 => "0001010011101100010000",
			979 => "0011110001101000001000",
			980 => "0001011001010000000100",
			981 => "0000000000111101101101",
			982 => "0000000000111101101101",
			983 => "0011001100110000000100",
			984 => "0000000000111101101101",
			985 => "0000000000111101101101",
			986 => "0000000000111101101101",
			987 => "0010101001111100010000",
			988 => "0011110001101000001000",
			989 => "0000111101001000000100",
			990 => "0000000000111110011001",
			991 => "0000000000111110011001",
			992 => "0011001100110000000100",
			993 => "1111111000111110011001",
			994 => "0000000000111110011001",
			995 => "0000101011001000000100",
			996 => "0000000000111110011001",
			997 => "0000000000111110011001",
			998 => "0010101001111100010000",
			999 => "0011001000000100000100",
			1000 => "1111111000111110111101",
			1001 => "0000000110001000001000",
			1002 => "0001001100101000000100",
			1003 => "0000000000111110111101",
			1004 => "0000001000111110111101",
			1005 => "1111111000111110111101",
			1006 => "0000001000111110111101",
			1007 => "0011001101101000000100",
			1008 => "1111111000111111100001",
			1009 => "0000111011000000000100",
			1010 => "1111111000111111100001",
			1011 => "0000100011111100000100",
			1012 => "0000001000111111100001",
			1013 => "0000110000100000000100",
			1014 => "1111111000111111100001",
			1015 => "0000001000111111100001",
			1016 => "0011001101101000000100",
			1017 => "0000000001000000000101",
			1018 => "0000111011000000000100",
			1019 => "0000000001000000000101",
			1020 => "0000101011100000000100",
			1021 => "0000000001000000000101",
			1022 => "0000110010010100000100",
			1023 => "0000000001000000000101",
			1024 => "0000000001000000000101",
			1025 => "0000110000100000010000",
			1026 => "0000100111000000001100",
			1027 => "0000111011000000000100",
			1028 => "0000000001000000101001",
			1029 => "0011010101011100000100",
			1030 => "0000000001000000101001",
			1031 => "0000000001000000101001",
			1032 => "0000000001000000101001",
			1033 => "0000000001000000101001",
			1034 => "0000111011000000000100",
			1035 => "0000000001000001001101",
			1036 => "0011001101101000000100",
			1037 => "0000000001000001001101",
			1038 => "0000101011001000000100",
			1039 => "0000000001000001001101",
			1040 => "0000011110011000000100",
			1041 => "0000000001000001001101",
			1042 => "0000000001000001001101",
			1043 => "0010101001111100010000",
			1044 => "0010111010000100000100",
			1045 => "1111111001000001111001",
			1046 => "0000111011000000000100",
			1047 => "1111111001000001111001",
			1048 => "0000001000011100000100",
			1049 => "0000001001000001111001",
			1050 => "1111111001000001111001",
			1051 => "0000010011010000000100",
			1052 => "0000001001000001111001",
			1053 => "0000001001000001111001",
			1054 => "0010111101101000001000",
			1055 => "0001001111100000000100",
			1056 => "1111111001000010100101",
			1057 => "0000000001000010100101",
			1058 => "0000111011000000000100",
			1059 => "0000000001000010100101",
			1060 => "0000100111111100000100",
			1061 => "0000001001000010100101",
			1062 => "0000110000100000000100",
			1063 => "0000000001000010100101",
			1064 => "0000000001000010100101",
			1065 => "0010111101101000001000",
			1066 => "0001001111100000000100",
			1067 => "0000000001000011010001",
			1068 => "0000000001000011010001",
			1069 => "0001001010000100000100",
			1070 => "0000000001000011010001",
			1071 => "0000101011001000000100",
			1072 => "0000000001000011010001",
			1073 => "0000110110100000000100",
			1074 => "0000000001000011010001",
			1075 => "0000000001000011010001",
			1076 => "0010100001101000001100",
			1077 => "0010101100110100000100",
			1078 => "0000000001000100000101",
			1079 => "0010100000111000000100",
			1080 => "0000000001000100000101",
			1081 => "0000000001000100000101",
			1082 => "0000100011111100001000",
			1083 => "0010111001000100000100",
			1084 => "0000000001000100000101",
			1085 => "0000000001000100000101",
			1086 => "0000110000100000000100",
			1087 => "0000000001000100000101",
			1088 => "0000000001000100000101",
			1089 => "0000110000100000010100",
			1090 => "0011001000000100001000",
			1091 => "0001000010001100000100",
			1092 => "1111111001000100110001",
			1093 => "0000000001000100110001",
			1094 => "0000000110001000001000",
			1095 => "0001000110000000000100",
			1096 => "1111111001000100110001",
			1097 => "0000001001000100110001",
			1098 => "1111111001000100110001",
			1099 => "0000001001000100110001",
			1100 => "0001010011101100010100",
			1101 => "0011110001101000001000",
			1102 => "0010101001010100000100",
			1103 => "0000000001000101011101",
			1104 => "0000000001000101011101",
			1105 => "0011001100110000000100",
			1106 => "0000000001000101011101",
			1107 => "0011001000101000000100",
			1108 => "0000000001000101011101",
			1109 => "0000000001000101011101",
			1110 => "0000000001000101011101",
			1111 => "0000111111100000010100",
			1112 => "0010110011001000001100",
			1113 => "0010111010000100000100",
			1114 => "1111111001000110010001",
			1115 => "0001111001010100000100",
			1116 => "0000000001000110010001",
			1117 => "1111111001000110010001",
			1118 => "0010101110111000000100",
			1119 => "1111111001000110010001",
			1120 => "0000001001000110010001",
			1121 => "0010101010011000000100",
			1122 => "0000001001000110010001",
			1123 => "0000001001000110010001",
			1124 => "0010101001111100010100",
			1125 => "0011001000000100001100",
			1126 => "0010111010000100000100",
			1127 => "1111111001000111000101",
			1128 => "0011000011000000000100",
			1129 => "0000001001000111000101",
			1130 => "1111111001000111000101",
			1131 => "0010101010011100000100",
			1132 => "1111111001000111000101",
			1133 => "0000001001000111000101",
			1134 => "0000010011010000000100",
			1135 => "0000001001000111000101",
			1136 => "0000001001000111000101",
			1137 => "0010111101101000001000",
			1138 => "0001001111100000000100",
			1139 => "1111111001000111111001",
			1140 => "0000000001000111111001",
			1141 => "0000111011000000000100",
			1142 => "1111111001000111111001",
			1143 => "0000101011001000001000",
			1144 => "0011011111011000000100",
			1145 => "0000001001000111111001",
			1146 => "0000000001000111111001",
			1147 => "0000110110100000000100",
			1148 => "1111111001000111111001",
			1149 => "0000001001000111111001",
			1150 => "0011001101101000000100",
			1151 => "1111111001001000100101",
			1152 => "0000111011000000000100",
			1153 => "0000000001001000100101",
			1154 => "0000011011101100001000",
			1155 => "0011110110110000000100",
			1156 => "0000001001001000100101",
			1157 => "0000000001001000100101",
			1158 => "0000001000100100000100",
			1159 => "0000000001001000100101",
			1160 => "0000000001001000100101",
			1161 => "0010101001111100010100",
			1162 => "0010111010000100000100",
			1163 => "1111111001001001010001",
			1164 => "0001101110010100001000",
			1165 => "0000101000000100000100",
			1166 => "0000000001001001010001",
			1167 => "0000000001001001010001",
			1168 => "0011001100110000000100",
			1169 => "0000000001001001010001",
			1170 => "0000000001001001010001",
			1171 => "0000000001001001010001",
			1172 => "0010101010011000011000",
			1173 => "0010111010000100001000",
			1174 => "0001001111100000000100",
			1175 => "1111111001001010000101",
			1176 => "0000000001001010000101",
			1177 => "0000000100110100001000",
			1178 => "0001000110000000000100",
			1179 => "1111111001001010000101",
			1180 => "0000001001001010000101",
			1181 => "0011011010000100000100",
			1182 => "0000000001001010000101",
			1183 => "1111111001001010000101",
			1184 => "0000001001001010000101",
			1185 => "0010111101101000001000",
			1186 => "0001001111100000000100",
			1187 => "1111111001001010111001",
			1188 => "0000000001001010111001",
			1189 => "0000111011000000000100",
			1190 => "0000000001001010111001",
			1191 => "0011110011101000001100",
			1192 => "0000010110110100000100",
			1193 => "0000001001001010111001",
			1194 => "0000001110011100000100",
			1195 => "0000000001001010111001",
			1196 => "0000000001001010111001",
			1197 => "0000000001001010111001",
			1198 => "0000111011000000000100",
			1199 => "0000000001001011101101",
			1200 => "0010111101101000001100",
			1201 => "0011111001110000001000",
			1202 => "0000100000000100000100",
			1203 => "0000000001001011101101",
			1204 => "0000000001001011101101",
			1205 => "0000000001001011101101",
			1206 => "0000101011001000000100",
			1207 => "0000000001001011101101",
			1208 => "0000010111011100000100",
			1209 => "0000000001001011101101",
			1210 => "0000000001001011101101",
			1211 => "0000111011000000000100",
			1212 => "0000000001001100100001",
			1213 => "0010111101101000001100",
			1214 => "0001101110000000001000",
			1215 => "0000100000000100000100",
			1216 => "0000000001001100100001",
			1217 => "0000000001001100100001",
			1218 => "0000000001001100100001",
			1219 => "0000101011001000000100",
			1220 => "0000000001001100100001",
			1221 => "0000010111011100000100",
			1222 => "0000000001001100100001",
			1223 => "0000000001001100100001",
			1224 => "0000110100000000010100",
			1225 => "0010111000111000010000",
			1226 => "0010101101111100001100",
			1227 => "0010101110010100000100",
			1228 => "1111111001001101011101",
			1229 => "0010001111001000000100",
			1230 => "1111111001001101011101",
			1231 => "0000000001001101011101",
			1232 => "0000000001001101011101",
			1233 => "0000000001001101011101",
			1234 => "0000000010101000000100",
			1235 => "0000100001001101011101",
			1236 => "0010111010000100000100",
			1237 => "0000011001001101011101",
			1238 => "0000011001001101011101",
			1239 => "0010111101101000001000",
			1240 => "0001001111100000000100",
			1241 => "1111111001001110011001",
			1242 => "0000000001001110011001",
			1243 => "0000111011000000000100",
			1244 => "1111111001001110011001",
			1245 => "0000101011001000001100",
			1246 => "0011001111011000000100",
			1247 => "0000001001001110011001",
			1248 => "0000100111111100000100",
			1249 => "0000001001001110011001",
			1250 => "0000000001001110011001",
			1251 => "0000110110100000000100",
			1252 => "1111111001001110011001",
			1253 => "0000001001001110011001",
			1254 => "0010111101101000001000",
			1255 => "0001001111100000000100",
			1256 => "1111111001001111010101",
			1257 => "0000000001001111010101",
			1258 => "0000111011000000000100",
			1259 => "1111111001001111010101",
			1260 => "0000101011001000001100",
			1261 => "0000010110110100000100",
			1262 => "0000001001001111010101",
			1263 => "0000010101010100000100",
			1264 => "0000000001001111010101",
			1265 => "0000001001001111010101",
			1266 => "0000110110100000000100",
			1267 => "1111111001001111010101",
			1268 => "0000001001001111010101",
			1269 => "0010101100110100000100",
			1270 => "1111111001010000010001",
			1271 => "0010111101101000010000",
			1272 => "0011111001110000000100",
			1273 => "0000000001010000010001",
			1274 => "0000000011011100000100",
			1275 => "1111111001010000010001",
			1276 => "0000001010000000000100",
			1277 => "0000000001010000010001",
			1278 => "1111111001010000010001",
			1279 => "0000101011001000001000",
			1280 => "0000100111111100000100",
			1281 => "0000001001010000010001",
			1282 => "0000001001010000010001",
			1283 => "0000000001010000010001",
			1284 => "0000111011000000000100",
			1285 => "0000000001010001000101",
			1286 => "0011001101101000000100",
			1287 => "0000000001010001000101",
			1288 => "0000100011111100000100",
			1289 => "0000000001010001000101",
			1290 => "0001100100001100001000",
			1291 => "0010000000110000000100",
			1292 => "0000000001010001000101",
			1293 => "0000000001010001000101",
			1294 => "0011110011101000000100",
			1295 => "0000000001010001000101",
			1296 => "0000000001010001000101",
			1297 => "0010110110000000001000",
			1298 => "0001011010011000000100",
			1299 => "1111111001010010001001",
			1300 => "0000000001010010001001",
			1301 => "0000111011000000000100",
			1302 => "1111111001010010001001",
			1303 => "0000101011001000010000",
			1304 => "0000010110110100001000",
			1305 => "0001111011000000000100",
			1306 => "0000001001010010001001",
			1307 => "0000001001010010001001",
			1308 => "0011001100110000000100",
			1309 => "0000000001010010001001",
			1310 => "0000001001010010001001",
			1311 => "0000110110100000000100",
			1312 => "1111111001010010001001",
			1313 => "0000001001010010001001",
			1314 => "0000111011000000000100",
			1315 => "0000000001010011000111",
			1316 => "0011001101101000000100",
			1317 => "0000000001010011000111",
			1318 => "0000100011111100000100",
			1319 => "0000000001010011000111",
			1320 => "0010111010000100001000",
			1321 => "0010001111011000000100",
			1322 => "0000000001010011000111",
			1323 => "0000000001010011000111",
			1324 => "0011110010001000000100",
			1325 => "0000000001010011000111",
			1326 => "0001100110110000000100",
			1327 => "0000000001010011000111",
			1328 => "0000000001010011000111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(455, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(899, initial_addr_3'length));
	end generate gen_rom_10;

	gen_rom_11: if SELECT_ROM = 11 generate
		bank <= (
			0 => "0000000001101100011000",
			1 => "0010111010100100001100",
			2 => "0000011000111100000100",
			3 => "0000000000000001110101",
			4 => "0011100011001000000100",
			5 => "0000000000000001110101",
			6 => "0000000000000001110101",
			7 => "0001101000111000001000",
			8 => "0001111111011000000100",
			9 => "0000000000000001110101",
			10 => "0000000000000001110101",
			11 => "0000000000000001110101",
			12 => "0011011011101100010100",
			13 => "0001100010001100000100",
			14 => "0000000000000001110101",
			15 => "0010010111011100000100",
			16 => "0000000000000001110101",
			17 => "0011110010000000001000",
			18 => "0001001111101000000100",
			19 => "0000000000000001110101",
			20 => "0000000000000001110101",
			21 => "0000000000000001110101",
			22 => "0011001001001000001000",
			23 => "0000011000111100000100",
			24 => "0000000000000001110101",
			25 => "0000000000000001110101",
			26 => "0000101110010000000100",
			27 => "0000000000000001110101",
			28 => "0000000000000001110101",
			29 => "0000010111100100100100",
			30 => "0000110101101100010000",
			31 => "0000100000111000001000",
			32 => "0011111001001000000100",
			33 => "0000000000000011111001",
			34 => "0000000000000011111001",
			35 => "0001011001001000000100",
			36 => "0000000000000011111001",
			37 => "0000000000000011111001",
			38 => "0001011010011100001100",
			39 => "0001101110111100001000",
			40 => "0010000101101100000100",
			41 => "0000000000000011111001",
			42 => "0000000000000011111001",
			43 => "0000000000000011111001",
			44 => "0011001001001000000100",
			45 => "0000000000000011111001",
			46 => "0000000000000011111001",
			47 => "0001000101101100011000",
			48 => "0010111001001000001100",
			49 => "0001100011001000001000",
			50 => "0001001001100000000100",
			51 => "0000000000000011111001",
			52 => "0000000000000011111001",
			53 => "0000000000000011111001",
			54 => "0011111000000000000100",
			55 => "0000000000000011111001",
			56 => "0011000110000000000100",
			57 => "0000000000000011111001",
			58 => "0000000000000011111001",
			59 => "0010000101011100000100",
			60 => "0000000000000011111001",
			61 => "0000000000000011111001",
			62 => "0000011000111100010100",
			63 => "0001011010000100001000",
			64 => "0010011100101000000100",
			65 => "0000000000000101111101",
			66 => "0000000000000101111101",
			67 => "0000111111011000000100",
			68 => "0000000000000101111101",
			69 => "0001111000111000000100",
			70 => "0000000000000101111101",
			71 => "0000000000000101111101",
			72 => "0011000101011100001100",
			73 => "0001011000011000000100",
			74 => "0000000000000101111101",
			75 => "0000111011000000000100",
			76 => "0000000000000101111101",
			77 => "0000000000000101111101",
			78 => "0000010111100100010000",
			79 => "0010101000000000001000",
			80 => "0001111010000100000100",
			81 => "0000000000000101111101",
			82 => "0000000000000101111101",
			83 => "0001001001011000000100",
			84 => "0000000000000101111101",
			85 => "0000000000000101111101",
			86 => "0001000110000000001100",
			87 => "0000000010110100001000",
			88 => "0000001011111000000100",
			89 => "0000000000000101111101",
			90 => "0000000000000101111101",
			91 => "0000000000000101111101",
			92 => "0000111000000000000100",
			93 => "0000000000000101111101",
			94 => "0000000000000101111101",
			95 => "0000000001101100100000",
			96 => "0011000111011100010000",
			97 => "0000000000111000001000",
			98 => "0010110110001100000100",
			99 => "0000000000001000001001",
			100 => "0000000000001000001001",
			101 => "0011110000111000000100",
			102 => "0000000000001000001001",
			103 => "0000000000001000001001",
			104 => "0001101000111000001000",
			105 => "0001111111011000000100",
			106 => "0000000000001000001001",
			107 => "0000000000001000001001",
			108 => "0001011110011000000100",
			109 => "0000000000001000001001",
			110 => "0000000000001000001001",
			111 => "0010001111111100100000",
			112 => "0001101001101100000100",
			113 => "0000000000001000001001",
			114 => "0001100100100100010000",
			115 => "0001011001000000001000",
			116 => "0001110101111000000100",
			117 => "0000000000001000001001",
			118 => "0000000000001000001001",
			119 => "0001111100010000000100",
			120 => "0000000000001000001001",
			121 => "0000000000001000001001",
			122 => "0011000011010000000100",
			123 => "0000000000001000001001",
			124 => "0010011001001000000100",
			125 => "0000000000001000001001",
			126 => "0000000000001000001001",
			127 => "0010111000101000000100",
			128 => "0000000000001000001001",
			129 => "0000000000001000001001",
			130 => "0001010110101100101100",
			131 => "0000000000110100010000",
			132 => "0010110110001100000100",
			133 => "0000000000001010100101",
			134 => "0000101010000100000100",
			135 => "0000000000001010100101",
			136 => "0010011100110000000100",
			137 => "0000000000001010100101",
			138 => "0000000000001010100101",
			139 => "0001101001101100000100",
			140 => "0000000000001010100101",
			141 => "0001100101001000001100",
			142 => "0010001111111100000100",
			143 => "0000000000001010100101",
			144 => "0010111100101000000100",
			145 => "0000000000001010100101",
			146 => "0000000000001010100101",
			147 => "0011000011010000000100",
			148 => "0000000000001010100101",
			149 => "0011011011101100000100",
			150 => "0000000000001010100101",
			151 => "0000000000001010100101",
			152 => "0011001001001000010100",
			153 => "0010000011010000001000",
			154 => "0000111001010100000100",
			155 => "0000000000001010100101",
			156 => "0000000000001010100101",
			157 => "0011111100001100000100",
			158 => "0000000000001010100101",
			159 => "0010110101011100000100",
			160 => "0000000000001010100101",
			161 => "0000000000001010100101",
			162 => "0010001001000100001000",
			163 => "0001001001011000000100",
			164 => "0000000000001010100101",
			165 => "0000000000001010100101",
			166 => "0001001101101000000100",
			167 => "0000000000001010100101",
			168 => "0000000000001010100101",
			169 => "0001001110011000100100",
			170 => "0000111100101000011100",
			171 => "0001001001100000001100",
			172 => "0000000011000000000100",
			173 => "0000000000001101001001",
			174 => "0001001001100100000100",
			175 => "0000000000001101001001",
			176 => "0000000000001101001001",
			177 => "0001011001001000001100",
			178 => "0011001101101000001000",
			179 => "0011101001000100000100",
			180 => "0000000000001101001001",
			181 => "0000000000001101001001",
			182 => "0000000000001101001001",
			183 => "0000000000001101001001",
			184 => "0001100101110100000100",
			185 => "0000000000001101001001",
			186 => "0000000000001101001001",
			187 => "0011001001001000011000",
			188 => "0011100001001000001000",
			189 => "0000011000011000000100",
			190 => "0000000000001101001001",
			191 => "0000000000001101001001",
			192 => "0000011000111100000100",
			193 => "0000000000001101001001",
			194 => "0010110101011100000100",
			195 => "0000000000001101001001",
			196 => "0011011010100100000100",
			197 => "0000000000001101001001",
			198 => "0000000000001101001001",
			199 => "0011010011010000001000",
			200 => "0001001001011000000100",
			201 => "0000000000001101001001",
			202 => "0000000000001101001001",
			203 => "0001000101101100001100",
			204 => "0011111000111000000100",
			205 => "0000000000001101001001",
			206 => "0011011100101000000100",
			207 => "0000000000001101001001",
			208 => "0000000000001101001001",
			209 => "0000000000001101001001",
			210 => "0011100001001000100000",
			211 => "0000011000011000010000",
			212 => "0010110110001100000100",
			213 => "0000000000001111100101",
			214 => "0000101101000100001000",
			215 => "0000000011000000000100",
			216 => "0000000000001111100101",
			217 => "0000000000001111100101",
			218 => "0000000000001111100101",
			219 => "0001001110011000001100",
			220 => "0000101100010000000100",
			221 => "0000000000001111100101",
			222 => "0000100001111100000100",
			223 => "0000000000001111100101",
			224 => "0000000000001111100101",
			225 => "0000000000001111100101",
			226 => "0011001001001000100100",
			227 => "0001001110011000001100",
			228 => "0010010111011100000100",
			229 => "0000000000001111100101",
			230 => "0001101111000100000100",
			231 => "0000000000001111100101",
			232 => "0000000000001111100101",
			233 => "0000011000111100000100",
			234 => "0000000000001111100101",
			235 => "0010110101011100001100",
			236 => "0011011111011100000100",
			237 => "0000000000001111100101",
			238 => "0010000011010000000100",
			239 => "0000000000001111100101",
			240 => "0000000000001111100101",
			241 => "0011011010100100000100",
			242 => "0000000000001111100101",
			243 => "0000000000001111100101",
			244 => "0000101110010000000100",
			245 => "0000000000001111100101",
			246 => "0000010001110000000100",
			247 => "0000000000001111100101",
			248 => "0000000000001111100101",
			249 => "0001001110011000100100",
			250 => "0011000110110100000100",
			251 => "0000000000010010001001",
			252 => "0010101010100100001100",
			253 => "0000001010100000001000",
			254 => "0000101010000100000100",
			255 => "0000000000010010001001",
			256 => "0000000000010010001001",
			257 => "0000000000010010001001",
			258 => "0001101101000100001100",
			259 => "0000001001011000000100",
			260 => "0000000000010010001001",
			261 => "0000000100110000000100",
			262 => "0000000000010010001001",
			263 => "0000000000010010001001",
			264 => "0001010110000000000100",
			265 => "0000000000010010001001",
			266 => "0000000000010010001001",
			267 => "0011001001001000011000",
			268 => "0011100001001000001000",
			269 => "0011000011010000000100",
			270 => "0000000000010010001001",
			271 => "0000000000010010001001",
			272 => "0000011000111100000100",
			273 => "0000000000010010001001",
			274 => "0010110101011100000100",
			275 => "0000000000010010001001",
			276 => "0011011010100100000100",
			277 => "0000000000010010001001",
			278 => "0000000000010010001001",
			279 => "0011010011010000001000",
			280 => "0001001001011000000100",
			281 => "0000000000010010001001",
			282 => "0000000000010010001001",
			283 => "0001000101101100001100",
			284 => "0011111000111000000100",
			285 => "0000000000010010001001",
			286 => "0011011100101000000100",
			287 => "0000000000010010001001",
			288 => "0000000000010010001001",
			289 => "0000000000010010001001",
			290 => "0001010110101100110100",
			291 => "0000110101101100011100",
			292 => "0001011110011000001100",
			293 => "0011111001001000000100",
			294 => "0000000000010100111101",
			295 => "0001001001100100000100",
			296 => "0000000000010100111101",
			297 => "0000000000010100111101",
			298 => "0010100110000000001100",
			299 => "0010000011001000000100",
			300 => "0000000000010100111101",
			301 => "0010000011100100000100",
			302 => "0000000000010100111101",
			303 => "0000000000010100111101",
			304 => "0000000000010100111101",
			305 => "0011110011010100010100",
			306 => "0000010111100100000100",
			307 => "0000000000010100111101",
			308 => "0011010101011100001000",
			309 => "0000101001111100000100",
			310 => "0000000000010100111101",
			311 => "0000000000010100111101",
			312 => "0000001001000000000100",
			313 => "0000000000010100111101",
			314 => "0000000000010100111101",
			315 => "0000000000010100111101",
			316 => "0011001001001000011000",
			317 => "0011111100001100000100",
			318 => "0000000000010100111101",
			319 => "0010000011010000001000",
			320 => "0000011001100100000100",
			321 => "0000000000010100111101",
			322 => "0000000000010100111101",
			323 => "0011010110110100000100",
			324 => "0000000000010100111101",
			325 => "0010110101011100000100",
			326 => "0000000000010100111101",
			327 => "0000000000010100111101",
			328 => "0010001001000100001000",
			329 => "0001011110010100000100",
			330 => "0000000000010100111101",
			331 => "0000000000010100111101",
			332 => "0001001101101000000100",
			333 => "0000000000010100111101",
			334 => "0000000000010100111101",
			335 => "0000010111100100110000",
			336 => "0011101111100000100000",
			337 => "0010110110001100000100",
			338 => "0000000000010111101001",
			339 => "0010001001000100010100",
			340 => "0001000101111000001100",
			341 => "0001011100000000001000",
			342 => "0001010011000000000100",
			343 => "0000000000010111101001",
			344 => "0000000000010111101001",
			345 => "0000000000010111101001",
			346 => "0011111101101100000100",
			347 => "0000000000010111101001",
			348 => "0000000000010111101001",
			349 => "0000001110010100000100",
			350 => "0000000000010111101001",
			351 => "0000000000010111101001",
			352 => "0000100100011100000100",
			353 => "0000000000010111101001",
			354 => "0001010001011000001000",
			355 => "0001101110111100000100",
			356 => "0000000000010111101001",
			357 => "0000000000010111101001",
			358 => "0000000000010111101001",
			359 => "0011101001000000011000",
			360 => "0010110011010000000100",
			361 => "0000000000010111101001",
			362 => "0010111010000100001100",
			363 => "0000000001101100001000",
			364 => "0000001011111000000100",
			365 => "0000000000010111101001",
			366 => "0000000000010111101001",
			367 => "0000000000010111101001",
			368 => "0010001111011000000100",
			369 => "0000000000010111101001",
			370 => "0000000000010111101001",
			371 => "0010010001010000001000",
			372 => "0010001001001100000100",
			373 => "0000000000010111101001",
			374 => "0000000000010111101001",
			375 => "0010100000111100000100",
			376 => "0000000000010111101001",
			377 => "0000000000010111101001",
			378 => "0000101110010001000100",
			379 => "0000110101101100100100",
			380 => "0001011110011000010100",
			381 => "0000011000111100000100",
			382 => "0000000000011001111101",
			383 => "0010100110110100001000",
			384 => "0001011000011000000100",
			385 => "0000000000011001111101",
			386 => "0000000000011001111101",
			387 => "0000001000101000000100",
			388 => "0000000000011001111101",
			389 => "0000000000011001111101",
			390 => "0010110101010100001000",
			391 => "0001011001001000000100",
			392 => "0000000000011001111101",
			393 => "0000000000011001111101",
			394 => "0010011000000000000100",
			395 => "0000000000011001111101",
			396 => "0000000000011001111101",
			397 => "0001000101101100001000",
			398 => "0000001011000000000100",
			399 => "0000000000011001111101",
			400 => "0000000000011001111101",
			401 => "0010110111011100001100",
			402 => "0011100001001000000100",
			403 => "0000000000011001111101",
			404 => "0011101001101100000100",
			405 => "0000000000011001111101",
			406 => "0000000000011001111101",
			407 => "0001111100010000001000",
			408 => "0011101100110100000100",
			409 => "0000000000011001111101",
			410 => "0000000000011001111101",
			411 => "0000000000011001111101",
			412 => "0010000011010000000100",
			413 => "0000000000011001111101",
			414 => "0000000000011001111101",
			415 => "0000010111100100111000",
			416 => "0011001010100100010100",
			417 => "0011011111011100001100",
			418 => "0010111101000000000100",
			419 => "0000000000011100100001",
			420 => "0000011001100100000100",
			421 => "0000000000011100100001",
			422 => "0000000000011100100001",
			423 => "0010000011010000000100",
			424 => "0000000000011100100001",
			425 => "0000000000011100100001",
			426 => "0001001011111000011100",
			427 => "0011110011010100011000",
			428 => "0010101001001100001100",
			429 => "0000001101000100001000",
			430 => "0000001000000100000100",
			431 => "0000000000011100100001",
			432 => "0000000000011100100001",
			433 => "0000000000011100100001",
			434 => "0010001001000100001000",
			435 => "0010010110000000000100",
			436 => "0000000000011100100001",
			437 => "0000000000011100100001",
			438 => "0000000000011100100001",
			439 => "0000000000011100100001",
			440 => "0000010110010000000100",
			441 => "0000000000011100100001",
			442 => "0000000000011100100001",
			443 => "0010010001010000010100",
			444 => "0010001001001100000100",
			445 => "0000000000011100100001",
			446 => "0001010001100100000100",
			447 => "0000000000011100100001",
			448 => "0001011100011100000100",
			449 => "0000000000011100100001",
			450 => "0001010011110100000100",
			451 => "0000000000011100100001",
			452 => "0000000000011100100001",
			453 => "0001001001001000000100",
			454 => "0000000000011100100001",
			455 => "0000000000011100100001",
			456 => "0011101010100001000000",
			457 => "0011000101010100100000",
			458 => "0001010110101100011000",
			459 => "0011001011101100000100",
			460 => "0000000000011111100101",
			461 => "0010000101101100010000",
			462 => "0011000011010000001000",
			463 => "0010101110011000000100",
			464 => "0000000000011111100101",
			465 => "0000001000011111100101",
			466 => "0000000110100000000100",
			467 => "0000000000011111100101",
			468 => "0000000000011111100101",
			469 => "0000000000011111100101",
			470 => "0011111111100100000100",
			471 => "0000000000011111100101",
			472 => "0000000000011111100101",
			473 => "0010001001000100010000",
			474 => "0011101100001100001000",
			475 => "0000001000101000000100",
			476 => "0000000000011111100101",
			477 => "0000001000011111100101",
			478 => "0011000101011100000100",
			479 => "0000000000011111100101",
			480 => "0000000000011111100101",
			481 => "0001000101101100001100",
			482 => "0000000001101100001000",
			483 => "0000001011000000000100",
			484 => "0000000000011111100101",
			485 => "0000000000011111100101",
			486 => "0000000000011111100101",
			487 => "0000000000011111100101",
			488 => "0010101000111000010000",
			489 => "0011000011010000001000",
			490 => "0011011101000000000100",
			491 => "0000000000011111100101",
			492 => "0000000000011111100101",
			493 => "0011110100001100000100",
			494 => "0000000000011111100101",
			495 => "0000000000011111100101",
			496 => "0010000011010000001000",
			497 => "0001010100101100000100",
			498 => "0000000000011111100101",
			499 => "0000000000011111100101",
			500 => "0011001001001000000100",
			501 => "1111111000011111100101",
			502 => "0000000100100000000100",
			503 => "0000000000011111100101",
			504 => "0000000000011111100101",
			505 => "0011100000100000110100",
			506 => "0001010110101100011000",
			507 => "0011000110110100000100",
			508 => "1111111000100001010001",
			509 => "0000101010000100000100",
			510 => "1111111000100001010001",
			511 => "0011100101111000000100",
			512 => "0000001000100001010001",
			513 => "0011001011101100000100",
			514 => "1111111000100001010001",
			515 => "0010101010100100000100",
			516 => "0000000000100001010001",
			517 => "0000000000100001010001",
			518 => "0010001001000100010100",
			519 => "0011001001001000010000",
			520 => "0010000011010000000100",
			521 => "0000001000100001010001",
			522 => "0000000001101100000100",
			523 => "0000000000100001010001",
			524 => "0000011000111100000100",
			525 => "0000000000100001010001",
			526 => "1111111000100001010001",
			527 => "0000001000100001010001",
			528 => "0001111011111000000100",
			529 => "1111111000100001010001",
			530 => "0000000000100001010001",
			531 => "1111111000100001010001",
			532 => "0001111000000100101100",
			533 => "0000101101000100011000",
			534 => "0010110110001100000100",
			535 => "1111111000100011101101",
			536 => "0000011000111100000100",
			537 => "0000010000100011101101",
			538 => "0011001010100100000100",
			539 => "0000000000100011101101",
			540 => "0010111010100100000100",
			541 => "0000001000100011101101",
			542 => "0001111111011000000100",
			543 => "0000001000100011101101",
			544 => "0000001000100011101101",
			545 => "0001001011101100000100",
			546 => "1111111000100011101101",
			547 => "0001011100000000001000",
			548 => "0011111101101100000100",
			549 => "0000000000100011101101",
			550 => "0000001000100011101101",
			551 => "0000001110100100000100",
			552 => "0000001000100011101101",
			553 => "1111111000100011101101",
			554 => "0000100111101000011100",
			555 => "0000001000101000000100",
			556 => "1111111000100011101101",
			557 => "0000111000100000010100",
			558 => "0011001001001000001100",
			559 => "0011011011101100000100",
			560 => "0000001000100011101101",
			561 => "0001100100000000000100",
			562 => "0000000000100011101101",
			563 => "1111111000100011101101",
			564 => "0010101101001000000100",
			565 => "0000000000100011101101",
			566 => "0000010000100011101101",
			567 => "1111111000100011101101",
			568 => "0010101010000100000100",
			569 => "0000000000100011101101",
			570 => "1111111000100011101101",
			571 => "0011101000100000011100",
			572 => "0010111010100100001100",
			573 => "0001100101111000000100",
			574 => "0000000000100110101001",
			575 => "0000000000111000000100",
			576 => "0000000000100110101001",
			577 => "0000000000100110101001",
			578 => "0001111111011000001000",
			579 => "0000000000110100000100",
			580 => "0000000000100110101001",
			581 => "0000000000100110101001",
			582 => "0001101100010000000100",
			583 => "0000000000100110101001",
			584 => "0000000000100110101001",
			585 => "0011001001001000110100",
			586 => "0010001001001100011000",
			587 => "0000111101101000001000",
			588 => "0001100010110000000100",
			589 => "0000000000100110101001",
			590 => "0000000000100110101001",
			591 => "0000010111100100001100",
			592 => "0011000111011100001000",
			593 => "0011000011010000000100",
			594 => "0000000000100110101001",
			595 => "0000000000100110101001",
			596 => "0000000000100110101001",
			597 => "0000000000100110101001",
			598 => "0010110101011100010000",
			599 => "0000000101000000000100",
			600 => "1111111000100110101001",
			601 => "0010001111111100001000",
			602 => "0000000100100000000100",
			603 => "0000000000100110101001",
			604 => "0000000000100110101001",
			605 => "0000000000100110101001",
			606 => "0011010111011100000100",
			607 => "0000000000100110101001",
			608 => "0011010101011100000100",
			609 => "0000000000100110101001",
			610 => "0000000000100110101001",
			611 => "0000010111100100001000",
			612 => "0001010010111000000100",
			613 => "0000000000100110101001",
			614 => "0000000000100110101001",
			615 => "0000100111100000000100",
			616 => "0000000000100110101001",
			617 => "0000000000100110101001",
			618 => "0001111000000001000000",
			619 => "0000000001101100101000",
			620 => "0010111010100100010000",
			621 => "0000000000111000001000",
			622 => "0010110110001100000100",
			623 => "1111111000101001100101",
			624 => "0000001000101001100101",
			625 => "0000010001110000000100",
			626 => "0000000000101001100101",
			627 => "1111111000101001100101",
			628 => "0000001000111000000100",
			629 => "1111111000101001100101",
			630 => "0010001001000100001000",
			631 => "0000001010001100000100",
			632 => "0000001000101001100101",
			633 => "0000001000101001100101",
			634 => "0000101001101100001000",
			635 => "0001101000111000000100",
			636 => "0000001000101001100101",
			637 => "0000001000101001100101",
			638 => "0000001000101001100101",
			639 => "0000010000011000001100",
			640 => "0000111001010100001000",
			641 => "0000101101010000000100",
			642 => "0000001000101001100101",
			643 => "1111111000101001100101",
			644 => "1111111000101001100101",
			645 => "0010100011000100001000",
			646 => "0011110000100000000100",
			647 => "1111111000101001100101",
			648 => "0000000000101001100101",
			649 => "0000000000101001100101",
			650 => "0000001100111000011100",
			651 => "0001101001011000001100",
			652 => "0001111000111000001000",
			653 => "0000000110001100000100",
			654 => "1111111000101001100101",
			655 => "0000000000101001100101",
			656 => "1111111000101001100101",
			657 => "0000110001001000001100",
			658 => "0001111100110000001000",
			659 => "0000011000011000000100",
			660 => "0000000000101001100101",
			661 => "1111111000101001100101",
			662 => "0000001000101001100101",
			663 => "1111111000101001100101",
			664 => "1111111000101001100101",
			665 => "0000101110010000110100",
			666 => "0011000110110100000100",
			667 => "0000000000101011110001",
			668 => "0010001001000100100000",
			669 => "0001011010011100011000",
			670 => "0001011111011000010000",
			671 => "0011000011010000001000",
			672 => "0001011100101000000100",
			673 => "0000000000101011110001",
			674 => "0000000000101011110001",
			675 => "0000001101000100000100",
			676 => "0000000000101011110001",
			677 => "0000000000101011110001",
			678 => "0011000011010000000100",
			679 => "0000000000101011110001",
			680 => "0000000000101011110001",
			681 => "0001001100101100000100",
			682 => "0000000000101011110001",
			683 => "0000000000101011110001",
			684 => "0001000101101100001100",
			685 => "0000100011000100000100",
			686 => "0000000000101011110001",
			687 => "0010010110000000000100",
			688 => "0000000000101011110001",
			689 => "0000000000101011110001",
			690 => "0000000000101011110001",
			691 => "0000010000011000010000",
			692 => "0010101000111000001000",
			693 => "0000100000001100000100",
			694 => "0000000000101011110001",
			695 => "0000000000101011110001",
			696 => "0010010011000000000100",
			697 => "0000000000101011110001",
			698 => "0000000000101011110001",
			699 => "0000000000101011110001",
			700 => "0001111000000100111000",
			701 => "0011111011111000011000",
			702 => "0010110110001100000100",
			703 => "1111111000101110010101",
			704 => "0001111111011000010000",
			705 => "0000001011111000000100",
			706 => "0000001000101110010101",
			707 => "0011111001010000001000",
			708 => "0000010011110000000100",
			709 => "0000001000101110010101",
			710 => "0000001000101110010101",
			711 => "0000001000101110010101",
			712 => "0000000000101110010101",
			713 => "0011000111011100010100",
			714 => "0000010000011000001100",
			715 => "0000001101010000001000",
			716 => "0001101001101100000100",
			717 => "0000000000101110010101",
			718 => "0000001000101110010101",
			719 => "1111111000101110010101",
			720 => "0010001001001100000100",
			721 => "0000000000101110010101",
			722 => "1111111000101110010101",
			723 => "0000101111110000000100",
			724 => "0000001000101110010101",
			725 => "0011101110001100000100",
			726 => "1111111000101110010101",
			727 => "0000001000101110010101",
			728 => "0000100000001100011000",
			729 => "0000001000101000000100",
			730 => "1111111000101110010101",
			731 => "0001001011111000010000",
			732 => "0011000011010000000100",
			733 => "1111111000101110010101",
			734 => "0000010111100100000100",
			735 => "0000001000101110010101",
			736 => "0001011011111000000100",
			737 => "0000000000101110010101",
			738 => "1111111000101110010101",
			739 => "1111111000101110010101",
			740 => "1111111000101110010101",
			741 => "0000100000001100111000",
			742 => "0001010110101100100000",
			743 => "0011000110110100000100",
			744 => "1111111000110000001001",
			745 => "0000101010000100000100",
			746 => "1111111000110000001001",
			747 => "0000100000111000001100",
			748 => "0010011100110000001000",
			749 => "0000010011110000000100",
			750 => "0000001000110000001001",
			751 => "0000000000110000001001",
			752 => "0000000000110000001001",
			753 => "0001111001000100000100",
			754 => "1111111000110000001001",
			755 => "0000000010000000000100",
			756 => "0000001000110000001001",
			757 => "0000000000110000001001",
			758 => "0010001001000100010000",
			759 => "0010110101011100001100",
			760 => "0001011010011100001000",
			761 => "0011000011010000000100",
			762 => "1111111000110000001001",
			763 => "0000000000110000001001",
			764 => "1111111000110000001001",
			765 => "0000001000110000001001",
			766 => "0001111101001000000100",
			767 => "1111111000110000001001",
			768 => "0000000000110000001001",
			769 => "1111111000110000001001",
			770 => "0011100000100000110000",
			771 => "0001011010011100101100",
			772 => "0010001001001100001100",
			773 => "0010110110001100000100",
			774 => "0000000000110001101101",
			775 => "0010101111011000000100",
			776 => "0000001000110001101101",
			777 => "0000000000110001101101",
			778 => "0011000011010000001000",
			779 => "0001101000000000000100",
			780 => "0000000000110001101101",
			781 => "1111111000110001101101",
			782 => "0001110101111000001100",
			783 => "0000101101000100001000",
			784 => "0010101111011100000100",
			785 => "0000000000110001101101",
			786 => "0000001000110001101101",
			787 => "0000000000110001101101",
			788 => "0001101000111000000100",
			789 => "1111111000110001101101",
			790 => "0010101000101000000100",
			791 => "0000000000110001101101",
			792 => "0000000000110001101101",
			793 => "1111111000110001101101",
			794 => "1111111000110001101101",
			795 => "0001001110011000100000",
			796 => "0010101010100100001100",
			797 => "0001011001100000001000",
			798 => "0000001010011100000100",
			799 => "0000000000110100101001",
			800 => "0000000000110100101001",
			801 => "0000000000110100101001",
			802 => "0001101101000100001100",
			803 => "0000000100110000001000",
			804 => "0000001011000000000100",
			805 => "0000000000110100101001",
			806 => "0000000000110100101001",
			807 => "0000000000110100101001",
			808 => "0010111110011000000100",
			809 => "0000000000110100101001",
			810 => "0000000000110100101001",
			811 => "0011000101010100001100",
			812 => "0001101111101000000100",
			813 => "0000000000110100101001",
			814 => "0010110111011100000100",
			815 => "0000000000110100101001",
			816 => "0000000000110100101001",
			817 => "0011011011101100001000",
			818 => "0001001011111000000100",
			819 => "0000000000110100101001",
			820 => "0000000000110100101001",
			821 => "0000101101100100010100",
			822 => "0010001001000100000100",
			823 => "0000000000110100101001",
			824 => "0001111011111000001000",
			825 => "0010101101001000000100",
			826 => "0000000000110100101001",
			827 => "0000000000110100101001",
			828 => "0000011110011000000100",
			829 => "0000000000110100101001",
			830 => "0000000000110100101001",
			831 => "0010010011001000001100",
			832 => "0001110110101100000100",
			833 => "0000000000110100101001",
			834 => "0001111101001000000100",
			835 => "0000000000110100101001",
			836 => "0000000000110100101001",
			837 => "0000010110010000000100",
			838 => "0000000000110100101001",
			839 => "0010001011000000000100",
			840 => "0000000000110100101001",
			841 => "0000000000110100101001",
			842 => "0001111100010001001000",
			843 => "0000000001101100101000",
			844 => "0000000011000000000100",
			845 => "1111111000110111100101",
			846 => "0011000111011100010100",
			847 => "0001100011001000001000",
			848 => "0000010001110000000100",
			849 => "0000001000110111100101",
			850 => "0000001000110111100101",
			851 => "0000010111100100001000",
			852 => "0000110101010100000100",
			853 => "1111111000110111100101",
			854 => "0000000000110111100101",
			855 => "1111111000110111100101",
			856 => "0010001111011000001100",
			857 => "0001011111011000001000",
			858 => "0010100110110100000100",
			859 => "0000001000110111100101",
			860 => "0000001000110111100101",
			861 => "0000001000110111100101",
			862 => "0000000000110111100101",
			863 => "0011011011101100010000",
			864 => "0000100000001100001100",
			865 => "0001100010001100000100",
			866 => "1111111000110111100101",
			867 => "0001001111101000000100",
			868 => "0000001000110111100101",
			869 => "1111111000110111100101",
			870 => "1111111000110111100101",
			871 => "0011001001001000001000",
			872 => "0010011001001000000100",
			873 => "0000000000110111100101",
			874 => "1111111000110111100101",
			875 => "0001001001000100000100",
			876 => "1111111000110111100101",
			877 => "0000000000110111100101",
			878 => "0011001101001000010100",
			879 => "0011101111100100010000",
			880 => "0010000101101100001000",
			881 => "0011001001001000000100",
			882 => "1111111000110111100101",
			883 => "0000001000110111100101",
			884 => "0011010101111000000100",
			885 => "1111111000110111100101",
			886 => "0000000000110111100101",
			887 => "1111111000110111100101",
			888 => "0000000000110111100101",
			889 => "0000100000001100110100",
			890 => "0001011010011100110000",
			891 => "0010001001001100001100",
			892 => "0010010101010100000100",
			893 => "0000000000111001010001",
			894 => "0001101100110100000100",
			895 => "0000000000111001010001",
			896 => "0000001000111001010001",
			897 => "0011000011010000001100",
			898 => "0001101000000000000100",
			899 => "0000000000111001010001",
			900 => "0000000110000100000100",
			901 => "1111111000111001010001",
			902 => "0000000000111001010001",
			903 => "0001110101111000001100",
			904 => "0000101101000100001000",
			905 => "0010101111011100000100",
			906 => "0000000000111001010001",
			907 => "0000001000111001010001",
			908 => "0000000000111001010001",
			909 => "0001101000111000000100",
			910 => "1111111000111001010001",
			911 => "0010101000101000000100",
			912 => "0000000000111001010001",
			913 => "0000000000111001010001",
			914 => "1111111000111001010001",
			915 => "1111111000111001010001",
			916 => "0011101010110100111100",
			917 => "0011000110110100000100",
			918 => "0000000000111011010101",
			919 => "0001010110101100011100",
			920 => "0001111000000100010000",
			921 => "0011001011101100000100",
			922 => "0000000000111011010101",
			923 => "0001001001100100000100",
			924 => "0000000000111011010101",
			925 => "0010010110000000000100",
			926 => "0000000000111011010101",
			927 => "0000000000111011010101",
			928 => "0001101010100000001000",
			929 => "0010101000011000000100",
			930 => "0000000000111011010101",
			931 => "0000000000111011010101",
			932 => "0000000000111011010101",
			933 => "0011001001001000010000",
			934 => "0011111100001100000100",
			935 => "0000000000111011010101",
			936 => "0010000011010000000100",
			937 => "0000000000111011010101",
			938 => "0010110101011100000100",
			939 => "0000000000111011010101",
			940 => "0000000000111011010101",
			941 => "0011010111011100000100",
			942 => "0000000000111011010101",
			943 => "0000010110110100000100",
			944 => "0000000000111011010101",
			945 => "0000000000111011010101",
			946 => "0001111000000000000100",
			947 => "0000000000111011010101",
			948 => "0000000000111011010101",
			949 => "0000100000001101000100",
			950 => "0001000011110000010000",
			951 => "0000000011000000000100",
			952 => "0000000000111101100001",
			953 => "0000101101101100000100",
			954 => "0000001000111101100001",
			955 => "0001101100110100000100",
			956 => "0000000000111101100001",
			957 => "0000000000111101100001",
			958 => "0000011000011000011000",
			959 => "0011001011101100000100",
			960 => "1111111000111101100001",
			961 => "0001011010011100001100",
			962 => "0010101001010100001000",
			963 => "0010010110000000000100",
			964 => "0000000000111101100001",
			965 => "0000000000111101100001",
			966 => "0000001000111101100001",
			967 => "0010010011000000000100",
			968 => "1111111000111101100001",
			969 => "0000000000111101100001",
			970 => "0001000101101100010100",
			971 => "0010100011001000001100",
			972 => "0001010011010000001000",
			973 => "0001111000111000000100",
			974 => "0000000000111101100001",
			975 => "0000000000111101100001",
			976 => "1111111000111101100001",
			977 => "0010010011001000000100",
			978 => "0000000000111101100001",
			979 => "0000001000111101100001",
			980 => "0011011010100100000100",
			981 => "0000000000111101100001",
			982 => "1111111000111101100001",
			983 => "1111111000111101100001",
			984 => "0011100000100000110100",
			985 => "0001011010011100101100",
			986 => "0010110110001100000100",
			987 => "1111111000111111001101",
			988 => "0010001001001100001100",
			989 => "0001101111100000001000",
			990 => "0000001010100000000100",
			991 => "0000001000111111001101",
			992 => "0000000000111111001101",
			993 => "0000001000111111001101",
			994 => "0011000011010000001100",
			995 => "0001100001010000000100",
			996 => "0000000000111111001101",
			997 => "0001110101111000000100",
			998 => "1111111000111111001101",
			999 => "0000000000111111001101",
			1000 => "0001110101111000001000",
			1001 => "0000101101000100000100",
			1002 => "0000001000111111001101",
			1003 => "0000000000111111001101",
			1004 => "0001010001001000000100",
			1005 => "0000000000111111001101",
			1006 => "0000000000111111001101",
			1007 => "0010010011001000000100",
			1008 => "1111111000111111001101",
			1009 => "0000000000111111001101",
			1010 => "1111111000111111001101",
			1011 => "0000100101001101001000",
			1012 => "0001111000000100101100",
			1013 => "0011000101010100100000",
			1014 => "0000010111100100011000",
			1015 => "0000101101000100001100",
			1016 => "0010110110001100000100",
			1017 => "1111111001000001100001",
			1018 => "0000000001101000000100",
			1019 => "0000001001000001100001",
			1020 => "0000001001000001100001",
			1021 => "0001101001101100000100",
			1022 => "1111111001000001100001",
			1023 => "0000111001010000000100",
			1024 => "0000001001000001100001",
			1025 => "1111111001000001100001",
			1026 => "0001000110001100000100",
			1027 => "0000000001000001100001",
			1028 => "1111111001000001100001",
			1029 => "0000101111110000001000",
			1030 => "0010100110001100000100",
			1031 => "0000000001000001100001",
			1032 => "0000001001000001100001",
			1033 => "0000000001000001100001",
			1034 => "0000001000101000000100",
			1035 => "1111111001000001100001",
			1036 => "0010110101011100001100",
			1037 => "0010000101011100000100",
			1038 => "0000000001000001100001",
			1039 => "0001011000111000000100",
			1040 => "0000000001000001100001",
			1041 => "1111111001000001100001",
			1042 => "0000110001001000001000",
			1043 => "0000100111100000000100",
			1044 => "0000001001000001100001",
			1045 => "0000000001000001100001",
			1046 => "1111111001000001100001",
			1047 => "1111111001000001100001",
			1048 => "0011100000100001000000",
			1049 => "0010001001000100100000",
			1050 => "0001010000111000011100",
			1051 => "0010101011000000010100",
			1052 => "0011000110110100000100",
			1053 => "0000000001000011100101",
			1054 => "0001010110101100001000",
			1055 => "0011110101110000000100",
			1056 => "0000000001000011100101",
			1057 => "0000001001000011100101",
			1058 => "0011000011010000000100",
			1059 => "0000000001000011100101",
			1060 => "0000000001000011100101",
			1061 => "0010110111011100000100",
			1062 => "0000000001000011100101",
			1063 => "0000001001000011100101",
			1064 => "0000000001000011100101",
			1065 => "0001000101101100011100",
			1066 => "0010111001001000010000",
			1067 => "0001101111101000001100",
			1068 => "0000100110011100001000",
			1069 => "0010101111011100000100",
			1070 => "0000000001000011100101",
			1071 => "0000000001000011100101",
			1072 => "0000000001000011100101",
			1073 => "0000000001000011100101",
			1074 => "0000001001011000000100",
			1075 => "0000000001000011100101",
			1076 => "0000000100110000000100",
			1077 => "0000001001000011100101",
			1078 => "0000000001000011100101",
			1079 => "1111111001000011100101",
			1080 => "1111111001000011100101",
			1081 => "0000011000111100010100",
			1082 => "0001011010000100001000",
			1083 => "0010011100101000000100",
			1084 => "0000000001000110101001",
			1085 => "0000000001000110101001",
			1086 => "0000111111011000000100",
			1087 => "0000000001000110101001",
			1088 => "0001111000111000000100",
			1089 => "0000000001000110101001",
			1090 => "0000000001000110101001",
			1091 => "0011000111011100010000",
			1092 => "0001010001100100000100",
			1093 => "0000000001000110101001",
			1094 => "0010110111011100001000",
			1095 => "0010010110000000000100",
			1096 => "0000000001000110101001",
			1097 => "0000000001000110101001",
			1098 => "0000000001000110101001",
			1099 => "0001011010011100110100",
			1100 => "0010101000000000011100",
			1101 => "0001111000000100010000",
			1102 => "0000000110100000001000",
			1103 => "0011101010000100000100",
			1104 => "0000000001000110101001",
			1105 => "0000000001000110101001",
			1106 => "0011111010011100000100",
			1107 => "0000000001000110101001",
			1108 => "0000000001000110101001",
			1109 => "0000011110011000001000",
			1110 => "0001011111011100000100",
			1111 => "0000000001000110101001",
			1112 => "0000000001000110101001",
			1113 => "0000000001000110101001",
			1114 => "0010000101101100001000",
			1115 => "0000001100111000000100",
			1116 => "0000000001000110101001",
			1117 => "0000000001000110101001",
			1118 => "0011001010000100001000",
			1119 => "0000111000000000000100",
			1120 => "0000000001000110101001",
			1121 => "0000000001000110101001",
			1122 => "0010100000111100000100",
			1123 => "0000000001000110101001",
			1124 => "0000000001000110101001",
			1125 => "0010111100101000000100",
			1126 => "0000000001000110101001",
			1127 => "0000111000100000000100",
			1128 => "0000000001000110101001",
			1129 => "0000000001000110101001",
			1130 => "0000100000001100111000",
			1131 => "0000101010000100000100",
			1132 => "1111111001001000011101",
			1133 => "0001000101101100011000",
			1134 => "0011000110110100000100",
			1135 => "1111111001001000011101",
			1136 => "0001101111000100010000",
			1137 => "0000101111100000001000",
			1138 => "0010011100110000000100",
			1139 => "0000001001001000011101",
			1140 => "1111111001001000011101",
			1141 => "0010101010100100000100",
			1142 => "1111111001001000011101",
			1143 => "0000001001001000011101",
			1144 => "1111111001001000011101",
			1145 => "0010001001000100010100",
			1146 => "0011001100101000001100",
			1147 => "0001011010011100001000",
			1148 => "0011000011010000000100",
			1149 => "0000000001001000011101",
			1150 => "0000000001001000011101",
			1151 => "1111111001001000011101",
			1152 => "0001010010111000000100",
			1153 => "0000001001001000011101",
			1154 => "1111111001001000011101",
			1155 => "0010010011001000000100",
			1156 => "1111111001001000011101",
			1157 => "1111111001001000011101",
			1158 => "1111111001001000011101",
			1159 => "0011100000100001001000",
			1160 => "0011001001001000101000",
			1161 => "0001010011110100100100",
			1162 => "0010001111111100010100",
			1163 => "0011000110110100000100",
			1164 => "0000000001001010110001",
			1165 => "0011110111010100001000",
			1166 => "0000000000110100000100",
			1167 => "0000000001001010110001",
			1168 => "0000000001001010110001",
			1169 => "0000000000000100000100",
			1170 => "0000000001001010110001",
			1171 => "0000000001001010110001",
			1172 => "0011101010011100001100",
			1173 => "0011000011010000000100",
			1174 => "0000000001001010110001",
			1175 => "0000001000111000000100",
			1176 => "0000000001001010110001",
			1177 => "0000000001001010110001",
			1178 => "0000000001001010110001",
			1179 => "0000000001001010110001",
			1180 => "0000010111100100010000",
			1181 => "0010101000000000001100",
			1182 => "0011000101101100001000",
			1183 => "0000111101000000000100",
			1184 => "0000000001001010110001",
			1185 => "0000000001001010110001",
			1186 => "0000000001001010110001",
			1187 => "0000000001001010110001",
			1188 => "0000000010110100001100",
			1189 => "0001101000111000001000",
			1190 => "0001111111011000000100",
			1191 => "0000000001001010110001",
			1192 => "0000000001001010110001",
			1193 => "0000000001001010110001",
			1194 => "0000000001001010110001",
			1195 => "0000000001001010110001",
			1196 => "0011110010000001000100",
			1197 => "0001011010011100111100",
			1198 => "0000110101101100100000",
			1199 => "0001011110011000010100",
			1200 => "0000011000111100000100",
			1201 => "0000000001001100111101",
			1202 => "0010100110110100001000",
			1203 => "0001011000011000000100",
			1204 => "0000000001001100111101",
			1205 => "0000000001001100111101",
			1206 => "0000100110100000000100",
			1207 => "0000000001001100111101",
			1208 => "0000000001001100111101",
			1209 => "0001011001001000000100",
			1210 => "0000000001001100111101",
			1211 => "0001010101101100000100",
			1212 => "0000000001001100111101",
			1213 => "0000000001001100111101",
			1214 => "0001000101101100001100",
			1215 => "0000001000100000000100",
			1216 => "0000000001001100111101",
			1217 => "0001011000000100000100",
			1218 => "0000000001001100111101",
			1219 => "0000000001001100111101",
			1220 => "0010000101101100001100",
			1221 => "0010011001000100001000",
			1222 => "0000000010110100000100",
			1223 => "0000000001001100111101",
			1224 => "0000000001001100111101",
			1225 => "0000000001001100111101",
			1226 => "0000000001001100111101",
			1227 => "0010111100101000000100",
			1228 => "0000000001001100111101",
			1229 => "0000000001001100111101",
			1230 => "0000000001001100111101",
			1231 => "0000001100111000111100",
			1232 => "0000101010000100000100",
			1233 => "1111111001001111000001",
			1234 => "0000001001111100011000",
			1235 => "0010110110001100000100",
			1236 => "1111111001001111000001",
			1237 => "0000011101000000001100",
			1238 => "0000011001100100000100",
			1239 => "0000001001001111000001",
			1240 => "0000010011110000000100",
			1241 => "0000001001001111000001",
			1242 => "0000001001001111000001",
			1243 => "0001000101010100000100",
			1244 => "0000001001001111000001",
			1245 => "1111111001001111000001",
			1246 => "0010000011010000000100",
			1247 => "0000001001001111000001",
			1248 => "0011001100101000010000",
			1249 => "0000010000011000001000",
			1250 => "0001110011001000000100",
			1251 => "0000000001001111000001",
			1252 => "0000000001001111000001",
			1253 => "0011100011000100000100",
			1254 => "0000000001001111000001",
			1255 => "1111111001001111000001",
			1256 => "0000110001001000001000",
			1257 => "0010101111011000000100",
			1258 => "0000000001001111000001",
			1259 => "0000001001001111000001",
			1260 => "1111111001001111000001",
			1261 => "0001010101101100000100",
			1262 => "0000000001001111000001",
			1263 => "1111111001001111000001",
			1264 => "0011100000100001001100",
			1265 => "0010001111111100100000",
			1266 => "0001011010011100011100",
			1267 => "0011000110110100000100",
			1268 => "1111111001010001011101",
			1269 => "0011110001010100010000",
			1270 => "0000100000111000001000",
			1271 => "0000000011000000000100",
			1272 => "0000000001010001011101",
			1273 => "0000001001010001011101",
			1274 => "0000111101101000000100",
			1275 => "1111111001010001011101",
			1276 => "0000000001010001011101",
			1277 => "0010111011101100000100",
			1278 => "0000000001010001011101",
			1279 => "0000001001010001011101",
			1280 => "1111111001010001011101",
			1281 => "0010110101011100010000",
			1282 => "0011100011000100001100",
			1283 => "0010111010100100000100",
			1284 => "1111111001010001011101",
			1285 => "0000001000111000000100",
			1286 => "0000000001010001011101",
			1287 => "0000001001010001011101",
			1288 => "1111111001010001011101",
			1289 => "0000010111110000001000",
			1290 => "0000111100101000000100",
			1291 => "0000000001010001011101",
			1292 => "0000001001010001011101",
			1293 => "0001000110000000001100",
			1294 => "0000001011111000000100",
			1295 => "0000000001010001011101",
			1296 => "0000000010110100000100",
			1297 => "0000001001010001011101",
			1298 => "0000000001010001011101",
			1299 => "0010100100101100000100",
			1300 => "0000000001010001011101",
			1301 => "1111111001010001011101",
			1302 => "1111111001010001011101",
			1303 => "0011110110100001001000",
			1304 => "0011001011101100001000",
			1305 => "0011111000000100000100",
			1306 => "0000000001010011110001",
			1307 => "0000000001010011110001",
			1308 => "0001011100000000011100",
			1309 => "0010101010100100001100",
			1310 => "0000001010100000001000",
			1311 => "0000001000000100000100",
			1312 => "0000000001010011110001",
			1313 => "0000000001010011110001",
			1314 => "0000000001010011110001",
			1315 => "0001000101101100001100",
			1316 => "0000001011000000000100",
			1317 => "0000000001010011110001",
			1318 => "0000001000110100000100",
			1319 => "0000000001010011110001",
			1320 => "0000000001010011110001",
			1321 => "0000000001010011110001",
			1322 => "0011000101011100010000",
			1323 => "0001100000100000001100",
			1324 => "0000010001110000001000",
			1325 => "0011100001111100000100",
			1326 => "0000000001010011110001",
			1327 => "0000000001010011110001",
			1328 => "0000000001010011110001",
			1329 => "0000000001010011110001",
			1330 => "0010001001000100001100",
			1331 => "0001000011000100001000",
			1332 => "0010101111101000000100",
			1333 => "0000000001010011110001",
			1334 => "0000000001010011110001",
			1335 => "0000000001010011110001",
			1336 => "0010011001010000000100",
			1337 => "0000000001010011110001",
			1338 => "0000000001010011110001",
			1339 => "0000000001010011110001",
			1340 => "0000100000001101001000",
			1341 => "0001011010011101000000",
			1342 => "0000110101101100100000",
			1343 => "0001011110011000010000",
			1344 => "0010111101000000000100",
			1345 => "0000000001010110000101",
			1346 => "0011000111011100000100",
			1347 => "0000000001010110000101",
			1348 => "0011011011101100000100",
			1349 => "0000000001010110000101",
			1350 => "0000000001010110000101",
			1351 => "0010001111011000000100",
			1352 => "0000000001010110000101",
			1353 => "0011010101101100000100",
			1354 => "0000000001010110000101",
			1355 => "0010000011100100000100",
			1356 => "0000000001010110000101",
			1357 => "0000000001010110000101",
			1358 => "0000010111100100001100",
			1359 => "0010000101101100001000",
			1360 => "0001100010001000000100",
			1361 => "0000000001010110000101",
			1362 => "0000000001010110000101",
			1363 => "0000000001010110000101",
			1364 => "0011000101010100000100",
			1365 => "0000000001010110000101",
			1366 => "0000001100110100001000",
			1367 => "0010111010000100000100",
			1368 => "0000000001010110000101",
			1369 => "0000000001010110000101",
			1370 => "0000000011011000000100",
			1371 => "0000000001010110000101",
			1372 => "0000000001010110000101",
			1373 => "0011001001001000000100",
			1374 => "0000000001010110000101",
			1375 => "0000000001010110000101",
			1376 => "0000000001010110000101",
			1377 => "0011100000100001010000",
			1378 => "0001000101101100111000",
			1379 => "0000110101101100100100",
			1380 => "0001000011110000010000",
			1381 => "0000000011000000000100",
			1382 => "0000000001011000101001",
			1383 => "0000001010100000000100",
			1384 => "0000001001011000101001",
			1385 => "0001110101111000000100",
			1386 => "1111111001011000101001",
			1387 => "0000000001011000101001",
			1388 => "0010100101101100010000",
			1389 => "0001010110001100001000",
			1390 => "0000111101000000000100",
			1391 => "0000000001011000101001",
			1392 => "0000000001011000101001",
			1393 => "0000111100101000000100",
			1394 => "1111111001011000101001",
			1395 => "0000000001011000101001",
			1396 => "0000000001011000101001",
			1397 => "0000010111100100000100",
			1398 => "0000001001011000101001",
			1399 => "0000000010110100001100",
			1400 => "0010011010000100000100",
			1401 => "0000000001011000101001",
			1402 => "0000001001000000000100",
			1403 => "0000000001011000101001",
			1404 => "0000001001011000101001",
			1405 => "0000000001011000101001",
			1406 => "0010001001000100010100",
			1407 => "0001101010011100000100",
			1408 => "0000000001011000101001",
			1409 => "0011001001001000001100",
			1410 => "0010000011010000000100",
			1411 => "0000000001011000101001",
			1412 => "0001011001011000000100",
			1413 => "0000000001011000101001",
			1414 => "1111111001011000101001",
			1415 => "0000000001011000101001",
			1416 => "1111111001011000101001",
			1417 => "1111111001011000101001",
			1418 => "0011100000100001100100",
			1419 => "0001001110011000110000",
			1420 => "0000111100101000100100",
			1421 => "0001001001100000010000",
			1422 => "0010001001001100000100",
			1423 => "0000001001011011110111",
			1424 => "0011011011101100000100",
			1425 => "0000000001011011110111",
			1426 => "0000100110100000000100",
			1427 => "0000000001011011110111",
			1428 => "0000000001011011110111",
			1429 => "0001011001001000001100",
			1430 => "0000000001011100001000",
			1431 => "0000001011000000000100",
			1432 => "0000000001011011110111",
			1433 => "0000000001011011110111",
			1434 => "1111111001011011110111",
			1435 => "0001111001010100000100",
			1436 => "0000000001011011110111",
			1437 => "0000000001011011110111",
			1438 => "0000010111100100000100",
			1439 => "0000001001011011110111",
			1440 => "0011010101010100000100",
			1441 => "0000000001011011110111",
			1442 => "0000000001011011110111",
			1443 => "0000010111100100011100",
			1444 => "0011001001001000010100",
			1445 => "0000000110100000000100",
			1446 => "0000000001011011110111",
			1447 => "0011110101001000001000",
			1448 => "0010101111101000000100",
			1449 => "1111111001011011110111",
			1450 => "0000000001011011110111",
			1451 => "0010001111111100000100",
			1452 => "0000000001011011110111",
			1453 => "0000000001011011110111",
			1454 => "0000101110010000000100",
			1455 => "0000001001011011110111",
			1456 => "0000000001011011110111",
			1457 => "0010111000000000010100",
			1458 => "0010001111111100000100",
			1459 => "0000000001011011110111",
			1460 => "0001000101011100001000",
			1461 => "0010100110000000000100",
			1462 => "0000000001011011110111",
			1463 => "0000000001011011110111",
			1464 => "0010101000000000000100",
			1465 => "0000000001011011110111",
			1466 => "1111111001011011110111",
			1467 => "0000000001011011110111",
			1468 => "1111111001011011110111",
			1469 => "0000000001101100011000",
			1470 => "0010111010100100001100",
			1471 => "0000011000111100000100",
			1472 => "0000000001011101101001",
			1473 => "0011100011001000000100",
			1474 => "0000000001011101101001",
			1475 => "0000000001011101101001",
			1476 => "0001101000111000001000",
			1477 => "0001111111011000000100",
			1478 => "0000000001011101101001",
			1479 => "0000000001011101101001",
			1480 => "0000000001011101101001",
			1481 => "0011011011101100010100",
			1482 => "0001100010001100000100",
			1483 => "0000000001011101101001",
			1484 => "0010010111011100000100",
			1485 => "0000000001011101101001",
			1486 => "0011110010000000001000",
			1487 => "0001001111101000000100",
			1488 => "0000000001011101101001",
			1489 => "0000000001011101101001",
			1490 => "0000000001011101101001",
			1491 => "0011001001001000001000",
			1492 => "0000011000111100000100",
			1493 => "0000000001011101101001",
			1494 => "0000000001011101101001",
			1495 => "0000101110010000000100",
			1496 => "0000000001011101101001",
			1497 => "0000000001011101101001",
			1498 => "0001010110101100100000",
			1499 => "0000000000110100001100",
			1500 => "0010110110001100000100",
			1501 => "0000000001011111100101",
			1502 => "0000101010000100000100",
			1503 => "0000000001011111100101",
			1504 => "0000000001011111100101",
			1505 => "0011110101110000000100",
			1506 => "0000000001011111100101",
			1507 => "0010010111011100000100",
			1508 => "0000000001011111100101",
			1509 => "0011110011010100001000",
			1510 => "0010001111111100000100",
			1511 => "0000000001011111100101",
			1512 => "0000000001011111100101",
			1513 => "0000000001011111100101",
			1514 => "0011001001001000010000",
			1515 => "0011100001011000000100",
			1516 => "0000000001011111100101",
			1517 => "0010000011010000000100",
			1518 => "0000000001011111100101",
			1519 => "0000011000111100000100",
			1520 => "0000000001011111100101",
			1521 => "0000000001011111100101",
			1522 => "0010001001000100001000",
			1523 => "0001001001011000000100",
			1524 => "0000000001011111100101",
			1525 => "0000000001011111100101",
			1526 => "0001001010000100000100",
			1527 => "0000000001011111100101",
			1528 => "0000000001011111100101",
			1529 => "0011001001001000110100",
			1530 => "0011100001001000010100",
			1531 => "0010111010100100001100",
			1532 => "0011111010000100000100",
			1533 => "0000000001100001110001",
			1534 => "0000110101101100000100",
			1535 => "0000000001100001110001",
			1536 => "0000000001100001110001",
			1537 => "0000001000111000000100",
			1538 => "0000000001100001110001",
			1539 => "0000000001100001110001",
			1540 => "0010000011010000001100",
			1541 => "0011011101000000000100",
			1542 => "0000000001100001110001",
			1543 => "0000001101010000000100",
			1544 => "0000000001100001110001",
			1545 => "0000000001100001110001",
			1546 => "0000011000111100001100",
			1547 => "0010011001000100001000",
			1548 => "0011010110110100000100",
			1549 => "0000000001100001110001",
			1550 => "0000000001100001110001",
			1551 => "0000000001100001110001",
			1552 => "0011011101000000000100",
			1553 => "0000000001100001110001",
			1554 => "0000000001100001110001",
			1555 => "0000101110010000001100",
			1556 => "0001101000111000001000",
			1557 => "0001111111011000000100",
			1558 => "0000000001100001110001",
			1559 => "0000000001100001110001",
			1560 => "0000000001100001110001",
			1561 => "0000010001110000000100",
			1562 => "0000000001100001110001",
			1563 => "0000000001100001110001",
			1564 => "0001111000000100101100",
			1565 => "0000101101000100011000",
			1566 => "0011001110011000001000",
			1567 => "0011011111011100000100",
			1568 => "0000000001100100000101",
			1569 => "1111111001100100000101",
			1570 => "0001011001010100001100",
			1571 => "0001100001010000001000",
			1572 => "0011111001010000000100",
			1573 => "0000011001100100000101",
			1574 => "0000011001100100000101",
			1575 => "0000100001100100000101",
			1576 => "0000010001100100000101",
			1577 => "0000010000011000001000",
			1578 => "0010101000000000000100",
			1579 => "0000010001100100000101",
			1580 => "1111111001100100000101",
			1581 => "0011111011110000001000",
			1582 => "0010011101101000000100",
			1583 => "1111111001100100000101",
			1584 => "0000000001100100000101",
			1585 => "0000000001100100000101",
			1586 => "0000100111101000011000",
			1587 => "0000001000101000000100",
			1588 => "1111111001100100000101",
			1589 => "0000101101100100001000",
			1590 => "0011001001001000000100",
			1591 => "0000001001100100000101",
			1592 => "0000011001100100000101",
			1593 => "0010001111111100000100",
			1594 => "0000001001100100000101",
			1595 => "0011001001001000000100",
			1596 => "1111111001100100000101",
			1597 => "0000000001100100000101",
			1598 => "0001010101101100000100",
			1599 => "0000000001100100000101",
			1600 => "1111111001100100000101",
			1601 => "0001111000000100101000",
			1602 => "0000101101000100010100",
			1603 => "0010110110001100000100",
			1604 => "1111111001100110010001",
			1605 => "0001011001010100001100",
			1606 => "0011001010100100000100",
			1607 => "0000001001100110010001",
			1608 => "0011101001010100000100",
			1609 => "0000010001100110010001",
			1610 => "0000010001100110010001",
			1611 => "0000000001100110010001",
			1612 => "0000010000011000001000",
			1613 => "0001110011000000000100",
			1614 => "1111111001100110010001",
			1615 => "0000001001100110010001",
			1616 => "0000101111110000000100",
			1617 => "0000001001100110010001",
			1618 => "0001101101101100000100",
			1619 => "1111111001100110010001",
			1620 => "0000000001100110010001",
			1621 => "0000100111101000011000",
			1622 => "0000001000101000000100",
			1623 => "1111111001100110010001",
			1624 => "0010100000111100010000",
			1625 => "0010010011001000001100",
			1626 => "0011000011010000000100",
			1627 => "1111111001100110010001",
			1628 => "0010000101101100000100",
			1629 => "0000010001100110010001",
			1630 => "0000000001100110010001",
			1631 => "0000010001100110010001",
			1632 => "1111111001100110010001",
			1633 => "0001010101101100000100",
			1634 => "0000000001100110010001",
			1635 => "1111111001100110010001",
			1636 => "0010001111111100101000",
			1637 => "0010110110001100001000",
			1638 => "0000000101000000000100",
			1639 => "0000000001101000100101",
			1640 => "0000000001101000100101",
			1641 => "0001011010011100011000",
			1642 => "0011110011010100010100",
			1643 => "0011110111010100010000",
			1644 => "0011110100101100001000",
			1645 => "0000000011000000000100",
			1646 => "0000000001101000100101",
			1647 => "0000000001101000100101",
			1648 => "0000010111110000000100",
			1649 => "0000000001101000100101",
			1650 => "0000000001101000100101",
			1651 => "0000000001101000100101",
			1652 => "0000000001101000100101",
			1653 => "0011100010001100000100",
			1654 => "0000000001101000100101",
			1655 => "0000000001101000100101",
			1656 => "0010110101011100010000",
			1657 => "0011101001011000001000",
			1658 => "0010101010000100000100",
			1659 => "0000000001101000100101",
			1660 => "0000000001101000100101",
			1661 => "0001000110001100000100",
			1662 => "0000000001101000100101",
			1663 => "0000000001101000100101",
			1664 => "0000101110010000010000",
			1665 => "0001101000111000001000",
			1666 => "0001111111011000000100",
			1667 => "0000000001101000100101",
			1668 => "0000000001101000100101",
			1669 => "0000110111011100000100",
			1670 => "0000000001101000100101",
			1671 => "0000000001101000100101",
			1672 => "0000000001101000100101",
			1673 => "0011001001001001000000",
			1674 => "0011100001001000011000",
			1675 => "0010111010100100010000",
			1676 => "0000000000111000001000",
			1677 => "0010110110001100000100",
			1678 => "0000000001101011001001",
			1679 => "0000000001101011001001",
			1680 => "0000110101101100000100",
			1681 => "0000000001101011001001",
			1682 => "0000000001101011001001",
			1683 => "0000001000111000000100",
			1684 => "0000000001101011001001",
			1685 => "0000000001101011001001",
			1686 => "0010000011010000001100",
			1687 => "0011011101000000000100",
			1688 => "0000000001101011001001",
			1689 => "0001111100010000000100",
			1690 => "0000000001101011001001",
			1691 => "0000000001101011001001",
			1692 => "0000011000111100001100",
			1693 => "0010111110011000000100",
			1694 => "0000000001101011001001",
			1695 => "0010110011010000000100",
			1696 => "0000000001101011001001",
			1697 => "0000000001101011001001",
			1698 => "0010110101011100001000",
			1699 => "0011011101000000000100",
			1700 => "0000000001101011001001",
			1701 => "0000000001101011001001",
			1702 => "0011011010100100000100",
			1703 => "0000000001101011001001",
			1704 => "0000000001101011001001",
			1705 => "0000101110010000001100",
			1706 => "0001101000111000001000",
			1707 => "0001111111011000000100",
			1708 => "0000000001101011001001",
			1709 => "0000000001101011001001",
			1710 => "0000000001101011001001",
			1711 => "0000010001110000000100",
			1712 => "0000000001101011001001",
			1713 => "0000000001101011001001",
			1714 => "0001111000000100101100",
			1715 => "0000101101101100010000",
			1716 => "0010110110001100000100",
			1717 => "1111111001101101011101",
			1718 => "0000011101000000001000",
			1719 => "0000011000111100000100",
			1720 => "0000011001101101011101",
			1721 => "0000010001101101011101",
			1722 => "0000001001101101011101",
			1723 => "0000011000011000010100",
			1724 => "0000100101001100010000",
			1725 => "0010101010100100000100",
			1726 => "1111111001101101011101",
			1727 => "0001010001011000001000",
			1728 => "0001110011000000000100",
			1729 => "0000001001101101011101",
			1730 => "0000011001101101011101",
			1731 => "1111111001101101011101",
			1732 => "1111111001101101011101",
			1733 => "0010110101010100000100",
			1734 => "1111111001101101011101",
			1735 => "0000000001101101011101",
			1736 => "0000100111101000011000",
			1737 => "0000001000101000000100",
			1738 => "1111111001101101011101",
			1739 => "0010100000111100010000",
			1740 => "0000100010110000000100",
			1741 => "0000010001101101011101",
			1742 => "0010001111111100000100",
			1743 => "0000010001101101011101",
			1744 => "0011100101110000000100",
			1745 => "1111111001101101011101",
			1746 => "0000001001101101011101",
			1747 => "1111111001101101011101",
			1748 => "0001010101101100000100",
			1749 => "0000000001101101011101",
			1750 => "1111111001101101011101",
			1751 => "0001011110011000001100",
			1752 => "0010111101000000000100",
			1753 => "0000000001101111101001",
			1754 => "0000000011000000000100",
			1755 => "0000000001101111101001",
			1756 => "0000000001101111101001",
			1757 => "0011000011010000010100",
			1758 => "0010000011010000001100",
			1759 => "0011001011101100000100",
			1760 => "0000000001101111101001",
			1761 => "0001101111000100000100",
			1762 => "0000000001101111101001",
			1763 => "0000000001101111101001",
			1764 => "0011101001010100000100",
			1765 => "0000000001101111101001",
			1766 => "0000000001101111101001",
			1767 => "0001110101111000001000",
			1768 => "0010100110000000000100",
			1769 => "0000000001101111101001",
			1770 => "0000000001101111101001",
			1771 => "0001100010111000001000",
			1772 => "0001000110001100000100",
			1773 => "0000000001101111101001",
			1774 => "0000000001101111101001",
			1775 => "0011011011101100001100",
			1776 => "0001001001010100001000",
			1777 => "0000000100011000000100",
			1778 => "0000000001101111101001",
			1779 => "0000000001101111101001",
			1780 => "0000000001101111101001",
			1781 => "0000101101100100000100",
			1782 => "0000000001101111101001",
			1783 => "0010010011001000000100",
			1784 => "0000000001101111101001",
			1785 => "0000000001101111101001",
			1786 => "0001111000000000111100",
			1787 => "0000000001101100100100",
			1788 => "0010111010100100010000",
			1789 => "0000000000111000001000",
			1790 => "0010110110001100000100",
			1791 => "1111111001110010011101",
			1792 => "0000001001110010011101",
			1793 => "0010000101011100000100",
			1794 => "0000000001110010011101",
			1795 => "1111111001110010011101",
			1796 => "0000001000111000000100",
			1797 => "1111111001110010011101",
			1798 => "0010001001000100001000",
			1799 => "0001011111011000000100",
			1800 => "0000001001110010011101",
			1801 => "0000001001110010011101",
			1802 => "0001011101101000000100",
			1803 => "0000001001110010011101",
			1804 => "0000000001110010011101",
			1805 => "0000010000011000001100",
			1806 => "0000111001010100001000",
			1807 => "0000101101010000000100",
			1808 => "0000001001110010011101",
			1809 => "1111111001110010011101",
			1810 => "1111111001110010011101",
			1811 => "0010100011000100001000",
			1812 => "0011110000100000000100",
			1813 => "1111111001110010011101",
			1814 => "0000000001110010011101",
			1815 => "0000000001110010011101",
			1816 => "0000001100111000011100",
			1817 => "0011101100101100001100",
			1818 => "0001111000111000001000",
			1819 => "0000010111100100000100",
			1820 => "1111111001110010011101",
			1821 => "0000000001110010011101",
			1822 => "1111111001110010011101",
			1823 => "0000110001001000001100",
			1824 => "0001111100110000001000",
			1825 => "0000011000011000000100",
			1826 => "0000000001110010011101",
			1827 => "1111111001110010011101",
			1828 => "0000001001110010011101",
			1829 => "1111111001110010011101",
			1830 => "1111111001110010011101",
			1831 => "0011001010100100010000",
			1832 => "0001100101111000000100",
			1833 => "0000000001110100110001",
			1834 => "0010000011010000001000",
			1835 => "0010001010100100000100",
			1836 => "0000000001110100110001",
			1837 => "0000000001110100110001",
			1838 => "0000000001110100110001",
			1839 => "0011101000100000010100",
			1840 => "0000001000111000000100",
			1841 => "0000000001110100110001",
			1842 => "0000000000110100001100",
			1843 => "0000110110001100001000",
			1844 => "0010110011010000000100",
			1845 => "0000000001110100110001",
			1846 => "0000000001110100110001",
			1847 => "0000000001110100110001",
			1848 => "0000000001110100110001",
			1849 => "0011111010100000001000",
			1850 => "0001010001010000000100",
			1851 => "0000000001110100110001",
			1852 => "0000000001110100110001",
			1853 => "0011011011101100001100",
			1854 => "0011110010000000001000",
			1855 => "0001001111101000000100",
			1856 => "0000000001110100110001",
			1857 => "0000000001110100110001",
			1858 => "0000000001110100110001",
			1859 => "0011001001001000001000",
			1860 => "0000011000111100000100",
			1861 => "0000000001110100110001",
			1862 => "0000000001110100110001",
			1863 => "0010101001011000001000",
			1864 => "0000000100011000000100",
			1865 => "0000000001110100110001",
			1866 => "0000000001110100110001",
			1867 => "0000000001110100110001",
			1868 => "0000010111100100110000",
			1869 => "0011101111100000100000",
			1870 => "0010110110001100000100",
			1871 => "0000000001110111101101",
			1872 => "0010001001000100010100",
			1873 => "0001010011000000001100",
			1874 => "0000101101101100001000",
			1875 => "0000000011000000000100",
			1876 => "0000000001110111101101",
			1877 => "0000000001110111101101",
			1878 => "0000000001110111101101",
			1879 => "0000100100011100000100",
			1880 => "0000000001110111101101",
			1881 => "0000000001110111101101",
			1882 => "0000001110010100000100",
			1883 => "0000000001110111101101",
			1884 => "0000000001110111101101",
			1885 => "0000100100011100000100",
			1886 => "0000000001110111101101",
			1887 => "0001010001011000001000",
			1888 => "0001101110111100000100",
			1889 => "0000000001110111101101",
			1890 => "0000000001110111101101",
			1891 => "0000000001110111101101",
			1892 => "0011101001000000100000",
			1893 => "0000011101000000010100",
			1894 => "0010110011010000001000",
			1895 => "0000000001101000000100",
			1896 => "0000000001110111101101",
			1897 => "0000000001110111101101",
			1898 => "0001111000000000001000",
			1899 => "0000000001101100000100",
			1900 => "0000000001110111101101",
			1901 => "0000000001110111101101",
			1902 => "0000000001110111101101",
			1903 => "0001000111011100001000",
			1904 => "0000001000100000000100",
			1905 => "0000000001110111101101",
			1906 => "0000000001110111101101",
			1907 => "0000000001110111101101",
			1908 => "0010010001010000001000",
			1909 => "0010001001001100000100",
			1910 => "0000000001110111101101",
			1911 => "1111111001110111101101",
			1912 => "0010100000111100000100",
			1913 => "0000000001110111101101",
			1914 => "0000000001110111101101",
			1915 => "0000100000001100100100",
			1916 => "0001010111110000000100",
			1917 => "0000001001111000111001",
			1918 => "0011001011101100000100",
			1919 => "1111111001111000111001",
			1920 => "0000001000000100000100",
			1921 => "1111111001111000111001",
			1922 => "0000101111100000001000",
			1923 => "0000011101000000000100",
			1924 => "0000001001111000111001",
			1925 => "0000000001111000111001",
			1926 => "0000010111100100001000",
			1927 => "0011001001001000000100",
			1928 => "0000000001111000111001",
			1929 => "0000001001111000111001",
			1930 => "0011000101010100000100",
			1931 => "1111111001111000111001",
			1932 => "0000000001111000111001",
			1933 => "1111111001111000111001",
			1934 => "0001111000000100101100",
			1935 => "0000101101000100011000",
			1936 => "0010110110001100000100",
			1937 => "1111111001111011010101",
			1938 => "0011100011000100010000",
			1939 => "0000011101000000001100",
			1940 => "0010100110010000000100",
			1941 => "0000010001111011010101",
			1942 => "0010111010100100000100",
			1943 => "0000001001111011010101",
			1944 => "0000010001111011010101",
			1945 => "0000001001111011010101",
			1946 => "0000000001111011010101",
			1947 => "0010001111111100010000",
			1948 => "0000100101001100001100",
			1949 => "0001101001101100000100",
			1950 => "0000000001111011010101",
			1951 => "0001011000000100000100",
			1952 => "0000010001111011010101",
			1953 => "0000000001111011010101",
			1954 => "1111111001111011010101",
			1955 => "1111111001111011010101",
			1956 => "0000100111101000011100",
			1957 => "0000001000101000000100",
			1958 => "1111111001111011010101",
			1959 => "0000101101100100001000",
			1960 => "0001000101011100000100",
			1961 => "0000010001111011010101",
			1962 => "0000001001111011010101",
			1963 => "0001000100101100001100",
			1964 => "0001001100101000000100",
			1965 => "1111111001111011010101",
			1966 => "0000011001100000000100",
			1967 => "0000010001111011010101",
			1968 => "0000000001111011010101",
			1969 => "1111111001111011010101",
			1970 => "0001010101101100000100",
			1971 => "0000000001111011010101",
			1972 => "1111111001111011010101",
			1973 => "0011001010100100010000",
			1974 => "0001100101111000000100",
			1975 => "0000000001111101110001",
			1976 => "0010000011010000001000",
			1977 => "0010001010100100000100",
			1978 => "0000000001111101110001",
			1979 => "0000000001111101110001",
			1980 => "0000000001111101110001",
			1981 => "0011101000100000010100",
			1982 => "0000001000111000000100",
			1983 => "0000000001111101110001",
			1984 => "0000000000110100001100",
			1985 => "0000110110001100001000",
			1986 => "0010110011010000000100",
			1987 => "0000000001111101110001",
			1988 => "0000000001111101110001",
			1989 => "0000000001111101110001",
			1990 => "0000000001111101110001",
			1991 => "0011111010100000001100",
			1992 => "0011000101011100000100",
			1993 => "0000000001111101110001",
			1994 => "0011000101101100000100",
			1995 => "0000000001111101110001",
			1996 => "0000000001111101110001",
			1997 => "0011011011101100001100",
			1998 => "0011110010000000001000",
			1999 => "0001001111101000000100",
			2000 => "0000000001111101110001",
			2001 => "0000000001111101110001",
			2002 => "0000000001111101110001",
			2003 => "0011001001001000001000",
			2004 => "0000011000111100000100",
			2005 => "0000000001111101110001",
			2006 => "0000000001111101110001",
			2007 => "0010101001011000001000",
			2008 => "0000000100011000000100",
			2009 => "0000000001111101110001",
			2010 => "0000000001111101110001",
			2011 => "0000000001111101110001",
			2012 => "0011101000100000011100",
			2013 => "0010111010100100001100",
			2014 => "0001100101111000000100",
			2015 => "0000000010000000110101",
			2016 => "0000000000111000000100",
			2017 => "0000000010000000110101",
			2018 => "0000000010000000110101",
			2019 => "0001111111011000001000",
			2020 => "0000000000110100000100",
			2021 => "0000000010000000110101",
			2022 => "0000000010000000110101",
			2023 => "0001101100010000000100",
			2024 => "0000000010000000110101",
			2025 => "0000000010000000110101",
			2026 => "0011001001001000110100",
			2027 => "0010001001001100010100",
			2028 => "0000111101101000001000",
			2029 => "0001100010110000000100",
			2030 => "0000000010000000110101",
			2031 => "0000000010000000110101",
			2032 => "0000010111100100001000",
			2033 => "0000011000111100000100",
			2034 => "0000000010000000110101",
			2035 => "0000000010000000110101",
			2036 => "0000000010000000110101",
			2037 => "0001011000000100010000",
			2038 => "0001011111011000001000",
			2039 => "0011010110110100000100",
			2040 => "0000000010000000110101",
			2041 => "0000000010000000110101",
			2042 => "0000001011011000000100",
			2043 => "0000000010000000110101",
			2044 => "0000000010000000110101",
			2045 => "0011001100101000000100",
			2046 => "1111111010000000110101",
			2047 => "0011010111011100001000",
			2048 => "0010001111111100000100",
			2049 => "0000000010000000110101",
			2050 => "0000000010000000110101",
			2051 => "0000000010000000110101",
			2052 => "0011010011010000001000",
			2053 => "0001001001011000000100",
			2054 => "0000000010000000110101",
			2055 => "0000000010000000110101",
			2056 => "0010010001010000000100",
			2057 => "0000000010000000110101",
			2058 => "0010100000111100000100",
			2059 => "0000000010000000110101",
			2060 => "0000000010000000110101",
			2061 => "0000100010110000100000",
			2062 => "0001010110101100011000",
			2063 => "0010110110001100000100",
			2064 => "0000000010000011010001",
			2065 => "0000101010000100000100",
			2066 => "0000000010000011010001",
			2067 => "0000000000110100001100",
			2068 => "0001111001010000001000",
			2069 => "0001000001110000000100",
			2070 => "0000000010000011010001",
			2071 => "0000000010000011010001",
			2072 => "0000000010000011010001",
			2073 => "0000000010000011010001",
			2074 => "0010010110000000000100",
			2075 => "0000000010000011010001",
			2076 => "0000000010000011010001",
			2077 => "0011001001001000100000",
			2078 => "0011011011101100011100",
			2079 => "0010010111011100000100",
			2080 => "0000000010000011010001",
			2081 => "0010000011010000001100",
			2082 => "0001000110000000000100",
			2083 => "0000000010000011010001",
			2084 => "0000111001010100000100",
			2085 => "0000000010000011010001",
			2086 => "0000000010000011010001",
			2087 => "0010101000111000001000",
			2088 => "0000100000001100000100",
			2089 => "0000000010000011010001",
			2090 => "0000000010000011010001",
			2091 => "0000000010000011010001",
			2092 => "0000000010000011010001",
			2093 => "0000010111100100001000",
			2094 => "0001010010111000000100",
			2095 => "0000000010000011010001",
			2096 => "0000000010000011010001",
			2097 => "0010010001001000000100",
			2098 => "0000000010000011010001",
			2099 => "0000000010000011010001",
			2100 => "0000100000001100110100",
			2101 => "0010001001000100011100",
			2102 => "0001010000111000011000",
			2103 => "0011000110110100000100",
			2104 => "1111111010000100111101",
			2105 => "0010100110010000000100",
			2106 => "0000001010000100111101",
			2107 => "0011001010100100001000",
			2108 => "0010001001001100000100",
			2109 => "0000000010000100111101",
			2110 => "1111111010000100111101",
			2111 => "0000001000111000000100",
			2112 => "1111111010000100111101",
			2113 => "0000000010000100111101",
			2114 => "1111111010000100111101",
			2115 => "0001000101101100010100",
			2116 => "0000100011000100001000",
			2117 => "0001011101000000000100",
			2118 => "0000000010000100111101",
			2119 => "1111111010000100111101",
			2120 => "0000000010110100001000",
			2121 => "0011001100101000000100",
			2122 => "0000000010000100111101",
			2123 => "0000001010000100111101",
			2124 => "1111111010000100111101",
			2125 => "1111111010000100111101",
			2126 => "1111111010000100111101",
			2127 => "0011001011101100000100",
			2128 => "0000000010000111000001",
			2129 => "0010001111111100100000",
			2130 => "0001011010011100011000",
			2131 => "0011110011010100010100",
			2132 => "0010101110011000001100",
			2133 => "0000001010100000001000",
			2134 => "0000001000000100000100",
			2135 => "0000000010000111000001",
			2136 => "0000000010000111000001",
			2137 => "0000000010000111000001",
			2138 => "0001010111011100000100",
			2139 => "0000000010000111000001",
			2140 => "0000000010000111000001",
			2141 => "0000000010000111000001",
			2142 => "0010110101011100000100",
			2143 => "0000000010000111000001",
			2144 => "0000000010000111000001",
			2145 => "0010110101011100010000",
			2146 => "0011100011000100001100",
			2147 => "0001111001000100000100",
			2148 => "0000000010000111000001",
			2149 => "0000001001000000000100",
			2150 => "0000000010000111000001",
			2151 => "0000000010000111000001",
			2152 => "0000000010000111000001",
			2153 => "0000101110010000001100",
			2154 => "0001101000111000001000",
			2155 => "0001111111011000000100",
			2156 => "0000000010000111000001",
			2157 => "0000000010000111000001",
			2158 => "0000000010000111000001",
			2159 => "0000000010000111000001",
			2160 => "0000100000001100110100",
			2161 => "0000001000000100000100",
			2162 => "1111111010001000101101",
			2163 => "0001001110011000010100",
			2164 => "0010111011101100001000",
			2165 => "0011011111011100000100",
			2166 => "0000000010001000101101",
			2167 => "1111111010001000101101",
			2168 => "0000001010011000000100",
			2169 => "0000001010001000101101",
			2170 => "0001101001101100000100",
			2171 => "1111111010001000101101",
			2172 => "0000001010001000101101",
			2173 => "0010001001000100010000",
			2174 => "0011001001001000001100",
			2175 => "0001011010011100001000",
			2176 => "0011000011010000000100",
			2177 => "0000000010001000101101",
			2178 => "0000000010001000101101",
			2179 => "1111111010001000101101",
			2180 => "0000001010001000101101",
			2181 => "0001000101101100001000",
			2182 => "0010101000000000000100",
			2183 => "0000000010001000101101",
			2184 => "0000001010001000101101",
			2185 => "1111111010001000101101",
			2186 => "1111111010001000101101",
			2187 => "0011110110100001000000",
			2188 => "0010110101011100101000",
			2189 => "0010001111111100011000",
			2190 => "0001011010011100010100",
			2191 => "0011000110110100000100",
			2192 => "0000000010001010110001",
			2193 => "0011110111010100001000",
			2194 => "0011110100101100000100",
			2195 => "0000000010001010110001",
			2196 => "0000000010001010110001",
			2197 => "0000000100001000000100",
			2198 => "0000000010001010110001",
			2199 => "0000000010001010110001",
			2200 => "0000000010001010110001",
			2201 => "0011110001011000001100",
			2202 => "0010101010000100001000",
			2203 => "0010101000011000000100",
			2204 => "0000000010001010110001",
			2205 => "0000000010001010110001",
			2206 => "0000000010001010110001",
			2207 => "0000000010001010110001",
			2208 => "0001101000111000001000",
			2209 => "0001111111011000000100",
			2210 => "0000000010001010110001",
			2211 => "0000000010001010110001",
			2212 => "0000111000100000001100",
			2213 => "0000001100111000001000",
			2214 => "0010100011000000000100",
			2215 => "0000000010001010110001",
			2216 => "0000000010001010110001",
			2217 => "0000000010001010110001",
			2218 => "0000000010001010110001",
			2219 => "0000000010001010110001",
			2220 => "0000100101001101001000",
			2221 => "0011001001001000110000",
			2222 => "0010001001001100001100",
			2223 => "0001101100110100001000",
			2224 => "0000100000111000000100",
			2225 => "0000000010001101000101",
			2226 => "0000000010001101000101",
			2227 => "0000000010001101000101",
			2228 => "0011100011000100010000",
			2229 => "0010111010100100001000",
			2230 => "0001101111011000000100",
			2231 => "0000000010001101000101",
			2232 => "0000000010001101000101",
			2233 => "0000001000111000000100",
			2234 => "0000000010001101000101",
			2235 => "0000000010001101000101",
			2236 => "0000100010110100001100",
			2237 => "0001001110011000000100",
			2238 => "0000000010001101000101",
			2239 => "0010101111101000000100",
			2240 => "1111111010001101000101",
			2241 => "0000000010001101000101",
			2242 => "0010001111111100000100",
			2243 => "0000000010001101000101",
			2244 => "0000000010001101000101",
			2245 => "0001101000111000001000",
			2246 => "0001111111011000000100",
			2247 => "0000000010001101000101",
			2248 => "0000000010001101000101",
			2249 => "0010101100010000001000",
			2250 => "0000001101100100000100",
			2251 => "0000000010001101000101",
			2252 => "0000000010001101000101",
			2253 => "0000000010000000000100",
			2254 => "0000000010001101000101",
			2255 => "0000001010001101000101",
			2256 => "1111111010001101000101",
			2257 => "0001010110101100110100",
			2258 => "0010110110001100001000",
			2259 => "0010010111011100000100",
			2260 => "0000000010010000000001",
			2261 => "0000000010010000000001",
			2262 => "0001101111000100101000",
			2263 => "0010101111111100010100",
			2264 => "0000001010100000001100",
			2265 => "0001110011001000000100",
			2266 => "0000000010010000000001",
			2267 => "0001100101111000000100",
			2268 => "0000000010010000000001",
			2269 => "0000000010010000000001",
			2270 => "0000010011110000000100",
			2271 => "0000000010010000000001",
			2272 => "0000000010010000000001",
			2273 => "0000001011000000000100",
			2274 => "0000000010010000000001",
			2275 => "0000000000110100001000",
			2276 => "0001110101101100000100",
			2277 => "0000000010010000000001",
			2278 => "0000000010010000000001",
			2279 => "0010011001000100000100",
			2280 => "0000000010010000000001",
			2281 => "0000000010010000000001",
			2282 => "0000000010010000000001",
			2283 => "0011001001001000011100",
			2284 => "0010000011010000001000",
			2285 => "0000111001010100000100",
			2286 => "0000000010010000000001",
			2287 => "0000000010010000000001",
			2288 => "0011111100001100000100",
			2289 => "0000000010010000000001",
			2290 => "0010110101011100001000",
			2291 => "0011010110110100000100",
			2292 => "0000000010010000000001",
			2293 => "0000000010010000000001",
			2294 => "0011011010100100000100",
			2295 => "0000000010010000000001",
			2296 => "0000000010010000000001",
			2297 => "0010001001000100001000",
			2298 => "0001001001011000000100",
			2299 => "0000000010010000000001",
			2300 => "0000000010010000000001",
			2301 => "0001001101101000000100",
			2302 => "0000000010010000000001",
			2303 => "0000000010010000000001",
			2304 => "0000100000001101000000",
			2305 => "0011000011010000010100",
			2306 => "0000000000111000001000",
			2307 => "0010110110001100000100",
			2308 => "0000000010010010000101",
			2309 => "0000000010010010000101",
			2310 => "0010000011010000000100",
			2311 => "0000000010010010000101",
			2312 => "0000000100110000000100",
			2313 => "0000000010010010000101",
			2314 => "0000000010010010000101",
			2315 => "0001010000111000101000",
			2316 => "0010101111111100010000",
			2317 => "0000001101000100001000",
			2318 => "0000001000111000000100",
			2319 => "0000000010010010000101",
			2320 => "0000000010010010000101",
			2321 => "0000010011110000000100",
			2322 => "0000000010010010000101",
			2323 => "0000000010010010000101",
			2324 => "0000011000011000001100",
			2325 => "0010001001000100001000",
			2326 => "0001010011000000000100",
			2327 => "0000000010010010000101",
			2328 => "0000000010010010000101",
			2329 => "0000000010010010000101",
			2330 => "0001011111101000001000",
			2331 => "0000001110100100000100",
			2332 => "0000000010010010000101",
			2333 => "0000000010010010000101",
			2334 => "0000000010010010000101",
			2335 => "0000000010010010000101",
			2336 => "0000000010010010000101",
			2337 => "0000100101001100110000",
			2338 => "0000101010000100000100",
			2339 => "1111111010010011101001",
			2340 => "0011111011111000010100",
			2341 => "0001010011000000010000",
			2342 => "0010110110001100000100",
			2343 => "1111111010010011101001",
			2344 => "0001111001010000001000",
			2345 => "0000101001101100000100",
			2346 => "0000001010010011101001",
			2347 => "0000000010010011101001",
			2348 => "1111111010010011101001",
			2349 => "0000000010010011101001",
			2350 => "0001010000111000010100",
			2351 => "0001111001000100000100",
			2352 => "1111111010010011101001",
			2353 => "0011001100101000001000",
			2354 => "0010000011010000000100",
			2355 => "0000001010010011101001",
			2356 => "0000000010010011101001",
			2357 => "0011000101101100000100",
			2358 => "0000001010010011101001",
			2359 => "0000000010010011101001",
			2360 => "1111111010010011101001",
			2361 => "1111111010010011101001",
			2362 => "0011101111100001000000",
			2363 => "0010001001000100101000",
			2364 => "0010110110001100000100",
			2365 => "0000000010010110110101",
			2366 => "0000100111100000011100",
			2367 => "0000111110011000010000",
			2368 => "0001111001001000001000",
			2369 => "0000101111101000000100",
			2370 => "0000000010010110110101",
			2371 => "0000000010010110110101",
			2372 => "0010100110010000000100",
			2373 => "0000000010010110110101",
			2374 => "0000000010010110110101",
			2375 => "0000011000011000001000",
			2376 => "0001001111101000000100",
			2377 => "0000001010010110110101",
			2378 => "0000000010010110110101",
			2379 => "0000000010010110110101",
			2380 => "0011100001010100000100",
			2381 => "0000000010010110110101",
			2382 => "0000000010010110110101",
			2383 => "0001000101101100010100",
			2384 => "0010100011000000010000",
			2385 => "0001010011010000001100",
			2386 => "0000000110100000001000",
			2387 => "0000001011000000000100",
			2388 => "0000000010010110110101",
			2389 => "0000000010010110110101",
			2390 => "0000000010010110110101",
			2391 => "0000000010010110110101",
			2392 => "0000000010010110110101",
			2393 => "0000000010010110110101",
			2394 => "0010101000111000010000",
			2395 => "0011000011010000001000",
			2396 => "0011011111011100000100",
			2397 => "0000000010010110110101",
			2398 => "0000000010010110110101",
			2399 => "0011110100001100000100",
			2400 => "0000000010010110110101",
			2401 => "0000000010010110110101",
			2402 => "0010010001001000010100",
			2403 => "0010000011010000001000",
			2404 => "0011010110110100000100",
			2405 => "0000000010010110110101",
			2406 => "0000000010010110110101",
			2407 => "0011001001001000000100",
			2408 => "1111111010010110110101",
			2409 => "0011000101101100000100",
			2410 => "0000000010010110110101",
			2411 => "0000000010010110110101",
			2412 => "0000000010010110110101",
			2413 => "0011100010011101010000",
			2414 => "0010110101011100110000",
			2415 => "0010011101101000101000",
			2416 => "0011000101010100011000",
			2417 => "0001010110101100010000",
			2418 => "0011001011101100001000",
			2419 => "0001101111011000000100",
			2420 => "0000000010011001100001",
			2421 => "0000000010011001100001",
			2422 => "0011110001010100000100",
			2423 => "0000000010011001100001",
			2424 => "0000000010011001100001",
			2425 => "0000010001110000000100",
			2426 => "0000000010011001100001",
			2427 => "0000000010011001100001",
			2428 => "0000000001111000001100",
			2429 => "0000111100101000001000",
			2430 => "0001011101000000000100",
			2431 => "0000000010011001100001",
			2432 => "0000000010011001100001",
			2433 => "0000000010011001100001",
			2434 => "0000000010011001100001",
			2435 => "0011001001001000000100",
			2436 => "0000000010011001100001",
			2437 => "0000000010011001100001",
			2438 => "0000010111100100001100",
			2439 => "0010100101011100001000",
			2440 => "0001011101000000000100",
			2441 => "0000000010011001100001",
			2442 => "0000000010011001100001",
			2443 => "0000000010011001100001",
			2444 => "0000000011101100001100",
			2445 => "0001101000111000001000",
			2446 => "0001111111011000000100",
			2447 => "0000000010011001100001",
			2448 => "0000000010011001100001",
			2449 => "0000000010011001100001",
			2450 => "0001111001010100000100",
			2451 => "0000000010011001100001",
			2452 => "0000000010011001100001",
			2453 => "0010001011000000000100",
			2454 => "1111111010011001100001",
			2455 => "0000000010011001100001",
			2456 => "0011101010110101000100",
			2457 => "0011001011101100001000",
			2458 => "0001100011001000000100",
			2459 => "0000000010011011110101",
			2460 => "0000000010011011110101",
			2461 => "0001010110101100100000",
			2462 => "0000001000111000001000",
			2463 => "0000111001100000000100",
			2464 => "0000000010011011110101",
			2465 => "0000000010011011110101",
			2466 => "0000001000110100001100",
			2467 => "0010101010100100001000",
			2468 => "0010100110010000000100",
			2469 => "0000000010011011110101",
			2470 => "0000000010011011110101",
			2471 => "0000000010011011110101",
			2472 => "0001111100010000001000",
			2473 => "0001111000000100000100",
			2474 => "0000000010011011110101",
			2475 => "0000000010011011110101",
			2476 => "0000000010011011110101",
			2477 => "0011001001001000010000",
			2478 => "0011111100001100000100",
			2479 => "0000000010011011110101",
			2480 => "0001100000100000000100",
			2481 => "0000000010011011110101",
			2482 => "0011011011101100000100",
			2483 => "0000000010011011110101",
			2484 => "0000000010011011110101",
			2485 => "0011010111011100000100",
			2486 => "0000000010011011110101",
			2487 => "0001110001010000000100",
			2488 => "0000000010011011110101",
			2489 => "0000000010011011110101",
			2490 => "0001111000000000000100",
			2491 => "0000000010011011110101",
			2492 => "0000000010011011110101",
			2493 => "0000100000001100110100",
			2494 => "0000101010000100000100",
			2495 => "1111111010011101100001",
			2496 => "0000001001111100010100",
			2497 => "0010111010000100010000",
			2498 => "0010110110001100000100",
			2499 => "1111111010011101100001",
			2500 => "0000010011110000001000",
			2501 => "0000101001010100000100",
			2502 => "0000001010011101100001",
			2503 => "0000001010011101100001",
			2504 => "0000001010011101100001",
			2505 => "0000000010011101100001",
			2506 => "0001010000111000011000",
			2507 => "0001011001001000001000",
			2508 => "0001100001111100000100",
			2509 => "1111111010011101100001",
			2510 => "0000000010011101100001",
			2511 => "0010001001000100001000",
			2512 => "0011000011010000000100",
			2513 => "0000000010011101100001",
			2514 => "0000001010011101100001",
			2515 => "0001000110000000000100",
			2516 => "0000000010011101100001",
			2517 => "1111111010011101100001",
			2518 => "1111111010011101100001",
			2519 => "1111111010011101100001",
			2520 => "0011101010110101000000",
			2521 => "0011001011101100001000",
			2522 => "0011111000000100000100",
			2523 => "0000000010011111101101",
			2524 => "0000000010011111101101",
			2525 => "0001011010011100110000",
			2526 => "0011110100000000011100",
			2527 => "0000100010110000010000",
			2528 => "0010111010100100001000",
			2529 => "0000100001111100000100",
			2530 => "0000000010011111101101",
			2531 => "0000000010011111101101",
			2532 => "0000001000111000000100",
			2533 => "0000000010011111101101",
			2534 => "0000000010011111101101",
			2535 => "0011011010100100000100",
			2536 => "0000000010011111101101",
			2537 => "0011010111011100000100",
			2538 => "0000000010011111101101",
			2539 => "0000000010011111101101",
			2540 => "0010001111111100001000",
			2541 => "0000000100001000000100",
			2542 => "0000000010011111101101",
			2543 => "0000000010011111101101",
			2544 => "0010001111011000001000",
			2545 => "0000000100110000000100",
			2546 => "0000000010011111101101",
			2547 => "0000000010011111101101",
			2548 => "0000000010011111101101",
			2549 => "0011001001001000000100",
			2550 => "0000000010011111101101",
			2551 => "0000000010011111101101",
			2552 => "0010101010000100000100",
			2553 => "0000000010011111101101",
			2554 => "0000000010011111101101",
			2555 => "0000100000001101000000",
			2556 => "0011001011101100001000",
			2557 => "0010100110001100000100",
			2558 => "0000000010100001110001",
			2559 => "1111111010100001110001",
			2560 => "0001001110011000011100",
			2561 => "0000001000000100000100",
			2562 => "1111111010100001110001",
			2563 => "0000111100101000001100",
			2564 => "0000001010100000000100",
			2565 => "0000001010100001110001",
			2566 => "0001101110010100000100",
			2567 => "1111111010100001110001",
			2568 => "0000000010100001110001",
			2569 => "0010101010000100000100",
			2570 => "0000001010100001110001",
			2571 => "0010101111011000000100",
			2572 => "0000000010100001110001",
			2573 => "0000001010100001110001",
			2574 => "0010001001000100010000",
			2575 => "0011001001001000001100",
			2576 => "0001011010011100001000",
			2577 => "0011000101010100000100",
			2578 => "0000000010100001110001",
			2579 => "0000000010100001110001",
			2580 => "1111111010100001110001",
			2581 => "0000001010100001110001",
			2582 => "0001000101101100001000",
			2583 => "0010101000000000000100",
			2584 => "1111111010100001110001",
			2585 => "0000001010100001110001",
			2586 => "1111111010100001110001",
			2587 => "1111111010100001110001",
			2588 => "0001010110101101000000",
			2589 => "0010110110001100001000",
			2590 => "0010010111011100000100",
			2591 => "0000000010100101000101",
			2592 => "0000000010100101000101",
			2593 => "0001101111000100110100",
			2594 => "0010101111111100011100",
			2595 => "0001011111011100001100",
			2596 => "0000000011000000000100",
			2597 => "0000000010100101000101",
			2598 => "0000001010001100000100",
			2599 => "0000000010100101000101",
			2600 => "0000000010100101000101",
			2601 => "0000111100101000001000",
			2602 => "0010000011001000000100",
			2603 => "0000000010100101000101",
			2604 => "0000000010100101000101",
			2605 => "0010000011100100000100",
			2606 => "0000000010100101000101",
			2607 => "0000000010100101000101",
			2608 => "0010010110000000001000",
			2609 => "0001110101101100000100",
			2610 => "0000000010100101000101",
			2611 => "0000000010100101000101",
			2612 => "0000000000110100001000",
			2613 => "0000001001000000000100",
			2614 => "0000000010100101000101",
			2615 => "0000000010100101000101",
			2616 => "0001111100110000000100",
			2617 => "0000000010100101000101",
			2618 => "0000000010100101000101",
			2619 => "0000000010100101000101",
			2620 => "0011001001001000011100",
			2621 => "0010000011010000001000",
			2622 => "0000001011001000000100",
			2623 => "0000000010100101000101",
			2624 => "0000000010100101000101",
			2625 => "0010110101011100001100",
			2626 => "0001100011110100000100",
			2627 => "0000000010100101000101",
			2628 => "0011010110110100000100",
			2629 => "0000000010100101000101",
			2630 => "0000000010100101000101",
			2631 => "0011111001110000000100",
			2632 => "0000000010100101000101",
			2633 => "0000000010100101000101",
			2634 => "0010001001000100001000",
			2635 => "0001001001011000000100",
			2636 => "0000000010100101000101",
			2637 => "0000000010100101000101",
			2638 => "0001001101101000000100",
			2639 => "0000000010100101000101",
			2640 => "0000000010100101000101",
			2641 => "0011100000100001010000",
			2642 => "0001001110011000100100",
			2643 => "0000111100101000100000",
			2644 => "0001001001100000010000",
			2645 => "0000000011000000000100",
			2646 => "1111111010100111101001",
			2647 => "0000001010100000000100",
			2648 => "0000001010100111101001",
			2649 => "0010100110110100000100",
			2650 => "1111111010100111101001",
			2651 => "0000000010100111101001",
			2652 => "0001111010000100001000",
			2653 => "0010101110011000000100",
			2654 => "0000000010100111101001",
			2655 => "0000000010100111101001",
			2656 => "0010000011001000000100",
			2657 => "1111111010100111101001",
			2658 => "0000000010100111101001",
			2659 => "0000001010100111101001",
			2660 => "0010001001000100011100",
			2661 => "0011001100101000010000",
			2662 => "0001011010011100001100",
			2663 => "0011001110011000000100",
			2664 => "1111111010100111101001",
			2665 => "0011101000100000000100",
			2666 => "0000001010100111101001",
			2667 => "0000000010100111101001",
			2668 => "1111111010100111101001",
			2669 => "0001000011000100001000",
			2670 => "0001011101001000000100",
			2671 => "0000000010100111101001",
			2672 => "0000001010100111101001",
			2673 => "1111111010100111101001",
			2674 => "0001000101101100001100",
			2675 => "0010101000000000001000",
			2676 => "0000011001100000000100",
			2677 => "0000000010100111101001",
			2678 => "1111111010100111101001",
			2679 => "0000001010100111101001",
			2680 => "1111111010100111101001",
			2681 => "1111111010100111101001",
			2682 => "0000001100111000111100",
			2683 => "0000101010000100000100",
			2684 => "1111111010101001101101",
			2685 => "0000001001111100011000",
			2686 => "0010110110001100000100",
			2687 => "1111111010101001101101",
			2688 => "0000011101000000001100",
			2689 => "0000011001100100000100",
			2690 => "0000001010101001101101",
			2691 => "0000010011110000000100",
			2692 => "0000001010101001101101",
			2693 => "0000001010101001101101",
			2694 => "0001000101010100000100",
			2695 => "0000001010101001101101",
			2696 => "1111111010101001101101",
			2697 => "0001010000111000011100",
			2698 => "0010001001000100010000",
			2699 => "0001010101010100001000",
			2700 => "0001001001100000000100",
			2701 => "0000000010101001101101",
			2702 => "1111111010101001101101",
			2703 => "0011000101010100000100",
			2704 => "0000000010101001101101",
			2705 => "0000001010101001101101",
			2706 => "0001001001000100001000",
			2707 => "0010000000110000000100",
			2708 => "1111111010101001101101",
			2709 => "0000001010101001101101",
			2710 => "1111111010101001101101",
			2711 => "1111111010101001101101",
			2712 => "0001010101101100000100",
			2713 => "0000000010101001101101",
			2714 => "1111111010101001101101",
			2715 => "0000100101001100111100",
			2716 => "0000101010000100000100",
			2717 => "1111111010101011101001",
			2718 => "0000101101000100011000",
			2719 => "0001011001010100010100",
			2720 => "0010110110001100000100",
			2721 => "1111111010101011101001",
			2722 => "0010111010100100001000",
			2723 => "0010001111111100000100",
			2724 => "0000001010101011101001",
			2725 => "1111111010101011101001",
			2726 => "0000001000111000000100",
			2727 => "1111111010101011101001",
			2728 => "0000001010101011101001",
			2729 => "0000000010101011101001",
			2730 => "0010110101011100010000",
			2731 => "0010001111111100001100",
			2732 => "0001101001101100000100",
			2733 => "1111111010101011101001",
			2734 => "0001001100010000000100",
			2735 => "0000001010101011101001",
			2736 => "1111111010101011101001",
			2737 => "1111111010101011101001",
			2738 => "0010101000000000001000",
			2739 => "0000110011010000000100",
			2740 => "0000000010101011101001",
			2741 => "1111111010101011101001",
			2742 => "0000110001001000000100",
			2743 => "0000001010101011101001",
			2744 => "1111111010101011101001",
			2745 => "1111111010101011101001",
			2746 => "0011100000100001001100",
			2747 => "0000010111100100101000",
			2748 => "0001001011111000100000",
			2749 => "0010110110001100000100",
			2750 => "0000000010101110000101",
			2751 => "0010001001000100010000",
			2752 => "0010110101011100001000",
			2753 => "0000111101001000000100",
			2754 => "0000000010101110000101",
			2755 => "1111111010101110000101",
			2756 => "0000001000101000000100",
			2757 => "0000000010101110000101",
			2758 => "0000001010101110000101",
			2759 => "0000000001011100001000",
			2760 => "0000001001001000000100",
			2761 => "0000000010101110000101",
			2762 => "0000000010101110000101",
			2763 => "1111111010101110000101",
			2764 => "0001110011001000000100",
			2765 => "0000000010101110000101",
			2766 => "1111111010101110000101",
			2767 => "0011000101010100001000",
			2768 => "0001000110001100000100",
			2769 => "0000000010101110000101",
			2770 => "1111111010101110000101",
			2771 => "0001111111011000001000",
			2772 => "0000101101000100000100",
			2773 => "0000001010101110000101",
			2774 => "0000000010101110000101",
			2775 => "0001101100110000000100",
			2776 => "1111111010101110000101",
			2777 => "0000000010110100001000",
			2778 => "0010101000101000000100",
			2779 => "0000001010101110000101",
			2780 => "0000000010101110000101",
			2781 => "0011111101000100000100",
			2782 => "1111111010101110000101",
			2783 => "0000000010101110000101",
			2784 => "1111111010101110000101",
			2785 => "0000100000001101000100",
			2786 => "0000101010000100000100",
			2787 => "1111111010110000010001",
			2788 => "0001010110101100100100",
			2789 => "0000000000110100010100",
			2790 => "0010110110001100000100",
			2791 => "1111111010110000010001",
			2792 => "0001000110110100001000",
			2793 => "0001101101101000000100",
			2794 => "0000001010110000010001",
			2795 => "0000001010110000010001",
			2796 => "0010111010100100000100",
			2797 => "0000000010110000010001",
			2798 => "0000001010110000010001",
			2799 => "0011110111010100000100",
			2800 => "1111111010110000010001",
			2801 => "0001101111000100001000",
			2802 => "0010001111111100000100",
			2803 => "0000001010110000010001",
			2804 => "0000000010110000010001",
			2805 => "1111111010110000010001",
			2806 => "0010001001000100010000",
			2807 => "0011001100101000001000",
			2808 => "0001000110101100000100",
			2809 => "0000000010110000010001",
			2810 => "1111111010110000010001",
			2811 => "0001000011000100000100",
			2812 => "0000001010110000010001",
			2813 => "1111111010110000010001",
			2814 => "0001111101001000001000",
			2815 => "0001111000000100000100",
			2816 => "1111111010110000010001",
			2817 => "1111111010110000010001",
			2818 => "0000000010110000010001",
			2819 => "1111111010110000010001",
			2820 => "0011100000100001011000",
			2821 => "0001001110011000100100",
			2822 => "0011000110110100000100",
			2823 => "1111111010110011000111",
			2824 => "0000101010000100000100",
			2825 => "0000000010110011000111",
			2826 => "0000111100101000010000",
			2827 => "0000001010100000001000",
			2828 => "0001011011101100000100",
			2829 => "0000001010110011000111",
			2830 => "0000000010110011000111",
			2831 => "0011110001011100000100",
			2832 => "1111111010110011000111",
			2833 => "0000000010110011000111",
			2834 => "0000010111100100000100",
			2835 => "0000001010110011000111",
			2836 => "0000011001100000000100",
			2837 => "0000000010110011000111",
			2838 => "0000000010110011000111",
			2839 => "0011001100101000011000",
			2840 => "0011011011101100010000",
			2841 => "0001011111011000000100",
			2842 => "0000000010110011000111",
			2843 => "0000111001010100001000",
			2844 => "0011000011010000000100",
			2845 => "0000000010110011000111",
			2846 => "0000001010110011000111",
			2847 => "1111111010110011000111",
			2848 => "0000010000011000000100",
			2849 => "0000000010110011000111",
			2850 => "1111111010110011000111",
			2851 => "0000001100110100001000",
			2852 => "0011011100101000000100",
			2853 => "0000000010110011000111",
			2854 => "1111111010110011000111",
			2855 => "0000100111100000000100",
			2856 => "0000001010110011000111",
			2857 => "0001100000100000001000",
			2858 => "0010010011001000000100",
			2859 => "1111111010110011000111",
			2860 => "0000000010110011000111",
			2861 => "0001001000100000000100",
			2862 => "0000001010110011000111",
			2863 => "0000000010110011000111",
			2864 => "1111111010110011000111",
			2865 => "0000000001101100011100",
			2866 => "0011000111011100010000",
			2867 => "0011101101001000001000",
			2868 => "0010110110001100000100",
			2869 => "0000000010110101001001",
			2870 => "0000000010110101001001",
			2871 => "0011111010011100000100",
			2872 => "0000000010110101001001",
			2873 => "0000000010110101001001",
			2874 => "0001101000111000001000",
			2875 => "0001111111011000000100",
			2876 => "0000000010110101001001",
			2877 => "0000000010110101001001",
			2878 => "0000000010110101001001",
			2879 => "0000010000011000010100",
			2880 => "0011101010100000001000",
			2881 => "0001111111011000000100",
			2882 => "0000000010110101001001",
			2883 => "0000000010110101001001",
			2884 => "0000101000110100000100",
			2885 => "0000000010110101001001",
			2886 => "0000100000001100000100",
			2887 => "0000000010110101001001",
			2888 => "0000000010110101001001",
			2889 => "0010111000101000010000",
			2890 => "0011101100001100001000",
			2891 => "0001100011110100000100",
			2892 => "0000000010110101001001",
			2893 => "0000000010110101001001",
			2894 => "0010000011010000000100",
			2895 => "0000000010110101001001",
			2896 => "0000000010110101001001",
			2897 => "0000000010110101001001",
			2898 => "0001010110101100100100",
			2899 => "0000000000110100010000",
			2900 => "0010110110001100000100",
			2901 => "0000000010110111001101",
			2902 => "0000101010000100000100",
			2903 => "0000000010110111001101",
			2904 => "0001000001110000000100",
			2905 => "0000000010110111001101",
			2906 => "0000000010110111001101",
			2907 => "0011110101110000000100",
			2908 => "0000000010110111001101",
			2909 => "0010010111011100000100",
			2910 => "0000000010110111001101",
			2911 => "0011110011010100001000",
			2912 => "0010001111111100000100",
			2913 => "0000000010110111001101",
			2914 => "0000000010110111001101",
			2915 => "0000000010110111001101",
			2916 => "0011001001001000010000",
			2917 => "0011100001011000000100",
			2918 => "0000000010110111001101",
			2919 => "0010000011010000000100",
			2920 => "0000000010110111001101",
			2921 => "0000011000111100000100",
			2922 => "0000000010110111001101",
			2923 => "0000000010110111001101",
			2924 => "0010001001000100001000",
			2925 => "0001001001011000000100",
			2926 => "0000000010110111001101",
			2927 => "0000000010110111001101",
			2928 => "0001001010000100000100",
			2929 => "0000000010110111001101",
			2930 => "0000000010110111001101",
			2931 => "0000000001101100100000",
			2932 => "0011000111011100010000",
			2933 => "0000000000111000001000",
			2934 => "0010110110001100000100",
			2935 => "0000000010111001011001",
			2936 => "0000000010111001011001",
			2937 => "0011110000111000000100",
			2938 => "0000000010111001011001",
			2939 => "0000000010111001011001",
			2940 => "0001101000111000001000",
			2941 => "0001111111011000000100",
			2942 => "0000000010111001011001",
			2943 => "0000000010111001011001",
			2944 => "0001011110011000000100",
			2945 => "0000000010111001011001",
			2946 => "0000000010111001011001",
			2947 => "0010001111111100100000",
			2948 => "0001101001101100000100",
			2949 => "0000000010111001011001",
			2950 => "0011100010011100010000",
			2951 => "0001011001000000001000",
			2952 => "0001110101111000000100",
			2953 => "0000000010111001011001",
			2954 => "0000000010111001011001",
			2955 => "0000001010111100000100",
			2956 => "0000000010111001011001",
			2957 => "0000000010111001011001",
			2958 => "0011000011010000000100",
			2959 => "0000000010111001011001",
			2960 => "0010011001001000000100",
			2961 => "0000000010111001011001",
			2962 => "0000000010111001011001",
			2963 => "0010111000101000000100",
			2964 => "0000000010111001011001",
			2965 => "0000000010111001011001",
			2966 => "0001010110101100101000",
			2967 => "0000000000110100010000",
			2968 => "0010110110001100000100",
			2969 => "0000000010111011101101",
			2970 => "0000101010000100000100",
			2971 => "0000000010111011101101",
			2972 => "0010011100110000000100",
			2973 => "0000000010111011101101",
			2974 => "0000000010111011101101",
			2975 => "0001101001101100000100",
			2976 => "0000000010111011101101",
			2977 => "0010010111011100000100",
			2978 => "0000000010111011101101",
			2979 => "0011110011010100001100",
			2980 => "0010001111111100000100",
			2981 => "0000000010111011101101",
			2982 => "0010111100101000000100",
			2983 => "0000000010111011101101",
			2984 => "0000000010111011101101",
			2985 => "0000000010111011101101",
			2986 => "0011001001001000010100",
			2987 => "0010000011010000001000",
			2988 => "0000111001010100000100",
			2989 => "0000000010111011101101",
			2990 => "0000000010111011101101",
			2991 => "0011111100001100000100",
			2992 => "0000000010111011101101",
			2993 => "0010110101011100000100",
			2994 => "0000000010111011101101",
			2995 => "0000000010111011101101",
			2996 => "0011010011010000001000",
			2997 => "0001001000100000000100",
			2998 => "0000000010111011101101",
			2999 => "0000000010111011101101",
			3000 => "0001001101101000000100",
			3001 => "0000000010111011101101",
			3002 => "0000000010111011101101",
			3003 => "0000101110010000110000",
			3004 => "0011000101010100011100",
			3005 => "0011011111011100000100",
			3006 => "0000000010111101011001",
			3007 => "0011101101001000001000",
			3008 => "0010111011101100000100",
			3009 => "0000000010111101011001",
			3010 => "0000000010111101011001",
			3011 => "0001011111011000000100",
			3012 => "0000000010111101011001",
			3013 => "0001010110101100000100",
			3014 => "0000000010111101011001",
			3015 => "0011111111100100000100",
			3016 => "0000000010111101011001",
			3017 => "0000000010111101011001",
			3018 => "0001001111101000010000",
			3019 => "0000001000101000000100",
			3020 => "0000000010111101011001",
			3021 => "0010101010100100001000",
			3022 => "0010101101000000000100",
			3023 => "0000000010111101011001",
			3024 => "0000000010111101011001",
			3025 => "0000000010111101011001",
			3026 => "0000000010111101011001",
			3027 => "0010000011010000000100",
			3028 => "0000000010111101011001",
			3029 => "0000000010111101011001",
			3030 => "0001111000000100101100",
			3031 => "0011110100101100010000",
			3032 => "0011001110011000001000",
			3033 => "0011011101000000000100",
			3034 => "1101101010111111101101",
			3035 => "1101100010111111101101",
			3036 => "0011000011010000000100",
			3037 => "1110100010111111101101",
			3038 => "1110101010111111101101",
			3039 => "0000010111100100010100",
			3040 => "0011000101010100010000",
			3041 => "0010101100010000001100",
			3042 => "0011111111100100001000",
			3043 => "0010101111111100000100",
			3044 => "1101100010111111101101",
			3045 => "1101111010111111101101",
			3046 => "1110010010111111101101",
			3047 => "1101100010111111101101",
			3048 => "1110011010111111101101",
			3049 => "0000101101000100000100",
			3050 => "1101110010111111101101",
			3051 => "1101100010111111101101",
			3052 => "0000100111101000011000",
			3053 => "0000001000101000000100",
			3054 => "1101100010111111101101",
			3055 => "0000000001101100000100",
			3056 => "1110100010111111101101",
			3057 => "0011001001001000001000",
			3058 => "0010000101011100000100",
			3059 => "1101111010111111101101",
			3060 => "1101100010111111101101",
			3061 => "0010101001011000000100",
			3062 => "1110001010111111101101",
			3063 => "1101110010111111101101",
			3064 => "0001010101101100000100",
			3065 => "1101101010111111101101",
			3066 => "1101100010111111101101",
			3067 => "0000010111100100110100",
			3068 => "0011001010100100010000",
			3069 => "0011011111011100001000",
			3070 => "0010111101000000000100",
			3071 => "0000000011000010001001",
			3072 => "0000000011000010001001",
			3073 => "0010000011010000000100",
			3074 => "0000000011000010001001",
			3075 => "0000000011000010001001",
			3076 => "0001001011111000011000",
			3077 => "0011110011010100010100",
			3078 => "0010101001001100001100",
			3079 => "0000001101000100001000",
			3080 => "0000001000000100000100",
			3081 => "0000000011000010001001",
			3082 => "0000000011000010001001",
			3083 => "0000000011000010001001",
			3084 => "0010001001000100000100",
			3085 => "0000000011000010001001",
			3086 => "0000000011000010001001",
			3087 => "0000000011000010001001",
			3088 => "0011001001001000000100",
			3089 => "0000000011000010001001",
			3090 => "0011000101101100000100",
			3091 => "0000000011000010001001",
			3092 => "0000000011000010001001",
			3093 => "0010010001010000010100",
			3094 => "0010001001001100000100",
			3095 => "0000000011000010001001",
			3096 => "0001010001100100000100",
			3097 => "0000000011000010001001",
			3098 => "0001011100011100000100",
			3099 => "0000000011000010001001",
			3100 => "0001010011110100000100",
			3101 => "0000000011000010001001",
			3102 => "0000000011000010001001",
			3103 => "0001001001001000000100",
			3104 => "0000000011000010001001",
			3105 => "0000000011000010001001",
			3106 => "0001011110011000001000",
			3107 => "0011111001001000000100",
			3108 => "0000000011000011110101",
			3109 => "0000000011000011110101",
			3110 => "0011000011010000001000",
			3111 => "0000000001101000000100",
			3112 => "0000000011000011110101",
			3113 => "0000000011000011110101",
			3114 => "0001110101111000001000",
			3115 => "0010100110000000000100",
			3116 => "0000000011000011110101",
			3117 => "0000000011000011110101",
			3118 => "0001100010111000001000",
			3119 => "0001000110001100000100",
			3120 => "0000000011000011110101",
			3121 => "0000000011000011110101",
			3122 => "0011011011101100001100",
			3123 => "0001001001010100001000",
			3124 => "0000000100011000000100",
			3125 => "0000000011000011110101",
			3126 => "0000000011000011110101",
			3127 => "0000000011000011110101",
			3128 => "0000101101100100000100",
			3129 => "0000000011000011110101",
			3130 => "0010010011001000000100",
			3131 => "0000000011000011110101",
			3132 => "0000000011000011110101",
			3133 => "0001000101101100101000",
			3134 => "0000110101101100100000",
			3135 => "0001001001100000001100",
			3136 => "0000000011000000000100",
			3137 => "0000000011000110001001",
			3138 => "0001001001100100000100",
			3139 => "0000000011000110001001",
			3140 => "0000000011000110001001",
			3141 => "0001011001001000001100",
			3142 => "0010001111011000001000",
			3143 => "0010001111001000000100",
			3144 => "0000000011000110001001",
			3145 => "0000000011000110001001",
			3146 => "0000000011000110001001",
			3147 => "0001010101101100000100",
			3148 => "0000000011000110001001",
			3149 => "0000000011000110001001",
			3150 => "0001101100100000000100",
			3151 => "0000000011000110001001",
			3152 => "0000000011000110001001",
			3153 => "0000011000011000100000",
			3154 => "0001101010011100000100",
			3155 => "0000000011000110001001",
			3156 => "0010101011000000010000",
			3157 => "0001100000100000001000",
			3158 => "0010010101101100000100",
			3159 => "0000000011000110001001",
			3160 => "0000000011000110001001",
			3161 => "0010000101011100000100",
			3162 => "0000000011000110001001",
			3163 => "0000000011000110001001",
			3164 => "0001010000111000001000",
			3165 => "0010110111011100000100",
			3166 => "0000000011000110001001",
			3167 => "0000000011000110001001",
			3168 => "0000000011000110001001",
			3169 => "0000000011000110001001",
			3170 => "0000101110010000110100",
			3171 => "0011000110110100000100",
			3172 => "0000000011001000001101",
			3173 => "0001110101111000011000",
			3174 => "0001010110101100010000",
			3175 => "0000011001100000001000",
			3176 => "0001000001110000000100",
			3177 => "0000000011001000001101",
			3178 => "0000000011001000001101",
			3179 => "0011000101011100000100",
			3180 => "0000000011001000001101",
			3181 => "0000000011001000001101",
			3182 => "0001001100000000000100",
			3183 => "0000000011001000001101",
			3184 => "0000000011001000001101",
			3185 => "0011001001001000010000",
			3186 => "0000100010110100001100",
			3187 => "0010110101011100001000",
			3188 => "0000001110111100000100",
			3189 => "0000000011001000001101",
			3190 => "0000000011001000001101",
			3191 => "0000000011001000001101",
			3192 => "0000000011001000001101",
			3193 => "0001101000111000000100",
			3194 => "0000000011001000001101",
			3195 => "0000000011001000001101",
			3196 => "0001010101101100000100",
			3197 => "0000000011001000001101",
			3198 => "0010010011001000000100",
			3199 => "0000000011001000001101",
			3200 => "0010011000000100000100",
			3201 => "0000000011001000001101",
			3202 => "0000000011001000001101",
			3203 => "0001111000000100101100",
			3204 => "0000101101000100011000",
			3205 => "0010110110001100000100",
			3206 => "1111111011001010101001",
			3207 => "0011100011000100010000",
			3208 => "0000011101000000001100",
			3209 => "0010100110010000000100",
			3210 => "0000010011001010101001",
			3211 => "0010111010100100000100",
			3212 => "0000001011001010101001",
			3213 => "0000001011001010101001",
			3214 => "0000001011001010101001",
			3215 => "0000000011001010101001",
			3216 => "0010001111111100010000",
			3217 => "0000100101001100001100",
			3218 => "0001101001101100000100",
			3219 => "0000000011001010101001",
			3220 => "0000110011001000000100",
			3221 => "0000010011001010101001",
			3222 => "0000000011001010101001",
			3223 => "1111111011001010101001",
			3224 => "1111111011001010101001",
			3225 => "0000100111101000011100",
			3226 => "0000001000101000000100",
			3227 => "1111111011001010101001",
			3228 => "0011001001001000001100",
			3229 => "0000111000101000001000",
			3230 => "0011000011010000000100",
			3231 => "1111111011001010101001",
			3232 => "0000001011001010101001",
			3233 => "1111111011001010101001",
			3234 => "0010100000111100001000",
			3235 => "0010101000000000000100",
			3236 => "0000001011001010101001",
			3237 => "0000010011001010101001",
			3238 => "0000000011001010101001",
			3239 => "0001010101101100000100",
			3240 => "0000000011001010101001",
			3241 => "1111111011001010101001",
			3242 => "0001010110101100111000",
			3243 => "0000110101101100100000",
			3244 => "0001011110011000010000",
			3245 => "0011111001001000000100",
			3246 => "0000000011001101100101",
			3247 => "0000001010100000000100",
			3248 => "0000000011001101100101",
			3249 => "0001101100011100000100",
			3250 => "0000000011001101100101",
			3251 => "0000000011001101100101",
			3252 => "0010100110000000001100",
			3253 => "0010000011001000000100",
			3254 => "0000000011001101100101",
			3255 => "0010000011100100000100",
			3256 => "0000000011001101100101",
			3257 => "0000000011001101100101",
			3258 => "0000000011001101100101",
			3259 => "0011110011010100010100",
			3260 => "0000010111100100000100",
			3261 => "0000000011001101100101",
			3262 => "0011010101011100001000",
			3263 => "0000101001111100000100",
			3264 => "0000000011001101100101",
			3265 => "0000000011001101100101",
			3266 => "0000001001000000000100",
			3267 => "0000000011001101100101",
			3268 => "0000000011001101100101",
			3269 => "0000000011001101100101",
			3270 => "0011001001001000011000",
			3271 => "0011111100001100000100",
			3272 => "0000000011001101100101",
			3273 => "0010000011010000001000",
			3274 => "0000011001100100000100",
			3275 => "0000000011001101100101",
			3276 => "0000000011001101100101",
			3277 => "0011010110110100000100",
			3278 => "0000000011001101100101",
			3279 => "0010110101011100000100",
			3280 => "0000000011001101100101",
			3281 => "0000000011001101100101",
			3282 => "0010001001000100001000",
			3283 => "0001011110010100000100",
			3284 => "0000000011001101100101",
			3285 => "0000000011001101100101",
			3286 => "0001001101101000000100",
			3287 => "0000000011001101100101",
			3288 => "0000000011001101100101",
			3289 => "0011110010000000110000",
			3290 => "0001011010011100101000",
			3291 => "0010000101101100010100",
			3292 => "0011000110110100000100",
			3293 => "0000000011001111001001",
			3294 => "0010001010100100000100",
			3295 => "0000000011001111001001",
			3296 => "0000000011000000000100",
			3297 => "0000000011001111001001",
			3298 => "0000011000011000000100",
			3299 => "0000000011001111001001",
			3300 => "0000000011001111001001",
			3301 => "0001000101101100010000",
			3302 => "0011000111011100000100",
			3303 => "0000000011001111001001",
			3304 => "0000001011111000000100",
			3305 => "0000000011001111001001",
			3306 => "0000000010110100000100",
			3307 => "0000000011001111001001",
			3308 => "0000000011001111001001",
			3309 => "0000000011001111001001",
			3310 => "0010111100101000000100",
			3311 => "0000000011001111001001",
			3312 => "0000000011001111001001",
			3313 => "0000000011001111001001",
			3314 => "0001111000000100101100",
			3315 => "0000101101000100011000",
			3316 => "0010110110001100000100",
			3317 => "1111111011010001100101",
			3318 => "0000011000111100000100",
			3319 => "0000010011010001100101",
			3320 => "0011001010100100000100",
			3321 => "0000000011010001100101",
			3322 => "0010111010100100000100",
			3323 => "0000001011010001100101",
			3324 => "0011111111101000000100",
			3325 => "0000001011010001100101",
			3326 => "0000010011010001100101",
			3327 => "0001001011101100000100",
			3328 => "1111111011010001100101",
			3329 => "0001011100000000001000",
			3330 => "0011111101101100000100",
			3331 => "0000000011010001100101",
			3332 => "0000001011010001100101",
			3333 => "0000001110100100000100",
			3334 => "0000001011010001100101",
			3335 => "1111111011010001100101",
			3336 => "0000100111101000011100",
			3337 => "0000001000101000000100",
			3338 => "1111111011010001100101",
			3339 => "0000111000100000010100",
			3340 => "0011001001001000001100",
			3341 => "0011011011101100000100",
			3342 => "0000001011010001100101",
			3343 => "0001100100000000000100",
			3344 => "0000000011010001100101",
			3345 => "1111111011010001100101",
			3346 => "0010101101001000000100",
			3347 => "0000001011010001100101",
			3348 => "0000010011010001100101",
			3349 => "1111111011010001100101",
			3350 => "0001010101101100000100",
			3351 => "0000000011010001100101",
			3352 => "1111111011010001100101",
			3353 => "0000010111100100110000",
			3354 => "0010110110001100001000",
			3355 => "0000000101000000000100",
			3356 => "0000000011010100000001",
			3357 => "0000000011010100000001",
			3358 => "0001101001011100100100",
			3359 => "0001011010011100011100",
			3360 => "0010101001001100001100",
			3361 => "0000001010100000001000",
			3362 => "0000000011000000000100",
			3363 => "0000000011010100000001",
			3364 => "0000000011010100000001",
			3365 => "0000000011010100000001",
			3366 => "0010000101101100001000",
			3367 => "0010010110000000000100",
			3368 => "0000000011010100000001",
			3369 => "0000000011010100000001",
			3370 => "0010010110000000000100",
			3371 => "0000000011010100000001",
			3372 => "0000000011010100000001",
			3373 => "0011001001001000000100",
			3374 => "0000000011010100000001",
			3375 => "0000000011010100000001",
			3376 => "0000000011010100000001",
			3377 => "0001000101101100010100",
			3378 => "0010111001001000001100",
			3379 => "0011101111011000001000",
			3380 => "0010000101101100000100",
			3381 => "0000000011010100000001",
			3382 => "0000000011010100000001",
			3383 => "0000000011010100000001",
			3384 => "0000001001011000000100",
			3385 => "0000000011010100000001",
			3386 => "0000000011010100000001",
			3387 => "0010001111111100001000",
			3388 => "0010000101011100000100",
			3389 => "0000000011010100000001",
			3390 => "0000000011010100000001",
			3391 => "0000000011010100000001",
			3392 => "0011101010100001000100",
			3393 => "0011000101010100011100",
			3394 => "0001010110101100010100",
			3395 => "0011001011101100000100",
			3396 => "0000000011010111001101",
			3397 => "0011110001010100001100",
			3398 => "0000101101000100001000",
			3399 => "0010101110011000000100",
			3400 => "0000000011010111001101",
			3401 => "0000000011010111001101",
			3402 => "0000000011010111001101",
			3403 => "0000000011010111001101",
			3404 => "0011111111100100000100",
			3405 => "1111111011010111001101",
			3406 => "0000000011010111001101",
			3407 => "0010001001000100011000",
			3408 => "0001000101010100010000",
			3409 => "0001110101111000000100",
			3410 => "0000000011010111001101",
			3411 => "0001111000111000000100",
			3412 => "0000000011010111001101",
			3413 => "0010101111011100000100",
			3414 => "0000000011010111001101",
			3415 => "0000000011010111001101",
			3416 => "0000100100011100000100",
			3417 => "0000001011010111001101",
			3418 => "0000000011010111001101",
			3419 => "0001000101101100001100",
			3420 => "0000000001101100001000",
			3421 => "0000001011000000000100",
			3422 => "0000000011010111001101",
			3423 => "0000000011010111001101",
			3424 => "0000000011010111001101",
			3425 => "0000000011010111001101",
			3426 => "0010101000111000010000",
			3427 => "0011000011010000001000",
			3428 => "0011011101000000000100",
			3429 => "0000000011010111001101",
			3430 => "1111111011010111001101",
			3431 => "0011110100001100000100",
			3432 => "0000000011010111001101",
			3433 => "0000000011010111001101",
			3434 => "0010000011010000001000",
			3435 => "0001010100101100000100",
			3436 => "0000000011010111001101",
			3437 => "0000000011010111001101",
			3438 => "0011001001001000000100",
			3439 => "1111111011010111001101",
			3440 => "0000000100100000000100",
			3441 => "0000000011010111001101",
			3442 => "0000000011010111001101",
			3443 => "0011100010011101000000",
			3444 => "0011001001001000100100",
			3445 => "0000111001010000100000",
			3446 => "0010001001001100001100",
			3447 => "0001101001101100001000",
			3448 => "0000100000111000000100",
			3449 => "0000000011011001100001",
			3450 => "0000000011011001100001",
			3451 => "0000001011011001100001",
			3452 => "0011001010100100000100",
			3453 => "1111111011011001100001",
			3454 => "0001100011000100001000",
			3455 => "0010100110110100000100",
			3456 => "0000000011011001100001",
			3457 => "0000000011011001100001",
			3458 => "0010011001000100000100",
			3459 => "0000000011011001100001",
			3460 => "0000000011011001100001",
			3461 => "1111111011011001100001",
			3462 => "0001101000111000001000",
			3463 => "0001111111011000000100",
			3464 => "0000000011011001100001",
			3465 => "0000000011011001100001",
			3466 => "0010101100010000001000",
			3467 => "0000000111001000000100",
			3468 => "0000000011011001100001",
			3469 => "0000000011011001100001",
			3470 => "0000111000100000001000",
			3471 => "0000000100100000000100",
			3472 => "0000001011011001100001",
			3473 => "0000000011011001100001",
			3474 => "0000000011011001100001",
			3475 => "0010101010000100000100",
			3476 => "0000000011011001100001",
			3477 => "0011001001010100000100",
			3478 => "1111111011011001100001",
			3479 => "0000000011011001100001",
			3480 => "0001111000000100101000",
			3481 => "0011001011101100000100",
			3482 => "0000000011011100100101",
			3483 => "0001011001010100011100",
			3484 => "0010101110011000001100",
			3485 => "0000001010100000001000",
			3486 => "0001111001001000000100",
			3487 => "0000000011011100100101",
			3488 => "0000000011011100100101",
			3489 => "0000000011011100100101",
			3490 => "0010010110000000001000",
			3491 => "0000011000011000000100",
			3492 => "0000000011011100100101",
			3493 => "0000000011011100100101",
			3494 => "0000001101000100000100",
			3495 => "0000000011011100100101",
			3496 => "0000000011011100100101",
			3497 => "0010111010100100000100",
			3498 => "0000000011011100100101",
			3499 => "0000000011011100100101",
			3500 => "0011001001001000011100",
			3501 => "0010000011010000001000",
			3502 => "0001010001010000000100",
			3503 => "0000000011011100100101",
			3504 => "0000000011011100100101",
			3505 => "0010100011001000010000",
			3506 => "0000110101101100001000",
			3507 => "0000110001100100000100",
			3508 => "0000000011011100100101",
			3509 => "0000000011011100100101",
			3510 => "0010000101011100000100",
			3511 => "0000000011011100100101",
			3512 => "0000000011011100100101",
			3513 => "0000000011011100100101",
			3514 => "0000010111100100010000",
			3515 => "0000111000000000001000",
			3516 => "0001011101000000000100",
			3517 => "0000000011011100100101",
			3518 => "0000000011011100100101",
			3519 => "0000111110111000000100",
			3520 => "0000000011011100100101",
			3521 => "0000000011011100100101",
			3522 => "0010011011111000001000",
			3523 => "0001111000000000000100",
			3524 => "0000000011011100100101",
			3525 => "0000000011011100100101",
			3526 => "0000111100101100000100",
			3527 => "0000000011011100100101",
			3528 => "0000000011011100100101",
			3529 => "0011001011101100000100",
			3530 => "0000000011011110101001",
			3531 => "0010001111111100100000",
			3532 => "0001011010011100011000",
			3533 => "0011110011010100010100",
			3534 => "0010101110011000001100",
			3535 => "0000001010100000001000",
			3536 => "0000001000000100000100",
			3537 => "0000000011011110101001",
			3538 => "0000000011011110101001",
			3539 => "0000000011011110101001",
			3540 => "0001010111011100000100",
			3541 => "0000000011011110101001",
			3542 => "0000000011011110101001",
			3543 => "0000000011011110101001",
			3544 => "0010110101011100000100",
			3545 => "0000000011011110101001",
			3546 => "0000000011011110101001",
			3547 => "0010110101011100010000",
			3548 => "0011100011000100001100",
			3549 => "0001111001000100000100",
			3550 => "0000000011011110101001",
			3551 => "0000001001000000000100",
			3552 => "0000000011011110101001",
			3553 => "0000000011011110101001",
			3554 => "0000000011011110101001",
			3555 => "0000101110010000001100",
			3556 => "0001101000111000001000",
			3557 => "0001111111011000000100",
			3558 => "0000000011011110101001",
			3559 => "0000000011011110101001",
			3560 => "0000000011011110101001",
			3561 => "0000000011011110101001",
			3562 => "0001111000000100110100",
			3563 => "0000101101101100011000",
			3564 => "0010110110001100000100",
			3565 => "1111111011100001000101",
			3566 => "0001010011001000010000",
			3567 => "0010001001001100000100",
			3568 => "0000001011100001000101",
			3569 => "0001101101101000000100",
			3570 => "0000001011100001000101",
			3571 => "0001111100101000000100",
			3572 => "0000001011100001000101",
			3573 => "0000001011100001000101",
			3574 => "0000000011100001000101",
			3575 => "0000011000011000010100",
			3576 => "0000100101001100010000",
			3577 => "0010101010100100000100",
			3578 => "1111111011100001000101",
			3579 => "0001000110101100001000",
			3580 => "0011000111011100000100",
			3581 => "0000001011100001000101",
			3582 => "0000001011100001000101",
			3583 => "1111111011100001000101",
			3584 => "1111111011100001000101",
			3585 => "0010110101010100000100",
			3586 => "1111111011100001000101",
			3587 => "0000000011100001000101",
			3588 => "0000100000001100011000",
			3589 => "0000001000101000000100",
			3590 => "1111111011100001000101",
			3591 => "0001001011111000010000",
			3592 => "0011000011010000000100",
			3593 => "1111111011100001000101",
			3594 => "0011011110011000000100",
			3595 => "0000001011100001000101",
			3596 => "0000000010110100000100",
			3597 => "0000001011100001000101",
			3598 => "0000000011100001000101",
			3599 => "1111111011100001000101",
			3600 => "1111111011100001000101",
			3601 => "0001111000000100110000",
			3602 => "0011001011101100000100",
			3603 => "0000000011100100011001",
			3604 => "0000010111100100011000",
			3605 => "0010101110011000001000",
			3606 => "0000001010100000000100",
			3607 => "0000000011100100011001",
			3608 => "0000000011100100011001",
			3609 => "0001010001011000001100",
			3610 => "0010000101101100001000",
			3611 => "0000100101001100000100",
			3612 => "0000000011100100011001",
			3613 => "0000000011100100011001",
			3614 => "0000000011100100011001",
			3615 => "0000000011100100011001",
			3616 => "0010110111011100001000",
			3617 => "0001011000000000000100",
			3618 => "0000000011100100011001",
			3619 => "0000000011100100011001",
			3620 => "0010000000110000001000",
			3621 => "0000000001101100000100",
			3622 => "0000000011100100011001",
			3623 => "0000000011100100011001",
			3624 => "0000000011100100011001",
			3625 => "0011001001001000011100",
			3626 => "0010000011010000001000",
			3627 => "0001010001010000000100",
			3628 => "0000000011100100011001",
			3629 => "0000000011100100011001",
			3630 => "0010100011001000010000",
			3631 => "0000110101101100001000",
			3632 => "0000110001100100000100",
			3633 => "0000000011100100011001",
			3634 => "0000000011100100011001",
			3635 => "0010000101011100000100",
			3636 => "0000000011100100011001",
			3637 => "0000000011100100011001",
			3638 => "0000000011100100011001",
			3639 => "0000010111100100010000",
			3640 => "0000111000000000001000",
			3641 => "0001111100110000000100",
			3642 => "0000000011100100011001",
			3643 => "0000000011100100011001",
			3644 => "0000111110111000000100",
			3645 => "0000000011100100011001",
			3646 => "0000000011100100011001",
			3647 => "0010011011111000001000",
			3648 => "0001111000000000000100",
			3649 => "0000000011100100011001",
			3650 => "0000000011100100011001",
			3651 => "0000111100101100000100",
			3652 => "0000000011100100011001",
			3653 => "0000000011100100011001",
			3654 => "0011101111100000111100",
			3655 => "0010001001000100100100",
			3656 => "0010110110001100000100",
			3657 => "0000000011100111011101",
			3658 => "0000100100011100011000",
			3659 => "0010100101011100001100",
			3660 => "0000000010001100001000",
			3661 => "0000000011000000000100",
			3662 => "0000000011100111011101",
			3663 => "0000000011100111011101",
			3664 => "0000000011100111011101",
			3665 => "0000011000011000001000",
			3666 => "0001001111101000000100",
			3667 => "0000001011100111011101",
			3668 => "0000000011100111011101",
			3669 => "0000000011100111011101",
			3670 => "0011100001010100000100",
			3671 => "0000000011100111011101",
			3672 => "0000000011100111011101",
			3673 => "0001000101101100010100",
			3674 => "0010100011000000010000",
			3675 => "0001010011010000001100",
			3676 => "0000000110100000001000",
			3677 => "0000001011000000000100",
			3678 => "0000000011100111011101",
			3679 => "0000000011100111011101",
			3680 => "0000000011100111011101",
			3681 => "0000000011100111011101",
			3682 => "0000000011100111011101",
			3683 => "0000000011100111011101",
			3684 => "0010101000111000010000",
			3685 => "0011000011010000001000",
			3686 => "0011011111011100000100",
			3687 => "0000000011100111011101",
			3688 => "0000000011100111011101",
			3689 => "0011110100001100000100",
			3690 => "0000000011100111011101",
			3691 => "0000000011100111011101",
			3692 => "0010010001001000010100",
			3693 => "0010000011010000001000",
			3694 => "0011010110110100000100",
			3695 => "0000000011100111011101",
			3696 => "0000000011100111011101",
			3697 => "0011001001001000000100",
			3698 => "1111111011100111011101",
			3699 => "0011000101101100000100",
			3700 => "0000000011100111011101",
			3701 => "0000000011100111011101",
			3702 => "0000000011100111011101",
			3703 => "0000010000011000100000",
			3704 => "0000110101101100001100",
			3705 => "0001011110011000001000",
			3706 => "0011000111011100000100",
			3707 => "0000000011101010110001",
			3708 => "0000000011101010110001",
			3709 => "0000000011101010110001",
			3710 => "0011110001010100000100",
			3711 => "0000000011101010110001",
			3712 => "0011100000100000001100",
			3713 => "0001001011111000001000",
			3714 => "0000101101010000000100",
			3715 => "0000000011101010110001",
			3716 => "0000000011101010110001",
			3717 => "0000000011101010110001",
			3718 => "0000000011101010110001",
			3719 => "0011101001000000100100",
			3720 => "0010111010100100001000",
			3721 => "0001000110110100000100",
			3722 => "0000000011101010110001",
			3723 => "0000000011101010110001",
			3724 => "0010111010000100001100",
			3725 => "0000101111110000001000",
			3726 => "0000001000111000000100",
			3727 => "0000000011101010110001",
			3728 => "0000000011101010110001",
			3729 => "0000000011101010110001",
			3730 => "0010001111011000000100",
			3731 => "0000000011101010110001",
			3732 => "0000111100101000001000",
			3733 => "0000110101010100000100",
			3734 => "0000000011101010110001",
			3735 => "0000000011101010110001",
			3736 => "0000000011101010110001",
			3737 => "0011001001001000010000",
			3738 => "0010000011010000000100",
			3739 => "0000000011101010110001",
			3740 => "0001011000000100001000",
			3741 => "0001010011001000000100",
			3742 => "0000000011101010110001",
			3743 => "0000000011101010110001",
			3744 => "1111111011101010110001",
			3745 => "0010100000111100010100",
			3746 => "0010101000101000001000",
			3747 => "0001110001001000000100",
			3748 => "0000000011101010110001",
			3749 => "0000000011101010110001",
			3750 => "0001111100101100000100",
			3751 => "0000000011101010110001",
			3752 => "0001110011110100000100",
			3753 => "0000000011101010110001",
			3754 => "0000000011101010110001",
			3755 => "0000000011101010110001",
			3756 => "0000100000001101000000",
			3757 => "0011000011010000010100",
			3758 => "0000000000111000001000",
			3759 => "0010110110001100000100",
			3760 => "0000000011101100110101",
			3761 => "0000000011101100110101",
			3762 => "0010000011010000000100",
			3763 => "0000000011101100110101",
			3764 => "0000000100110000000100",
			3765 => "0000000011101100110101",
			3766 => "0000000011101100110101",
			3767 => "0001010000111000101000",
			3768 => "0010101111111100010000",
			3769 => "0000001101000100001000",
			3770 => "0000001000111000000100",
			3771 => "0000000011101100110101",
			3772 => "0000000011101100110101",
			3773 => "0000010011110000000100",
			3774 => "0000000011101100110101",
			3775 => "0000000011101100110101",
			3776 => "0000011000011000001100",
			3777 => "0010001001000100001000",
			3778 => "0001010011000000000100",
			3779 => "0000000011101100110101",
			3780 => "0000000011101100110101",
			3781 => "0000000011101100110101",
			3782 => "0001011111101000001000",
			3783 => "0000001110100100000100",
			3784 => "0000000011101100110101",
			3785 => "0000000011101100110101",
			3786 => "0000000011101100110101",
			3787 => "0000000011101100110101",
			3788 => "0000000011101100110101",
			3789 => "0011100000100001000100",
			3790 => "0001001110011000011000",
			3791 => "0011000110110100000100",
			3792 => "1111111011101111000001",
			3793 => "0000101010000100000100",
			3794 => "0000000011101111000001",
			3795 => "0000101111100000000100",
			3796 => "0000001011101111000001",
			3797 => "0000111100101000001000",
			3798 => "0001101110010100000100",
			3799 => "1111111011101111000001",
			3800 => "0000000011101111000001",
			3801 => "0000001011101111000001",
			3802 => "0010001001000100011100",
			3803 => "0011001001001000010100",
			3804 => "0011101000100000001000",
			3805 => "0010111010100100000100",
			3806 => "0000000011101111000001",
			3807 => "0000001011101111000001",
			3808 => "0000011000111100000100",
			3809 => "0000000011101111000001",
			3810 => "0011110101001000000100",
			3811 => "1111111011101111000001",
			3812 => "0000000011101111000001",
			3813 => "0011000101101100000100",
			3814 => "0000001011101111000001",
			3815 => "1111111011101111000001",
			3816 => "0001000101101100001100",
			3817 => "0010101000000000001000",
			3818 => "0000011001100000000100",
			3819 => "0000000011101111000001",
			3820 => "0000000011101111000001",
			3821 => "0000000011101111000001",
			3822 => "1111111011101111000001",
			3823 => "1111111011101111000001",
			3824 => "0000100000001100110100",
			3825 => "0001011010011100101100",
			3826 => "0001010001001000101000",
			3827 => "0000010111100100010100",
			3828 => "0010110110001100000100",
			3829 => "1111111011110000101101",
			3830 => "0000101101000100001000",
			3831 => "0000000011000000000100",
			3832 => "0000000011110000101101",
			3833 => "0000001011110000101101",
			3834 => "0011111101101100000100",
			3835 => "0000000011110000101101",
			3836 => "0000000011110000101101",
			3837 => "0001000101101100001100",
			3838 => "0010101000000000001000",
			3839 => "0001011110011000000100",
			3840 => "0000000011110000101101",
			3841 => "0000000011110000101101",
			3842 => "0000001011110000101101",
			3843 => "0001000110000000000100",
			3844 => "0000000011110000101101",
			3845 => "1111111011110000101101",
			3846 => "0000001011110000101101",
			3847 => "0010010101111000000100",
			3848 => "1111111011110000101101",
			3849 => "0000000011110000101101",
			3850 => "1111111011110000101101",
			3851 => "0011100010011101010000",
			3852 => "0010110101011100110000",
			3853 => "0010011101101000101000",
			3854 => "0011000101010100011000",
			3855 => "0001010110101100010000",
			3856 => "0011001011101100001000",
			3857 => "0001101111011000000100",
			3858 => "0000000011110011011001",
			3859 => "0000000011110011011001",
			3860 => "0010000101101100000100",
			3861 => "0000000011110011011001",
			3862 => "0000000011110011011001",
			3863 => "0000010001110000000100",
			3864 => "0000000011110011011001",
			3865 => "0000000011110011011001",
			3866 => "0000000001111000001100",
			3867 => "0000111100101000001000",
			3868 => "0000000010000000000100",
			3869 => "0000000011110011011001",
			3870 => "0000000011110011011001",
			3871 => "0000000011110011011001",
			3872 => "0000000011110011011001",
			3873 => "0011001001001000000100",
			3874 => "0000000011110011011001",
			3875 => "0000000011110011011001",
			3876 => "0000010111100100001100",
			3877 => "0010100101011100001000",
			3878 => "0001011101000000000100",
			3879 => "0000000011110011011001",
			3880 => "0000000011110011011001",
			3881 => "0000000011110011011001",
			3882 => "0000000011101100001100",
			3883 => "0001101000111000001000",
			3884 => "0001111111011000000100",
			3885 => "0000000011110011011001",
			3886 => "0000000011110011011001",
			3887 => "0000000011110011011001",
			3888 => "0001111001010100000100",
			3889 => "0000000011110011011001",
			3890 => "0000000011110011011001",
			3891 => "0010001011000000000100",
			3892 => "1111111011110011011001",
			3893 => "0000000011110011011001",
			3894 => "0011110010000000111000",
			3895 => "0010101001011000110100",
			3896 => "0010000101101100011000",
			3897 => "0010101011000000010100",
			3898 => "0001010001011000010000",
			3899 => "0000000101000000001000",
			3900 => "0001111000000100000100",
			3901 => "0000000011110101001101",
			3902 => "1111111011110101001101",
			3903 => "0001100101110000000100",
			3904 => "0000000011110101001101",
			3905 => "0000001011110101001101",
			3906 => "0000000011110101001101",
			3907 => "0000001011110101001101",
			3908 => "0010110101011100001100",
			3909 => "0001100011001000001000",
			3910 => "0011101010100100000100",
			3911 => "0000000011110101001101",
			3912 => "0000000011110101001101",
			3913 => "1111111011110101001101",
			3914 => "0001101000111000001000",
			3915 => "0001111111011000000100",
			3916 => "0000000011110101001101",
			3917 => "0000000011110101001101",
			3918 => "0000000010110100000100",
			3919 => "0000001011110101001101",
			3920 => "0000000011110101001101",
			3921 => "1111111011110101001101",
			3922 => "1111111011110101001101",
			3923 => "0000100101001101010000",
			3924 => "0011001001001000111000",
			3925 => "0010000101101100101000",
			3926 => "0000101101000100010000",
			3927 => "0010110110001100000100",
			3928 => "0000000011110111110001",
			3929 => "0000010111100100001000",
			3930 => "0000110110001100000100",
			3931 => "0000000011110111110001",
			3932 => "0000001011110111110001",
			3933 => "0000000011110111110001",
			3934 => "0000000101000000010000",
			3935 => "0001001110011000001000",
			3936 => "0000010001110000000100",
			3937 => "0000000011110111110001",
			3938 => "0000000011110111110001",
			3939 => "0010101111101000000100",
			3940 => "0000000011110111110001",
			3941 => "0000000011110111110001",
			3942 => "0011011011101100000100",
			3943 => "0000000011110111110001",
			3944 => "0000000011110111110001",
			3945 => "0001100011001000001000",
			3946 => "0000001000101000000100",
			3947 => "0000000011110111110001",
			3948 => "0000000011110111110001",
			3949 => "0001000110001100000100",
			3950 => "0000000011110111110001",
			3951 => "0000000011110111110001",
			3952 => "0001101000111000001000",
			3953 => "0001111111011000000100",
			3954 => "0000000011110111110001",
			3955 => "0000000011110111110001",
			3956 => "0010101100010000001000",
			3957 => "0000001101100100000100",
			3958 => "0000000011110111110001",
			3959 => "0000000011110111110001",
			3960 => "0000000010000000000100",
			3961 => "0000000011110111110001",
			3962 => "0000001011110111110001",
			3963 => "1111111011110111110001",
			3964 => "0000100000001100111000",
			3965 => "0000101010000100000100",
			3966 => "1111111011111001100101",
			3967 => "0001000101101100011000",
			3968 => "0011000110110100000100",
			3969 => "1111111011111001100101",
			3970 => "0001101111000100010000",
			3971 => "0000101111100000001000",
			3972 => "0010011100110000000100",
			3973 => "0000001011111001100101",
			3974 => "1111111011111001100101",
			3975 => "0010101010100100000100",
			3976 => "1111111011111001100101",
			3977 => "0000001011111001100101",
			3978 => "1111111011111001100101",
			3979 => "0010001001000100010100",
			3980 => "0011001100101000001100",
			3981 => "0001011010011100001000",
			3982 => "0011000011010000000100",
			3983 => "0000000011111001100101",
			3984 => "0000001011111001100101",
			3985 => "1111111011111001100101",
			3986 => "0001010010111000000100",
			3987 => "0000001011111001100101",
			3988 => "1111111011111001100101",
			3989 => "0010010011001000000100",
			3990 => "1111111011111001100101",
			3991 => "1111111011111001100101",
			3992 => "1111111011111001100101",
			3993 => "0011100000100001000000",
			3994 => "0010001111111100100000",
			3995 => "0001011010011100011100",
			3996 => "0011000110110100000100",
			3997 => "1111111011111011101001",
			3998 => "0011110001010100010000",
			3999 => "0000100000111000001000",
			4000 => "0000000011000000000100",
			4001 => "0000000011111011101001",
			4002 => "0000001011111011101001",
			4003 => "0011000111011100000100",
			4004 => "0000000011111011101001",
			4005 => "0000000011111011101001",
			4006 => "0010111011101100000100",
			4007 => "0000000011111011101001",
			4008 => "0000001011111011101001",
			4009 => "1111111011111011101001",
			4010 => "0010111010100100000100",
			4011 => "1111111011111011101001",
			4012 => "0001111111011000001000",
			4013 => "0011101001011000000100",
			4014 => "0000001011111011101001",
			4015 => "0000000011111011101001",
			4016 => "0011001001001000001000",
			4017 => "0010101001100000000100",
			4018 => "0000000011111011101001",
			4019 => "1111111011111011101001",
			4020 => "0001101100010000000100",
			4021 => "1111111011111011101001",
			4022 => "0000101110010000000100",
			4023 => "0000000011111011101001",
			4024 => "0000000011111011101001",
			4025 => "1111111011111011101001",
			4026 => "0011100000100000111100",
			4027 => "0001010000111000111000",
			4028 => "0000010111100100011000",
			4029 => "0000101111100000001000",
			4030 => "0000000011000000000100",
			4031 => "1111111011111101100101",
			4032 => "0000001011111101100101",
			4033 => "0001010101010100000100",
			4034 => "1111111011111101100101",
			4035 => "0001001110011000000100",
			4036 => "0000001011111101100101",
			4037 => "0010110101011100000100",
			4038 => "0000000011111101100101",
			4039 => "0000001011111101100101",
			4040 => "0011000101010100001000",
			4041 => "0001000110001100000100",
			4042 => "0000000011111101100101",
			4043 => "1111111011111101100101",
			4044 => "0001111100000000001000",
			4045 => "0000000001101100000100",
			4046 => "0000001011111101100101",
			4047 => "1111111011111101100101",
			4048 => "0011101111100000001000",
			4049 => "0010101000111000000100",
			4050 => "1111111011111101100101",
			4051 => "0000000011111101100101",
			4052 => "0001011100101100000100",
			4053 => "0000001011111101100101",
			4054 => "1111111011111101100101",
			4055 => "1111111011111101100101",
			4056 => "1111111011111101100101",
			4057 => "0000100101001101001000",
			4058 => "0001111000000100101100",
			4059 => "0011000101010100100000",
			4060 => "0000010111100100011000",
			4061 => "0000101101000100001100",
			4062 => "0010110110001100000100",
			4063 => "1111111011111111111001",
			4064 => "0000000001101000000100",
			4065 => "0000001011111111111001",
			4066 => "0000001011111111111001",
			4067 => "0001101001101100000100",
			4068 => "1111111011111111111001",
			4069 => "0001011010011100000100",
			4070 => "0000000011111111111001",
			4071 => "0000000011111111111001",
			4072 => "0001101000000000000100",
			4073 => "0000000011111111111001",
			4074 => "1111111011111111111001",
			4075 => "0000101111110000001000",
			4076 => "0010100110001100000100",
			4077 => "0000000011111111111001",
			4078 => "0000001011111111111001",
			4079 => "0000000011111111111001",
			4080 => "0000001000101000000100",
			4081 => "1111111011111111111001",
			4082 => "0001000100101100010100",
			4083 => "0010011001001000000100",
			4084 => "1111111011111111111001",
			4085 => "0011111010100000001000",
			4086 => "0000001101100100000100",
			4087 => "0000000011111111111001",
			4088 => "1111111011111111111001",
			4089 => "0010110101011100000100",
			4090 => "0000000011111111111001",
			4091 => "0000001011111111111001",
			4092 => "1111111011111111111001",
			4093 => "1111111011111111111001",
			4094 => "0000100000001101000000",
			4095 => "0000101010000100000100",
			4096 => "1111111100000001111101",
			4097 => "0001010110101100100000",
			4098 => "0000000000110100010000",
			4099 => "0010110110001100000100",
			4100 => "1111111100000001111101",
			4101 => "0000011000111100000100",
			4102 => "0000001100000001111101",
			4103 => "0010111010100100000100",
			4104 => "0000000100000001111101",
			4105 => "0000001100000001111101",
			4106 => "0011110111010100000100",
			4107 => "1111111100000001111101",
			4108 => "0001101111000100001000",
			4109 => "0010001111111100000100",
			4110 => "0000001100000001111101",
			4111 => "0000000100000001111101",
			4112 => "1111111100000001111101",
			4113 => "0010001001000100010000",
			4114 => "0011001100101000001000",
			4115 => "0001011010011100000100",
			4116 => "0000000100000001111101",
			4117 => "1111111100000001111101",
			4118 => "0001000011000100000100",
			4119 => "0000001100000001111101",
			4120 => "1111111100000001111101",
			4121 => "0001111000000100000100",
			4122 => "1111111100000001111101",
			4123 => "0001111101001000000100",
			4124 => "1111111100000001111101",
			4125 => "1111111100000001111101",
			4126 => "1111111100000001111101",
			4127 => "0000100000001101001000",
			4128 => "0011001001001000110000",
			4129 => "0000111001010000101100",
			4130 => "0010001001001100001100",
			4131 => "0001101001101100001000",
			4132 => "0000100000111000000100",
			4133 => "0000000100000100010001",
			4134 => "0000000100000100010001",
			4135 => "0000000100000100010001",
			4136 => "0001100011000100010000",
			4137 => "0010111010100100001000",
			4138 => "0011100011001000000100",
			4139 => "0000000100000100010001",
			4140 => "0000000100000100010001",
			4141 => "0000001000111000000100",
			4142 => "0000000100000100010001",
			4143 => "0000001100000100010001",
			4144 => "0000000101000000001000",
			4145 => "0001111111011000000100",
			4146 => "1111111100000100010001",
			4147 => "0000000100000100010001",
			4148 => "0011100111010100000100",
			4149 => "0000000100000100010001",
			4150 => "0000000100000100010001",
			4151 => "1111111100000100010001",
			4152 => "0001101000111000001000",
			4153 => "0001111111011000000100",
			4154 => "0000000100000100010001",
			4155 => "0000000100000100010001",
			4156 => "0000110001001000001100",
			4157 => "0010101100010000001000",
			4158 => "0000000111001000000100",
			4159 => "0000000100000100010001",
			4160 => "0000000100000100010001",
			4161 => "0000001100000100010001",
			4162 => "0000000100000100010001",
			4163 => "1111111100000100010001",
			4164 => "0011100000100001001000",
			4165 => "0010001001000100101000",
			4166 => "0001010000111000100100",
			4167 => "0010101011000000011100",
			4168 => "0010001001001100010000",
			4169 => "0001101001000000001000",
			4170 => "0001101100000000000100",
			4171 => "0000000100000110100101",
			4172 => "0000000100000110100101",
			4173 => "0000101101010000000100",
			4174 => "0000001100000110100101",
			4175 => "0000000100000110100101",
			4176 => "0011001010100100000100",
			4177 => "0000000100000110100101",
			4178 => "0011100011000100000100",
			4179 => "0000000100000110100101",
			4180 => "0000000100000110100101",
			4181 => "0010110111011100000100",
			4182 => "0000000100000110100101",
			4183 => "0000001100000110100101",
			4184 => "0000000100000110100101",
			4185 => "0001000101101100011100",
			4186 => "0010111001001000010000",
			4187 => "0001101111101000001100",
			4188 => "0000100110011100001000",
			4189 => "0010101111011100000100",
			4190 => "0000000100000110100101",
			4191 => "0000000100000110100101",
			4192 => "0000000100000110100101",
			4193 => "0000000100000110100101",
			4194 => "0000001001011000000100",
			4195 => "0000000100000110100101",
			4196 => "0000000100110000000100",
			4197 => "0000000100000110100101",
			4198 => "0000000100000110100101",
			4199 => "1111111100000110100101",
			4200 => "1111111100000110100101",
			4201 => "0011100000100001010000",
			4202 => "0011001001001000110000",
			4203 => "0001010011110100101100",
			4204 => "0010001111111100011100",
			4205 => "0000110101101100001100",
			4206 => "0001011110011000001000",
			4207 => "0011000111011100000100",
			4208 => "0000000100001001001001",
			4209 => "0000000100001001001001",
			4210 => "0000000100001001001001",
			4211 => "0011110111010100001000",
			4212 => "0011101000100000000100",
			4213 => "0000000100001001001001",
			4214 => "0000000100001001001001",
			4215 => "0000000000000100000100",
			4216 => "0000001100001001001001",
			4217 => "0000000100001001001001",
			4218 => "0011101010011100001100",
			4219 => "0011000011010000000100",
			4220 => "0000000100001001001001",
			4221 => "0010001001000100000100",
			4222 => "0000000100001001001001",
			4223 => "0000000100001001001001",
			4224 => "0000000100001001001001",
			4225 => "0000000100001001001001",
			4226 => "0000010111100100010000",
			4227 => "0010101000000000001100",
			4228 => "0011000101101100001000",
			4229 => "0001001000011000000100",
			4230 => "0000000100001001001001",
			4231 => "0000000100001001001001",
			4232 => "0000000100001001001001",
			4233 => "0000000100001001001001",
			4234 => "0000000010110100001100",
			4235 => "0001101000111000001000",
			4236 => "0001111111011000000100",
			4237 => "0000000100001001001001",
			4238 => "0000000100001001001001",
			4239 => "0000000100001001001001",
			4240 => "0000000100001001001001",
			4241 => "0000000100001001001001",
			4242 => "0011100000100001000100",
			4243 => "0010101001011001000000",
			4244 => "0010001001001100010000",
			4245 => "0010110110001100000100",
			4246 => "0000000100001011010111",
			4247 => "0010011100101000000100",
			4248 => "0000001100001011010111",
			4249 => "0000111111011000000100",
			4250 => "0000000100001011010111",
			4251 => "0000000100001011010111",
			4252 => "0011000111011100010100",
			4253 => "0000000100011100010000",
			4254 => "0011101101001000001000",
			4255 => "0001110111011100000100",
			4256 => "0000000100001011010111",
			4257 => "0000000100001011010111",
			4258 => "0001111111011000000100",
			4259 => "1111111100001011010111",
			4260 => "0000000100001011010111",
			4261 => "0000000100001011010111",
			4262 => "0000000001101100010000",
			4263 => "0001101000111000001000",
			4264 => "0001111111011000000100",
			4265 => "0000000100001011010111",
			4266 => "1111111100001011010111",
			4267 => "0010101111111100000100",
			4268 => "0000000100001011010111",
			4269 => "0000001100001011010111",
			4270 => "0011111101101100000100",
			4271 => "1111111100001011010111",
			4272 => "0011001001001000000100",
			4273 => "0000000100001011010111",
			4274 => "0000001100001011010111",
			4275 => "1111111100001011010111",
			4276 => "1111111100001011010111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1469, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2865, initial_addr_3'length));
	end generate gen_rom_11;

	gen_rom_12: if SELECT_ROM = 12 generate
		bank <= (
			0 => "0000001000111000000100",
			1 => "0000001000000000001101",
			2 => "1111111000000000001101",
			3 => "0000001000111000000100",
			4 => "0000000000000000011001",
			5 => "0000000000000000011001",
			6 => "0000001000111000001000",
			7 => "0010000101011100000100",
			8 => "0000001000000000101101",
			9 => "0000010000000000101101",
			10 => "1111111000000000101101",
			11 => "0000001000111000001000",
			12 => "0010000101011100000100",
			13 => "0000000000000001000001",
			14 => "0000001000000001000001",
			15 => "1111111000000001000001",
			16 => "0000001000111000001000",
			17 => "0001010001100100000100",
			18 => "0000000000000001010101",
			19 => "0000001000000001010101",
			20 => "1111111000000001010101",
			21 => "0000001000111000001000",
			22 => "0010110101010100000100",
			23 => "0000000000000001101001",
			24 => "0000001000000001101001",
			25 => "1111111000000001101001",
			26 => "0000001000111000001000",
			27 => "0010000101011100000100",
			28 => "0000000000000001111101",
			29 => "0000001000000001111101",
			30 => "1111111000000001111101",
			31 => "0000001000111000001000",
			32 => "0010000101011100000100",
			33 => "0000000000000010010001",
			34 => "0000000000000010010001",
			35 => "1111111000000010010001",
			36 => "0000101000000100001000",
			37 => "0000111001100000000100",
			38 => "0000000000000010100101",
			39 => "0000000000000010100101",
			40 => "0000000000000010100101",
			41 => "0000001000111000001000",
			42 => "0010000101011100000100",
			43 => "0000000000000010111001",
			44 => "0000000000000010111001",
			45 => "0000000000000010111001",
			46 => "0000101000000100001000",
			47 => "0010101000011000000100",
			48 => "0000000000000011001101",
			49 => "0000000000000011001101",
			50 => "0000000000000011001101",
			51 => "0000001000111000001000",
			52 => "0010101000011000000100",
			53 => "0000000000000011100001",
			54 => "0000000000000011100001",
			55 => "0000000000000011100001",
			56 => "0000001000111000001000",
			57 => "0010110101010100000100",
			58 => "0000000000000011110101",
			59 => "0000000000000011110101",
			60 => "0000000000000011110101",
			61 => "0000001000111000001000",
			62 => "0010000101011100000100",
			63 => "0000000000000100001001",
			64 => "0000000000000100001001",
			65 => "0000000000000100001001",
			66 => "0000001000111000001000",
			67 => "0010000101011100000100",
			68 => "0000000000000100011101",
			69 => "0000000000000100011101",
			70 => "0000000000000100011101",
			71 => "0000001000111000001000",
			72 => "0010000101011100000100",
			73 => "0000000000000100110001",
			74 => "0000000000000100110001",
			75 => "0000000000000100110001",
			76 => "0000001000111000001000",
			77 => "0010101000011000000100",
			78 => "0000000000000101000101",
			79 => "0000000000000101000101",
			80 => "0000000000000101000101",
			81 => "0000001000111000001000",
			82 => "0010000101011100000100",
			83 => "0000000000000101011001",
			84 => "0000000000000101011001",
			85 => "0000000000000101011001",
			86 => "0000001000111000001000",
			87 => "0000100011000000000100",
			88 => "1110111000000101101101",
			89 => "1110110000000101101101",
			90 => "1110001000000101101101",
			91 => "0000001000000100001000",
			92 => "0010000101011100000100",
			93 => "0000001000000110001001",
			94 => "0000001000000110001001",
			95 => "0000001101001000000100",
			96 => "0000000000000110001001",
			97 => "1111111000000110001001",
			98 => "0000001000000100000100",
			99 => "0000001000000110100101",
			100 => "0010011100101100000100",
			101 => "1111111000000110100101",
			102 => "0010111000111000000100",
			103 => "0000000000000110100101",
			104 => "1111111000000110100101",
			105 => "0000101010000100000100",
			106 => "0000001000000111000001",
			107 => "0010110011001000000100",
			108 => "1111111000000111000001",
			109 => "0000001001111100000100",
			110 => "0000001000000111000001",
			111 => "1111111000000111000001",
			112 => "0000101010000100000100",
			113 => "0000001000000111011101",
			114 => "0010110011001000000100",
			115 => "1111111000000111011101",
			116 => "0000001001111100000100",
			117 => "0000001000000111011101",
			118 => "1111111000000111011101",
			119 => "0000101010000100000100",
			120 => "0000001000000111111001",
			121 => "0010110011000000000100",
			122 => "1111111000000111111001",
			123 => "0000001001111100000100",
			124 => "0000000000000111111001",
			125 => "0000000000000111111001",
			126 => "0000101010000100000100",
			127 => "0000000000001000010101",
			128 => "0010110011001000000100",
			129 => "1111111000001000010101",
			130 => "0000001001111100000100",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0000101010000100000100",
			134 => "0000000000001000110001",
			135 => "0010110011001000000100",
			136 => "1111111000001000110001",
			137 => "0000001001111100000100",
			138 => "0000000000001000110001",
			139 => "0000000000001000110001",
			140 => "0000101010000100000100",
			141 => "0000000000001001001101",
			142 => "0010110011001000000100",
			143 => "0000000000001001001101",
			144 => "0000001001111100000100",
			145 => "0000000000001001001101",
			146 => "0000000000001001001101",
			147 => "0000001000000100000100",
			148 => "0000000000001001101001",
			149 => "0010011100101100000100",
			150 => "0000000000001001101001",
			151 => "0011000110101100000100",
			152 => "0000000000001001101001",
			153 => "0000000000001001101001",
			154 => "0000101010000100000100",
			155 => "0000000000001010000101",
			156 => "0010110011000000000100",
			157 => "0000000000001010000101",
			158 => "0000001001111100000100",
			159 => "0000000000001010000101",
			160 => "0000000000001010000101",
			161 => "0000101010000100000100",
			162 => "0000000000001010100001",
			163 => "0010110011000000000100",
			164 => "0000000000001010100001",
			165 => "0000001001111100000100",
			166 => "0000000000001010100001",
			167 => "0000000000001010100001",
			168 => "0000101010000100000100",
			169 => "0000000000001010111101",
			170 => "0010110011000000000100",
			171 => "0000000000001010111101",
			172 => "0000001001111100000100",
			173 => "0000000000001010111101",
			174 => "0000000000001010111101",
			175 => "0000101010000100000100",
			176 => "0000000000001011011001",
			177 => "0010010001010000000100",
			178 => "0000000000001011011001",
			179 => "0010000110101100000100",
			180 => "0000000000001011011001",
			181 => "0000000000001011011001",
			182 => "0000001000000100001000",
			183 => "0010110101010100000100",
			184 => "0000001000001011111101",
			185 => "0000001000001011111101",
			186 => "0010011100101100000100",
			187 => "1111111000001011111101",
			188 => "0010101000100000000100",
			189 => "0000000000001011111101",
			190 => "1111111000001011111101",
			191 => "0000001000000100001000",
			192 => "0010000101011100000100",
			193 => "0000000000001100100001",
			194 => "0000001000001100100001",
			195 => "0010010110011100000100",
			196 => "1111111000001100100001",
			197 => "0010010001001000000100",
			198 => "0000000000001100100001",
			199 => "1111111000001100100001",
			200 => "0000001000000100001000",
			201 => "0000101010000100000100",
			202 => "0000001000001101000101",
			203 => "0000000000001101000101",
			204 => "0010011100101100000100",
			205 => "1111111000001101000101",
			206 => "0011000110101100000100",
			207 => "0000000000001101000101",
			208 => "1111111000001101000101",
			209 => "0000101010000100000100",
			210 => "0000001000001101101001",
			211 => "0010110011001000001000",
			212 => "0011010011000000000100",
			213 => "1111111000001101101001",
			214 => "0000000000001101101001",
			215 => "0000001001111100000100",
			216 => "0000000000001101101001",
			217 => "0000000000001101101001",
			218 => "0000101010000100000100",
			219 => "0000001000001110010101",
			220 => "0010110011001000001100",
			221 => "0010110011000000000100",
			222 => "1111111000001110010101",
			223 => "0010110101111000000100",
			224 => "0000000000001110010101",
			225 => "0000000000001110010101",
			226 => "0000001001111100000100",
			227 => "0000001000001110010101",
			228 => "0000000000001110010101",
			229 => "0000101010000100000100",
			230 => "0000001000001111000001",
			231 => "0010110011001000001100",
			232 => "0010110011000000000100",
			233 => "1111111000001111000001",
			234 => "0010110101111000000100",
			235 => "0000000000001111000001",
			236 => "0000000000001111000001",
			237 => "0000001001111100000100",
			238 => "0000000000001111000001",
			239 => "0000000000001111000001",
			240 => "0000101010000100000100",
			241 => "0000001000001111110111",
			242 => "0010110011001000010000",
			243 => "0010110011000000000100",
			244 => "1111111000001111110111",
			245 => "0010110101111000001000",
			246 => "0011010011000000000100",
			247 => "0000000000001111110111",
			248 => "0000000000001111110111",
			249 => "0000000000001111110111",
			250 => "0000001001111100000100",
			251 => "0000000000001111110111",
			252 => "0000000000001111110111",
			253 => "0000001000111000000100",
			254 => "0000000000010000000001",
			255 => "1111111000010000000001",
			256 => "0000001000111000001000",
			257 => "0001111000000000000100",
			258 => "0000010000010000010101",
			259 => "0000011000010000010101",
			260 => "1111111000010000010101",
			261 => "0000001000000100000100",
			262 => "0000001000010000101001",
			263 => "0000001101001000000100",
			264 => "0000000000010000101001",
			265 => "1111111000010000101001",
			266 => "0000001000111000001000",
			267 => "0010000101011100000100",
			268 => "0000000000010000111101",
			269 => "0000001000010000111101",
			270 => "1111111000010000111101",
			271 => "0000001000111000001000",
			272 => "0001010001100100000100",
			273 => "0000000000010001010001",
			274 => "0000001000010001010001",
			275 => "1111111000010001010001",
			276 => "0000001000111000001000",
			277 => "0010000101011100000100",
			278 => "0000000000010001100101",
			279 => "0000001000010001100101",
			280 => "1111111000010001100101",
			281 => "0000001000111000001000",
			282 => "0010000101011100000100",
			283 => "0000000000010001111001",
			284 => "0000001000010001111001",
			285 => "1111111000010001111001",
			286 => "0000001000111000001000",
			287 => "0010000101011100000100",
			288 => "0000000000010010001101",
			289 => "0000000000010010001101",
			290 => "1111111000010010001101",
			291 => "0000101000000100001000",
			292 => "0000111001100000000100",
			293 => "0000000000010010100001",
			294 => "0000000000010010100001",
			295 => "0000000000010010100001",
			296 => "0000001000111000001000",
			297 => "0010000101011100000100",
			298 => "0000000000010010110101",
			299 => "0000000000010010110101",
			300 => "0000000000010010110101",
			301 => "0000001000111000001000",
			302 => "0010110101010100000100",
			303 => "0000000000010011001001",
			304 => "0000000000010011001001",
			305 => "0000000000010011001001",
			306 => "0000001000111000001000",
			307 => "0010101000011000000100",
			308 => "0000000000010011011101",
			309 => "0000000000010011011101",
			310 => "0000000000010011011101",
			311 => "0000001000111000001000",
			312 => "0010101000011000000100",
			313 => "0000000000010011110001",
			314 => "0000000000010011110001",
			315 => "0000000000010011110001",
			316 => "0000001000111000001000",
			317 => "0010000101011100000100",
			318 => "0000000000010100000101",
			319 => "0000000000010100000101",
			320 => "0000000000010100000101",
			321 => "0000001000111000001000",
			322 => "0010110101010100000100",
			323 => "0000000000010100011001",
			324 => "0000000000010100011001",
			325 => "0000000000010100011001",
			326 => "0000001000111000001000",
			327 => "0010000101011100000100",
			328 => "0000000000010100101101",
			329 => "0000000000010100101101",
			330 => "0000000000010100101101",
			331 => "0000001000111000001000",
			332 => "0010101000011000000100",
			333 => "0000000000010101000001",
			334 => "0000000000010101000001",
			335 => "0000000000010101000001",
			336 => "0000001000111000001000",
			337 => "0010000101011100000100",
			338 => "0000000000010101010101",
			339 => "0000000000010101010101",
			340 => "0000000000010101010101",
			341 => "0000101000000100001000",
			342 => "0001010001100100000100",
			343 => "0000001000010101110001",
			344 => "0000001000010101110001",
			345 => "0000001000101000000100",
			346 => "1111111000010101110001",
			347 => "1111111000010101110001",
			348 => "0000001000000100001000",
			349 => "0000101010000100000100",
			350 => "0000001000010110001101",
			351 => "0000001000010110001101",
			352 => "0000100110101100000100",
			353 => "0000000000010110001101",
			354 => "1111111000010110001101",
			355 => "0000001000000100000100",
			356 => "0000001000010110101001",
			357 => "0010011100101100000100",
			358 => "1111111000010110101001",
			359 => "0010111000111000000100",
			360 => "0000000000010110101001",
			361 => "1111111000010110101001",
			362 => "0000101010000100000100",
			363 => "0000001000010111000101",
			364 => "0010110011001000000100",
			365 => "1111111000010111000101",
			366 => "0000001001111100000100",
			367 => "0000001000010111000101",
			368 => "1111111000010111000101",
			369 => "0000101010000100000100",
			370 => "0000001000010111100001",
			371 => "0010110011001000000100",
			372 => "1111111000010111100001",
			373 => "0000001001111100000100",
			374 => "0000001000010111100001",
			375 => "1111111000010111100001",
			376 => "0000101010000100000100",
			377 => "0000000000010111111101",
			378 => "0010110011000000000100",
			379 => "1111111000010111111101",
			380 => "0000001001111100000100",
			381 => "0000000000010111111101",
			382 => "0000000000010111111101",
			383 => "0000101010000100000100",
			384 => "0000000000011000011001",
			385 => "0010110011000000000100",
			386 => "1111111000011000011001",
			387 => "0000001001111100000100",
			388 => "0000000000011000011001",
			389 => "0000000000011000011001",
			390 => "0000101010000100000100",
			391 => "0000000000011000110101",
			392 => "0010110011001000000100",
			393 => "1111111000011000110101",
			394 => "0000001001111100000100",
			395 => "0000000000011000110101",
			396 => "0000000000011000110101",
			397 => "0000101010000100000100",
			398 => "0000000000011001010001",
			399 => "0010110011001000000100",
			400 => "0000000000011001010001",
			401 => "0000001001111100000100",
			402 => "0000000000011001010001",
			403 => "0000000000011001010001",
			404 => "0000101010000100000100",
			405 => "0000000000011001101101",
			406 => "0010110011000000000100",
			407 => "0000000000011001101101",
			408 => "0000001001111100000100",
			409 => "0000000000011001101101",
			410 => "0000000000011001101101",
			411 => "0000101010000100000100",
			412 => "0000000000011010001001",
			413 => "0010110011000000000100",
			414 => "0000000000011010001001",
			415 => "0000001001111100000100",
			416 => "0000000000011010001001",
			417 => "0000000000011010001001",
			418 => "0000101010000100000100",
			419 => "0000000000011010100101",
			420 => "0010110011000000000100",
			421 => "0000000000011010100101",
			422 => "0000001001111100000100",
			423 => "0000000000011010100101",
			424 => "0000000000011010100101",
			425 => "0000101010000100000100",
			426 => "0000000000011011000001",
			427 => "0010110011000000000100",
			428 => "0000000000011011000001",
			429 => "0000001001111100000100",
			430 => "0000000000011011000001",
			431 => "0000000000011011000001",
			432 => "0000101010000100000100",
			433 => "0000000000011011011101",
			434 => "0010110011001000000100",
			435 => "0000000000011011011101",
			436 => "0010001100110000000100",
			437 => "0000000000011011011101",
			438 => "0000000000011011011101",
			439 => "0000001000000100001000",
			440 => "0000111001100000000100",
			441 => "0000001000011100000001",
			442 => "0000001000011100000001",
			443 => "0010011100101100000100",
			444 => "1111111000011100000001",
			445 => "0000111011111000000100",
			446 => "0000000000011100000001",
			447 => "1111111000011100000001",
			448 => "0000001000000100001000",
			449 => "0000101010000100000100",
			450 => "0000001000011100100101",
			451 => "0000000000011100100101",
			452 => "0010011100101100000100",
			453 => "1111111000011100100101",
			454 => "0000010011010000000100",
			455 => "0000000000011100100101",
			456 => "1111111000011100100101",
			457 => "0000001000000100001000",
			458 => "0000101010000100000100",
			459 => "0000001000011101001001",
			460 => "0000000000011101001001",
			461 => "0010011100101100000100",
			462 => "1111111000011101001001",
			463 => "0001111010011100000100",
			464 => "0000000000011101001001",
			465 => "1111111000011101001001",
			466 => "0000101010000100000100",
			467 => "0000001000011101110101",
			468 => "0010110011001000001100",
			469 => "0010110011000000000100",
			470 => "1111111000011101110101",
			471 => "0010110101111000000100",
			472 => "0000000000011101110101",
			473 => "0000000000011101110101",
			474 => "0000001001111100000100",
			475 => "0000001000011101110101",
			476 => "1111111000011101110101",
			477 => "0000101010000100000100",
			478 => "0000001000011110100001",
			479 => "0010110011001000001100",
			480 => "0010110011000000000100",
			481 => "1111111000011110100001",
			482 => "0010110101111000000100",
			483 => "0000000000011110100001",
			484 => "0000000000011110100001",
			485 => "0000001001111100000100",
			486 => "0000001000011110100001",
			487 => "0000000000011110100001",
			488 => "0000101010000100000100",
			489 => "0000001000011111001111",
			490 => "0010110011001000001100",
			491 => "0010110011000000000100",
			492 => "1111111000011111001111",
			493 => "0010110101111000000100",
			494 => "0000000000011111001111",
			495 => "0000000000011111001111",
			496 => "0000001001111100000100",
			497 => "0000000000011111001111",
			498 => "0000000000011111001111",
			499 => "0000001000111000000100",
			500 => "0000000000011111011001",
			501 => "0000000000011111011001",
			502 => "0000001000000100000100",
			503 => "0000010000011111101101",
			504 => "0000001101001000000100",
			505 => "0000000000011111101101",
			506 => "1111111000011111101101",
			507 => "0000001000111000001000",
			508 => "0010000101011100000100",
			509 => "0000000000100000000001",
			510 => "0000001000100000000001",
			511 => "1111111000100000000001",
			512 => "0000001000111000001000",
			513 => "0010000101011100000100",
			514 => "0000000000100000010101",
			515 => "0000001000100000010101",
			516 => "1111111000100000010101",
			517 => "0000001000111000001000",
			518 => "0010000101011100000100",
			519 => "0000000000100000101001",
			520 => "0000001000100000101001",
			521 => "1111111000100000101001",
			522 => "0000001000111000001000",
			523 => "0010000101011100000100",
			524 => "0000000000100000111101",
			525 => "0000001000100000111101",
			526 => "1111111000100000111101",
			527 => "0000001000111000001000",
			528 => "0011011011101100000100",
			529 => "0000000000100001010001",
			530 => "0000001000100001010001",
			531 => "1111111000100001010001",
			532 => "0000001000111000001000",
			533 => "0010000101011100000100",
			534 => "0000000000100001100101",
			535 => "0000000000100001100101",
			536 => "0000000000100001100101",
			537 => "0000001000111000001000",
			538 => "0010000101011100000100",
			539 => "0000000000100001111001",
			540 => "0000000000100001111001",
			541 => "0000000000100001111001",
			542 => "0000001000111000001000",
			543 => "0010110101010100000100",
			544 => "0000000000100010001101",
			545 => "0000000000100010001101",
			546 => "0000000000100010001101",
			547 => "0000001000111000001000",
			548 => "0010101000011000000100",
			549 => "0000000000100010100001",
			550 => "0000000000100010100001",
			551 => "0000000000100010100001",
			552 => "0000001000111000001000",
			553 => "0010110101010100000100",
			554 => "0000000000100010110101",
			555 => "0000000000100010110101",
			556 => "0000000000100010110101",
			557 => "0000001000111000001000",
			558 => "0010101000011000000100",
			559 => "0000000000100011001001",
			560 => "0000000000100011001001",
			561 => "0000000000100011001001",
			562 => "0000001000111000001000",
			563 => "0010000101011100000100",
			564 => "0000000000100011011101",
			565 => "0000000000100011011101",
			566 => "0000000000100011011101",
			567 => "0000001000111000001000",
			568 => "0010110101010100000100",
			569 => "0000000000100011110001",
			570 => "0000000000100011110001",
			571 => "0000000000100011110001",
			572 => "0000001000111000001000",
			573 => "0010101000011000000100",
			574 => "0000000000100100000101",
			575 => "0000000000100100000101",
			576 => "0000000000100100000101",
			577 => "0000001000111000001000",
			578 => "0010101000011000000100",
			579 => "0000000000100100011001",
			580 => "0000000000100100011001",
			581 => "0000000000100100011001",
			582 => "0000001000111000001000",
			583 => "0010000101011100000100",
			584 => "0000000000100100101101",
			585 => "0000000000100100101101",
			586 => "0000000000100100101101",
			587 => "0000101000000100001000",
			588 => "0010000101011100000100",
			589 => "0000001000100101001001",
			590 => "0000001000100101001001",
			591 => "0000001000101000000100",
			592 => "1111111000100101001001",
			593 => "1111111000100101001001",
			594 => "0000001000000100001000",
			595 => "0000101010000100000100",
			596 => "0000001000100101100101",
			597 => "0000001000100101100101",
			598 => "0000100110101100000100",
			599 => "0000000000100101100101",
			600 => "1111111000100101100101",
			601 => "0000101010000100000100",
			602 => "0000001000100110000001",
			603 => "0010110011001000000100",
			604 => "1111111000100110000001",
			605 => "0000001001111100000100",
			606 => "0000001000100110000001",
			607 => "1111111000100110000001",
			608 => "0000101010000100000100",
			609 => "0000001000100110011101",
			610 => "0010110011001000000100",
			611 => "1111111000100110011101",
			612 => "0000001001111100000100",
			613 => "0000001000100110011101",
			614 => "1111111000100110011101",
			615 => "0000101010000100000100",
			616 => "0000001000100110111001",
			617 => "0010110011001000000100",
			618 => "1111111000100110111001",
			619 => "0000001001111100000100",
			620 => "0000001000100110111001",
			621 => "1111111000100110111001",
			622 => "0000101010000100000100",
			623 => "0000000000100111010101",
			624 => "0010010001010000000100",
			625 => "1111111000100111010101",
			626 => "0000001010011000000100",
			627 => "0000000000100111010101",
			628 => "0000000000100111010101",
			629 => "0000101010000100000100",
			630 => "0000000000100111110001",
			631 => "0010110011000000000100",
			632 => "1111111000100111110001",
			633 => "0000001001111100000100",
			634 => "0000000000100111110001",
			635 => "0000000000100111110001",
			636 => "0000101010000100000100",
			637 => "0000000000101000001101",
			638 => "0010110011001000000100",
			639 => "1111111000101000001101",
			640 => "0000001001111100000100",
			641 => "0000000000101000001101",
			642 => "0000000000101000001101",
			643 => "0000101010000100000100",
			644 => "0000000000101000101001",
			645 => "0010110011001000000100",
			646 => "0000000000101000101001",
			647 => "0000001001111100000100",
			648 => "0000000000101000101001",
			649 => "0000000000101000101001",
			650 => "0000101010000100000100",
			651 => "0000000000101001000101",
			652 => "0010110011000000000100",
			653 => "0000000000101001000101",
			654 => "0000001001111100000100",
			655 => "0000000000101001000101",
			656 => "0000000000101001000101",
			657 => "0000101010000100000100",
			658 => "0000000000101001100001",
			659 => "0010110011000000000100",
			660 => "0000000000101001100001",
			661 => "0000001001111100000100",
			662 => "0000000000101001100001",
			663 => "0000000000101001100001",
			664 => "0000101010000100000100",
			665 => "0000000000101001111101",
			666 => "0010110011000000000100",
			667 => "0000000000101001111101",
			668 => "0000001001111100000100",
			669 => "0000000000101001111101",
			670 => "0000000000101001111101",
			671 => "0000101010000100000100",
			672 => "0000000000101010011001",
			673 => "0010010001010000000100",
			674 => "0000000000101010011001",
			675 => "0010000110101100000100",
			676 => "0000000000101010011001",
			677 => "0000000000101010011001",
			678 => "0000101010000100000100",
			679 => "0000000000101010110101",
			680 => "0010110011001000000100",
			681 => "0000000000101010110101",
			682 => "0010001100110000000100",
			683 => "0000000000101010110101",
			684 => "0000000000101010110101",
			685 => "0000001000000100001000",
			686 => "0010000101011100000100",
			687 => "0000001000101011011001",
			688 => "0000001000101011011001",
			689 => "0010010110011100000100",
			690 => "1111111000101011011001",
			691 => "0010010001001000000100",
			692 => "0000000000101011011001",
			693 => "1111111000101011011001",
			694 => "0000001000000100001000",
			695 => "0010101000011000000100",
			696 => "0000000000101011111101",
			697 => "0000001000101011111101",
			698 => "0010011100101100000100",
			699 => "1111111000101011111101",
			700 => "0000010011010000000100",
			701 => "0000000000101011111101",
			702 => "1111111000101011111101",
			703 => "0000001000000100001000",
			704 => "0010101000011000000100",
			705 => "0000000000101100100001",
			706 => "0000000000101100100001",
			707 => "0010011100101100000100",
			708 => "0000000000101100100001",
			709 => "0011000110101100000100",
			710 => "0000000000101100100001",
			711 => "0000000000101100100001",
			712 => "0000101010000100000100",
			713 => "0000001000101101001101",
			714 => "0010110011001000001100",
			715 => "0010110011000000000100",
			716 => "1111111000101101001101",
			717 => "0010110101111000000100",
			718 => "0000000000101101001101",
			719 => "0000000000101101001101",
			720 => "0000001001111100000100",
			721 => "0000001000101101001101",
			722 => "1111111000101101001101",
			723 => "0000101010000100000100",
			724 => "0000001000101101111001",
			725 => "0010110011001000001100",
			726 => "0010110011000000000100",
			727 => "1111111000101101111001",
			728 => "0010110101111000000100",
			729 => "0000000000101101111001",
			730 => "0000000000101101111001",
			731 => "0000001001111100000100",
			732 => "0000000000101101111001",
			733 => "0000000000101101111001",
			734 => "0000101010000100000100",
			735 => "0000000000101110100111",
			736 => "0010110011001000001100",
			737 => "0011010011000000000100",
			738 => "1111111000101110100111",
			739 => "0011010101111000000100",
			740 => "0000000000101110100111",
			741 => "0000000000101110100111",
			742 => "0000001001111100000100",
			743 => "0000000000101110100111",
			744 => "0000000000101110100111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(253, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(499, initial_addr_3'length));
	end generate gen_rom_12;

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
