-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom_centroids is
    generic(ADDRESS_BITS: positive := 8;
            DATA_LENGTH:  positive := 13);
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0));

end rom_centroids;

architecture Behavioral of rom_centroids is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin
	bank <= (
		0 => "1000100000011",
		1 => "1000110001011",
		2 => "0000111101001",
		3 => "0010110000100",
		4 => "0100110110001",
		215 => "0000011011100",
		5 => "0110001000101",
		6 => "0000000110101",
		7 => "0011010111000",
		8 => "0110110101000",
		9 => "1100011111011",
		10 => "0010010101111",
		171 => "0001110010111",
		198 => "0000101001101",
		12 => "0010001010010",
		13 => "0011101111000",
		14 => "0010000111101",
		15 => "0000011110001",
		16 => "0100000000010",
		17 => "0000100000110",
		117 => "0100110000111",
		18 => "0011101100110",
		20 => "0001010010110",
		21 => "0001011101000",
		22 => "0011011000101",
		23 => "0101000111010",
		234 => "0011111011010",
		24 => "1101000000001",
		25 => "0111000100100",
		26 => "0011001010111",
		27 => "0110101101110",
		28 => "0001011110111",
		29 => "0001101111011",
		30 => "0000100101100",
		31 => "0010110100111",
		32 => "0100011001000",
		33 => "0100100001011",
		34 => "0011011111111",
		35 => "0000001110010",
		36 => "0111001100011",
		131 => "0100110011101",
		38 => "0001111110111",
		39 => "0100000111100",
		41 => "0110011000001",
		42 => "0001110001010",
		43 => "0001000011100",
		44 => "0101101110111",
		45 => "0011110100101",
		89 => "0011011001111",
		47 => "0010000000110",
		49 => "1011101110100",
		50 => "0100010011010",
		51 => "0101110011101",
		52 => "0010000101010",
		53 => "0110010000001",
		54 => "0110101010101",
		70 => "0010111110111",
		56 => "0011000000100",
		57 => "1101001100110",
		58 => "0001000110000",
		134 => "0011001101101",
		225 => "0100000001101",
		62 => "0111111000110",
		63 => "0010000011001",
		141 => "0101011101101",
		64 => "0010011010010",
		65 => "0011010101010",
		66 => "0010110011101",
		67 => "0110001100100",
		68 => "0011100001110",
		69 => "0010010010010",
		55 => "0010100001111",
		71 => "1010101101101",
		74 => "0100001011100",
		244 => "0100000100011",
		75 => "0000111001000",
		77 => "0000101000011",
		79 => "0000110000111",
		80 => "0101100100001",
		81 => "0001011011001",
		82 => "0100000010110",
		83 => "1000101100011",
		84 => "0000110100010",
		200 => "0000000100100",
		76 => "1001010110010",
		86 => "1001011011110",
		87 => "0000011111011",
		249 => "0100111011011",
		88 => "1000100101010",
		46 => "0101110101110",
		139 => "0001110110000",
		248 => "0110010010111",
		184 => "0110011110110",
		92 => "0100001001101",
		95 => "1100110000101",
		96 => "0000001000100",
		97 => "0010101000110",
		98 => "0001101001000",
		99 => "0101101001100",
		100 => "0100011011101",
		40 => "1010111110011",
		104 => "0011110111000",
		105 => "0011001000100",
		106 => "0000010010001",
		107 => "0100111001010",
		108 => "0111010101010",
		109 => "0011011101110",
		110 => "0101010011100",
		111 => "0100101010010",
		143 => "0010011100101",
		113 => "0001101101001",
		114 => "0010111010000",
		115 => "1100000011101",
		116 => "0011010011111",
		252 => "1010000101011",
		118 => "0100101000010",
		119 => "0110100101110",
		73 => "1001111101000",
		121 => "0000010100000",
		103 => "0001011001010",
		123 => "0000111011001",
		124 => "0011100111011",
		125 => "0001001000100",
		126 => "0010001111010",
		127 => "0100001101010",
		102 => "0001010001010",
		191 => "0000100001111",
		128 => "0011000010111",
		129 => "0101011011101",
		130 => "0101110001100",
		37 => "0101010000010",
		132 => "0000110010010",
		133 => "0001001100111",
		60 => "0101101100001",
		135 => "0101100000001",
		136 => "0100111101110",
		137 => "0001001010111",
		138 => "0101001001010",
		90 => "1101000110001",
		140 => "0001111000011",
		72 => "1001100110101",
		142 => "0010011110000",
		112 => "0001110100010",
		237 => "0100011111100",
		221 => "0110110001000",
		145 => "0001001111000",
		146 => "0011000101010",
		147 => "0110000001101",
		148 => "0100000101111",
		149 => "0011101010110",
		255 => "1010110101111",
		150 => "0000011100111",
		151 => "0100001110100",
		152 => "0100011101101",
		153 => "0000101110110",
		154 => "0001100100011",
		155 => "1001001010000",
		157 => "0011000110110",
		48 => "0101001011101",
		159 => "0000110110111",
		160 => "0010001011111",
		172 => "0001010101001",
		161 => "0100101110110",
		162 => "0100001111110",
		163 => "0011010010010",
		164 => "1001000001111",
		165 => "0011101001001",
		167 => "0011001111001",
		168 => "0000111111001",
		169 => "0001000001010",
		170 => "1000011100010",
		11 => "0110111110101",
		19 => "0111100000010",
		173 => "0101111100000",
		174 => "0010111011011",
		175 => "0010110110110",
		176 => "0011000010000",
		177 => "0010010100010",
		178 => "0110101000010",
		179 => "0000101101100",
		181 => "0001100111000",
		182 => "1000111100111",
		189 => "0011100101111",
		91 => "0010100110011",
		185 => "0111101101111",
		186 => "0000011000000",
		187 => "0101000000001",
		188 => "0101010110011",
		93 => "0011100011101",
		190 => "0100111000001",
		158 => "0000001111111",
		192 => "0100100110000",
		193 => "0001100001001",
		194 => "0010010111110",
		245 => "0100101100011",
		195 => "0101100110011",
		156 => "0010100000100",
		197 => "0100010110010",
		94 => "1100010010000",
		199 => "0001010111001",
		183 => "0011011011111",
		201 => "0011111100111",
		202 => "0010110001111",
		203 => "0010101010100",
		204 => "0010100101001",
		206 => "0101000011000",
		207 => "0110111001010",
		208 => "1000000001000",
		211 => "1011010110110",
		212 => "0001111011000",
		213 => "0010110111110",
		214 => "0000101100001",
		180 => "1100111000001",
		216 => "0010100011011",
		217 => "1010100010000",
		218 => "0000010110000",
		247 => "0011010000110",
		219 => "0101000101011",
		59 => "0110011010110",
		222 => "0010101110100",
		223 => "0000100111010",
		61 => "0110010101110",
		205 => "0000001100010",
		226 => "1000110110011",
		120 => "0011111110101",
		228 => "0100010001011",
		229 => "0000100010111",
		230 => "1000001101100",
		231 => "0000000010111",
		232 => "0000001010001",
		233 => "0101100010010",
		209 => "0011111001010",
		235 => "0011110001111",
		236 => "0010111101001",
		224 => "0101011000111",
		144 => "0110100010111",
		238 => "0110000101000",
		239 => "0010001101100",
		240 => "0000101111101",
		241 => "0001111100110",
		122 => "0000100100000",
		242 => "0001101011000",
		85 => "0101111110100",
		243 => "0000011001110",
		210 => "0101111000101",
		78 => "1000010111011",
		246 => "1001110000111",
		196 => "0100100011101",
		227 => "0010101100011",
		166 => "0000101010111",
		250 => "0101001101100",
		251 => "1001010010101",
		220 => "1011111000011",
		253 => "1010010011010",
		254 => "1100100111110",
		101 => "1010001011101",
		others => (others => '0')
	);

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
