-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive;
            DATA_LENGTH:  positive;
            SELECT_ROM:  integer := 0); -- Select which ROM to use
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0);
         initial_addr_2: out std_logic_vector (ADDRESS_BITS - 1 downto 0);
         initial_addr_3: out std_logic_vector (ADDRESS_BITS - 1 downto 0));
end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin

	gen_rom_0: if SELECT_ROM = 0 generate
		bank <= (
			0 => x"0d00170c",
			1 => x"08001f04",
			2 => x"fe63005d",
			3 => x"05002204",
			4 => x"0130005d",
			5 => x"fe74005d",
			6 => x"0f006504",
			7 => x"fe6a005d",
			8 => x"0500561c",
			9 => x"07003f10",
			10 => x"0000d304",
			11 => x"023b005d",
			12 => x"09002004",
			13 => x"fe35005d",
			14 => x"02013704",
			15 => x"009e005d",
			16 => x"ff0d005d",
			17 => x"05003508",
			18 => x"0a003104",
			19 => x"01ae005d",
			20 => x"002d005d",
			21 => x"01b8005d",
			22 => x"fe5d005d",
			23 => x"0d001710",
			24 => x"05002208",
			25 => x"0a002704",
			26 => x"fff300e9",
			27 => x"001f00e9",
			28 => x"09002304",
			29 => x"ff9900e9",
			30 => x"000300e9",
			31 => x"04002b1c",
			32 => x"0f006504",
			33 => x"ffcf00e9",
			34 => x"00014610",
			35 => x"09001e04",
			36 => x"ffec00e9",
			37 => x"0a003104",
			38 => x"008e00e9",
			39 => x"08002304",
			40 => x"ffda00e9",
			41 => x"004c00e9",
			42 => x"0d001f04",
			43 => x"ffa900e9",
			44 => x"004800e9",
			45 => x"04002e0c",
			46 => x"01001908",
			47 => x"00012904",
			48 => x"fffe00e9",
			49 => x"ff9a00e9",
			50 => x"001000e9",
			51 => x"03004008",
			52 => x"00010404",
			53 => x"fff500e9",
			54 => x"006e00e9",
			55 => x"01001704",
			56 => x"ffc600e9",
			57 => x"000100e9",
			58 => x"01001220",
			59 => x"08002210",
			60 => x"01000e04",
			61 => x"fe480175",
			62 => x"0b001508",
			63 => x"0d001504",
			64 => x"fe4d0175",
			65 => x"00ad0175",
			66 => x"fe450175",
			67 => x"0c001b08",
			68 => x"09002004",
			69 => x"ffd70175",
			70 => x"03480175",
			71 => x"0c001d04",
			72 => x"fff30175",
			73 => x"fe480175",
			74 => x"0f008208",
			75 => x"09002404",
			76 => x"005f0175",
			77 => x"fe490175",
			78 => x"0300411c",
			79 => x"0d001904",
			80 => x"ffc10175",
			81 => x"05003910",
			82 => x"07004008",
			83 => x"02013704",
			84 => x"02250175",
			85 => x"fecc0175",
			86 => x"04002704",
			87 => x"02d20175",
			88 => x"02580175",
			89 => x"0c001c04",
			90 => x"02430175",
			91 => x"02ad0175",
			92 => x"fecd0175",
			93 => x"01001438",
			94 => x"01001224",
			95 => x"01000e08",
			96 => x"08002304",
			97 => x"fe3e0219",
			98 => x"fed10219",
			99 => x"0f008c0c",
			100 => x"0c001908",
			101 => x"07002404",
			102 => x"fe460219",
			103 => x"003c0219",
			104 => x"fe3e0219",
			105 => x"08002208",
			106 => x"0a002d04",
			107 => x"00750219",
			108 => x"fe350219",
			109 => x"0f00c204",
			110 => x"03060219",
			111 => x"fffe0219",
			112 => x"0f008208",
			113 => x"06006504",
			114 => x"fe410219",
			115 => x"ff530219",
			116 => x"00011f04",
			117 => x"03c20219",
			118 => x"05003804",
			119 => x"fe2b0219",
			120 => x"029e0219",
			121 => x"0f009308",
			122 => x"0c002404",
			123 => x"ff400219",
			124 => x"fe400219",
			125 => x"09002404",
			126 => x"00ea0219",
			127 => x"08002604",
			128 => x"02b90219",
			129 => x"0d001c04",
			130 => x"04070219",
			131 => x"04002104",
			132 => x"02a80219",
			133 => x"03700219",
			134 => x"0d001914",
			135 => x"05002208",
			136 => x"0a002704",
			137 => x"ffe802cd",
			138 => x"002b02cd",
			139 => x"0e00a508",
			140 => x"0a002704",
			141 => x"fffc02cd",
			142 => x"ff8302cd",
			143 => x"000602cd",
			144 => x"0c001e1c",
			145 => x"0e008d10",
			146 => x"06009908",
			147 => x"06005e04",
			148 => x"ffea02cd",
			149 => x"009a02cd",
			150 => x"0f00b904",
			151 => x"ff9702cd",
			152 => x"ffe402cd",
			153 => x"02013904",
			154 => x"00a602cd",
			155 => x"0e009c04",
			156 => x"ffab02cd",
			157 => x"001f02cd",
			158 => x"01001718",
			159 => x"0500380c",
			160 => x"05003308",
			161 => x"01001404",
			162 => x"ffde02cd",
			163 => x"002902cd",
			164 => x"ff3c02cd",
			165 => x"05005308",
			166 => x"0f00ba04",
			167 => x"000102cd",
			168 => x"004f02cd",
			169 => x"ffc702cd",
			170 => x"0e00950c",
			171 => x"00013108",
			172 => x"06008a04",
			173 => x"ffee02cd",
			174 => x"003e02cd",
			175 => x"ffc202cd",
			176 => x"0b001f04",
			177 => x"fffa02cd",
			178 => x"009402cd",
			179 => x"01001434",
			180 => x"01001224",
			181 => x"01001018",
			182 => x"08002310",
			183 => x"01000e04",
			184 => x"df540379",
			185 => x"0f008c04",
			186 => x"df550379",
			187 => x"0600a804",
			188 => x"e1b90379",
			189 => x"df5a0379",
			190 => x"09002604",
			191 => x"e1b90379",
			192 => x"df570379",
			193 => x"0f008204",
			194 => x"df550379",
			195 => x"00012e04",
			196 => x"e4180379",
			197 => x"e0320379",
			198 => x"0f008208",
			199 => x"09002604",
			200 => x"e0280379",
			201 => x"df560379",
			202 => x"05003804",
			203 => x"e1e30379",
			204 => x"e8990379",
			205 => x"06008508",
			206 => x"07003004",
			207 => x"e0280379",
			208 => x"df560379",
			209 => x"04002108",
			210 => x"0b001d04",
			211 => x"e3240379",
			212 => x"e9230379",
			213 => x"08002604",
			214 => x"e8420379",
			215 => x"0100170c",
			216 => x"05003804",
			217 => x"e8a20379",
			218 => x"05004204",
			219 => x"ec0d0379",
			220 => x"e98d0379",
			221 => x"ec150379",
			222 => x"01001220",
			223 => x"08002210",
			224 => x"01000e04",
			225 => x"fe5d0405",
			226 => x"0200e908",
			227 => x"06006f04",
			228 => x"fe650405",
			229 => x"01df0405",
			230 => x"fe590405",
			231 => x"0c001d0c",
			232 => x"09002004",
			233 => x"ff590405",
			234 => x"05003404",
			235 => x"00060405",
			236 => x"01fa0405",
			237 => x"fe630405",
			238 => x"06005e04",
			239 => x"fe620405",
			240 => x"03004620",
			241 => x"0d001f14",
			242 => x"0f00aa04",
			243 => x"021c0405",
			244 => x"04002108",
			245 => x"04002004",
			246 => x"006f0405",
			247 => x"fe470405",
			248 => x"07003704",
			249 => x"ff980405",
			250 => x"01840405",
			251 => x"03002e08",
			252 => x"03002d04",
			253 => x"01cf0405",
			254 => x"00190405",
			255 => x"01cf0405",
			256 => x"fe0c0405",
			257 => x"08002320",
			258 => x"0f00bb18",
			259 => x"01000e04",
			260 => x"ff5c04c1",
			261 => x"0f00820c",
			262 => x"0a002a08",
			263 => x"01001204",
			264 => x"ffe404c1",
			265 => x"003d04c1",
			266 => x"ff7404c1",
			267 => x"0f00a904",
			268 => x"009e04c1",
			269 => x"001404c1",
			270 => x"0e00a504",
			271 => x"ff1804c1",
			272 => x"000a04c1",
			273 => x"02012b24",
			274 => x"01001a18",
			275 => x"0700330c",
			276 => x"0000db08",
			277 => x"0000a204",
			278 => x"ffcb04c1",
			279 => x"009104c1",
			280 => x"ff7004c1",
			281 => x"03004608",
			282 => x"06008504",
			283 => x"ffeb04c1",
			284 => x"011404c1",
			285 => x"ffbe04c1",
			286 => x"0f00c208",
			287 => x"00010c04",
			288 => x"ffe604c1",
			289 => x"002b04c1",
			290 => x"ff7004c1",
			291 => x"01001910",
			292 => x"0c001c04",
			293 => x"004904c1",
			294 => x"05003804",
			295 => x"ff4004c1",
			296 => x"0600b704",
			297 => x"ffc404c1",
			298 => x"007d04c1",
			299 => x"01001a04",
			300 => x"00cc04c1",
			301 => x"01001c04",
			302 => x"ffcb04c1",
			303 => x"004504c1",
			304 => x"01001220",
			305 => x"08002210",
			306 => x"01000e04",
			307 => x"fe4d0555",
			308 => x"0b001708",
			309 => x"09001d04",
			310 => x"fe4c0555",
			311 => x"01640555",
			312 => x"fe4d0555",
			313 => x"0c001d0c",
			314 => x"07002c04",
			315 => x"fe4e0555",
			316 => x"0f00c204",
			317 => x"03560555",
			318 => x"001f0555",
			319 => x"fe4d0555",
			320 => x"0f008708",
			321 => x"0b001c04",
			322 => x"ff480555",
			323 => x"fe4f0555",
			324 => x"0d001904",
			325 => x"ffab0555",
			326 => x"0a00471c",
			327 => x"0500380c",
			328 => x"00011f04",
			329 => x"03020555",
			330 => x"07004004",
			331 => x"00a30555",
			332 => x"02420555",
			333 => x"07003b08",
			334 => x"0e008b04",
			335 => x"028e0555",
			336 => x"012f0555",
			337 => x"0c001e04",
			338 => x"02b90555",
			339 => x"02660555",
			340 => x"00730555",
			341 => x"08002320",
			342 => x"06009518",
			343 => x"06008010",
			344 => x"0d001804",
			345 => x"ff9d0601",
			346 => x"0a003108",
			347 => x"0a002804",
			348 => x"fff70601",
			349 => x"00380601",
			350 => x"ffe30601",
			351 => x"01000c04",
			352 => x"fff20601",
			353 => x"005f0601",
			354 => x"04002a04",
			355 => x"ff650601",
			356 => x"002a0601",
			357 => x"0a00432c",
			358 => x"05003820",
			359 => x"07004018",
			360 => x"0400200c",
			361 => x"09002504",
			362 => x"00920601",
			363 => x"0d001f04",
			364 => x"ffcb0601",
			365 => x"00190601",
			366 => x"01001404",
			367 => x"ff730601",
			368 => x"0f00c204",
			369 => x"007e0601",
			370 => x"ffc20601",
			371 => x"0d002404",
			372 => x"00780601",
			373 => x"00000601",
			374 => x"0f00b808",
			375 => x"03003304",
			376 => x"001a0601",
			377 => x"ffd50601",
			378 => x"00ad0601",
			379 => x"01001808",
			380 => x"07004104",
			381 => x"ffb70601",
			382 => x"00020601",
			383 => x"00070601",
			384 => x"05003420",
			385 => x"08002718",
			386 => x"0200ca0c",
			387 => x"0e005b04",
			388 => x"ffe006bd",
			389 => x"0d001504",
			390 => x"fff006bd",
			391 => x"004406bd",
			392 => x"0a002708",
			393 => x"07002c04",
			394 => x"fff806bd",
			395 => x"000806bd",
			396 => x"ff9f06bd",
			397 => x"0e008a04",
			398 => x"ffde06bd",
			399 => x"004706bd",
			400 => x"0a003b24",
			401 => x"02013718",
			402 => x"01000e04",
			403 => x"ffe806bd",
			404 => x"01001a0c",
			405 => x"0600b908",
			406 => x"04002d04",
			407 => x"007706bd",
			408 => x"fffc06bd",
			409 => x"fffb06bd",
			410 => x"03003104",
			411 => x"000906bd",
			412 => x"ffee06bd",
			413 => x"02014108",
			414 => x"0600bf04",
			415 => x"ffc706bd",
			416 => x"fffe06bd",
			417 => x"003306bd",
			418 => x"0600b718",
			419 => x"01001710",
			420 => x"07003308",
			421 => x"07003104",
			422 => x"ffee06bd",
			423 => x"001006bd",
			424 => x"07004004",
			425 => x"ffa906bd",
			426 => x"000006bd",
			427 => x"00012104",
			428 => x"fffe06bd",
			429 => x"000d06bd",
			430 => x"002b06bd",
			431 => x"0100121c",
			432 => x"08002314",
			433 => x"01000e04",
			434 => x"fe530759",
			435 => x"0f008204",
			436 => x"fe560759",
			437 => x"0e007c04",
			438 => x"02170759",
			439 => x"07003504",
			440 => x"fe490759",
			441 => x"00080759",
			442 => x"0c001d04",
			443 => x"01c10759",
			444 => x"fe550759",
			445 => x"0f008208",
			446 => x"09002304",
			447 => x"00910759",
			448 => x"fe560759",
			449 => x"07003f18",
			450 => x"02013714",
			451 => x"0d001904",
			452 => x"ff8a0759",
			453 => x"00011f08",
			454 => x"07003804",
			455 => x"02c80759",
			456 => x"01f80759",
			457 => x"01001404",
			458 => x"ffec0759",
			459 => x"01ab0759",
			460 => x"feb50759",
			461 => x"00011e04",
			462 => x"011c0759",
			463 => x"05003508",
			464 => x"02013404",
			465 => x"02220759",
			466 => x"01230759",
			467 => x"08002704",
			468 => x"02970759",
			469 => x"021a0759",
			470 => x"0800231c",
			471 => x"01000e04",
			472 => x"fe6107dd",
			473 => x"09001d04",
			474 => x"fe5807dd",
			475 => x"0c001a0c",
			476 => x"0a002d04",
			477 => x"017207dd",
			478 => x"07003004",
			479 => x"fe5307dd",
			480 => x"00a607dd",
			481 => x"0f009304",
			482 => x"fe6a07dd",
			483 => x"ff8b07dd",
			484 => x"0f007504",
			485 => x"fe6a07dd",
			486 => x"03004620",
			487 => x"05003810",
			488 => x"03002704",
			489 => x"01b607dd",
			490 => x"07004408",
			491 => x"02012704",
			492 => x"00be07dd",
			493 => x"ff2b07dd",
			494 => x"01aa07dd",
			495 => x"07003b08",
			496 => x"09002604",
			497 => x"004107dd",
			498 => x"01ae07dd",
			499 => x"0c001e04",
			500 => x"020e07dd",
			501 => x"01af07dd",
			502 => x"fe3a07dd",
			503 => x"0e00944c",
			504 => x"0f00c034",
			505 => x"04002218",
			506 => x"09001e0c",
			507 => x"04002004",
			508 => x"ffc708a1",
			509 => x"0000c504",
			510 => x"001c08a1",
			511 => x"fff708a1",
			512 => x"06006504",
			513 => x"ffe508a1",
			514 => x"0a003104",
			515 => x"007308a1",
			516 => x"fffe08a1",
			517 => x"08002410",
			518 => x"0f00b90c",
			519 => x"0d001b04",
			520 => x"ff8008a1",
			521 => x"0d001c04",
			522 => x"000d08a1",
			523 => x"ffff08a1",
			524 => x"000208a1",
			525 => x"03004608",
			526 => x"0e008504",
			527 => x"ffee08a1",
			528 => x"005908a1",
			529 => x"ffd808a1",
			530 => x"08002914",
			531 => x"04001d08",
			532 => x"0a002c04",
			533 => x"fff908a1",
			534 => x"000f08a1",
			535 => x"0b001808",
			536 => x"0b001704",
			537 => x"fff908a1",
			538 => x"000f08a1",
			539 => x"ff7908a1",
			540 => x"000d08a1",
			541 => x"01001710",
			542 => x"05003808",
			543 => x"0600b704",
			544 => x"001f08a1",
			545 => x"ff9908a1",
			546 => x"0600b704",
			547 => x"fffc08a1",
			548 => x"004c08a1",
			549 => x"0d001f04",
			550 => x"000108a1",
			551 => x"007608a1",
			552 => x"0d00170c",
			553 => x"09002304",
			554 => x"fe800945",
			555 => x"08001d04",
			556 => x"ff6f0945",
			557 => x"006b0945",
			558 => x"07003e38",
			559 => x"0f00c224",
			560 => x"08002618",
			561 => x"0c001908",
			562 => x"09001e04",
			563 => x"feac0945",
			564 => x"00d80945",
			565 => x"07003a08",
			566 => x"09002304",
			567 => x"fe6f0945",
			568 => x"ffa90945",
			569 => x"01001004",
			570 => x"ff6e0945",
			571 => x"018b0945",
			572 => x"09002c08",
			573 => x"00010c04",
			574 => x"006f0945",
			575 => x"01990945",
			576 => x"fec20945",
			577 => x"04002108",
			578 => x"0f00d204",
			579 => x"fdf20945",
			580 => x"ffe50945",
			581 => x"0600af04",
			582 => x"01120945",
			583 => x"08002604",
			584 => x"fe5e0945",
			585 => x"00e70945",
			586 => x"03002e08",
			587 => x"03002d04",
			588 => x"015d0945",
			589 => x"feb70945",
			590 => x"03005304",
			591 => x"01980945",
			592 => x"ff2b0945",
			593 => x"08002640",
			594 => x"02011c28",
			595 => x"0b001e24",
			596 => x"09001e0c",
			597 => x"05002208",
			598 => x"0a002704",
			599 => x"fff20a11",
			600 => x"00220a11",
			601 => x"ffb40a11",
			602 => x"0d00170c",
			603 => x"05002404",
			604 => x"00050a11",
			605 => x"09002304",
			606 => x"ffcb0a11",
			607 => x"00040a11",
			608 => x"0f006504",
			609 => x"ffe20a11",
			610 => x"04003404",
			611 => x"008b0a11",
			612 => x"ffef0a11",
			613 => x"ffbb0a11",
			614 => x"05003a10",
			615 => x"0e00a30c",
			616 => x"0a003108",
			617 => x"0a002f04",
			618 => x"ffe30a11",
			619 => x"00110a11",
			620 => x"ff570a11",
			621 => x"00110a11",
			622 => x"0600a904",
			623 => x"ffd80a11",
			624 => x"003f0a11",
			625 => x"04002110",
			626 => x"0300270c",
			627 => x"08002704",
			628 => x"fff80a11",
			629 => x"0b002504",
			630 => x"00340a11",
			631 => x"fffa0a11",
			632 => x"ffc30a11",
			633 => x"01001408",
			634 => x"0200e304",
			635 => x"00020a11",
			636 => x"ffeb0a11",
			637 => x"08002d08",
			638 => x"03004404",
			639 => x"00d20a11",
			640 => x"fffd0a11",
			641 => x"0e009504",
			642 => x"ffdb0a11",
			643 => x"00230a11",
			644 => x"08002320",
			645 => x"0f00bb18",
			646 => x"01000e04",
			647 => x"ff630add",
			648 => x"0f00820c",
			649 => x"0a002a08",
			650 => x"01001204",
			651 => x"ffe50add",
			652 => x"003d0add",
			653 => x"ff7a0add",
			654 => x"0f00a904",
			655 => x"00940add",
			656 => x"00130add",
			657 => x"0e00a504",
			658 => x"ff200add",
			659 => x"000a0add",
			660 => x"02012b30",
			661 => x"01001a24",
			662 => x"06009d18",
			663 => x"03002d08",
			664 => x"0000ae04",
			665 => x"ffdb0add",
			666 => x"009f0add",
			667 => x"01001408",
			668 => x"0000d804",
			669 => x"00050add",
			670 => x"ff5c0add",
			671 => x"05004304",
			672 => x"003c0add",
			673 => x"00010add",
			674 => x"04003308",
			675 => x"02012704",
			676 => x"01260add",
			677 => x"004a0add",
			678 => x"ffe70add",
			679 => x"0f00c208",
			680 => x"00010c04",
			681 => x"ffe70add",
			682 => x"002a0add",
			683 => x"ff770add",
			684 => x"0700400c",
			685 => x"03002e04",
			686 => x"ff5e0add",
			687 => x"03003104",
			688 => x"00cf0add",
			689 => x"ff680add",
			690 => x"0c002104",
			691 => x"00c80add",
			692 => x"0c002304",
			693 => x"ffc40add",
			694 => x"00500add",
			695 => x"01001220",
			696 => x"08002210",
			697 => x"01000e04",
			698 => x"fe5a0b79",
			699 => x"04001e04",
			700 => x"fe5b0b79",
			701 => x"03002a04",
			702 => x"011a0b79",
			703 => x"fe5d0b79",
			704 => x"0c001d0c",
			705 => x"07002c04",
			706 => x"fe680b79",
			707 => x"0f00be04",
			708 => x"01f60b79",
			709 => x"004e0b79",
			710 => x"fe5e0b79",
			711 => x"0f006504",
			712 => x"fe5c0b79",
			713 => x"0a004a28",
			714 => x"0d001f14",
			715 => x"0f00aa04",
			716 => x"025e0b79",
			717 => x"07003708",
			718 => x"0f00bf04",
			719 => x"ff690b79",
			720 => x"fe230b79",
			721 => x"03002a04",
			722 => x"ffd00b79",
			723 => x"01780b79",
			724 => x"01001708",
			725 => x"05003904",
			726 => x"00940b79",
			727 => x"01db0b79",
			728 => x"03002e08",
			729 => x"0e009d04",
			730 => x"01430b79",
			731 => x"01db0b79",
			732 => x"01e50b79",
			733 => x"fe1e0b79",
			734 => x"08002330",
			735 => x"0e008928",
			736 => x"07002f18",
			737 => x"0a002a14",
			738 => x"0400200c",
			739 => x"0c001704",
			740 => x"ff8b0c4d",
			741 => x"0c001904",
			742 => x"00310c4d",
			743 => x"ffe40c4d",
			744 => x"05002d04",
			745 => x"007d0c4d",
			746 => x"fff00c4d",
			747 => x"ff470c4d",
			748 => x"0400360c",
			749 => x"00012508",
			750 => x"01000e04",
			751 => x"fff50c4d",
			752 => x"00c40c4d",
			753 => x"ffd70c4d",
			754 => x"ffce0c4d",
			755 => x"0e00a504",
			756 => x"fef30c4d",
			757 => x"00290c4d",
			758 => x"0a003b24",
			759 => x"00014618",
			760 => x"0e008a0c",
			761 => x"0f00b008",
			762 => x"0f006504",
			763 => x"ffc00c4d",
			764 => x"00a50c4d",
			765 => x"ff980c4d",
			766 => x"0c001e04",
			767 => x"012b0c4d",
			768 => x"08002904",
			769 => x"ffa50c4d",
			770 => x"00d30c4d",
			771 => x"0d001f04",
			772 => x"ff3a0c4d",
			773 => x"04002704",
			774 => x"00ab0c4d",
			775 => x"fff00c4d",
			776 => x"0600b714",
			777 => x"0100170c",
			778 => x"00012a08",
			779 => x"00010804",
			780 => x"ffe10c4d",
			781 => x"00170c4d",
			782 => x"ff220c4d",
			783 => x"00011604",
			784 => x"fff40c4d",
			785 => x"002d0c4d",
			786 => x"00720c4d",
			787 => x"0a003b3c",
			788 => x"05003930",
			789 => x"0d002128",
			790 => x"0201371c",
			791 => x"03002f10",
			792 => x"03002a08",
			793 => x"01001604",
			794 => x"003b0cf1",
			795 => x"ff700cf1",
			796 => x"09002104",
			797 => x"ffbc0cf1",
			798 => x"00c80cf1",
			799 => x"01001708",
			800 => x"03003304",
			801 => x"ff690cf1",
			802 => x"000d0cf1",
			803 => x"00350cf1",
			804 => x"0f00dd04",
			805 => x"ff470cf1",
			806 => x"0f00e704",
			807 => x"003c0cf1",
			808 => x"ffc10cf1",
			809 => x"00011404",
			810 => x"ffe90cf1",
			811 => x"00950cf1",
			812 => x"0d001704",
			813 => x"ffdf0cf1",
			814 => x"0b002304",
			815 => x"00a70cf1",
			816 => x"00010cf1",
			817 => x"0600b714",
			818 => x"00013a10",
			819 => x"0d001b04",
			820 => x"ff980cf1",
			821 => x"04003e08",
			822 => x"00010f04",
			823 => x"fff10cf1",
			824 => x"007d0cf1",
			825 => x"ffcf0cf1",
			826 => x"ff610cf1",
			827 => x"00320cf1",
			828 => x"0d001b34",
			829 => x"0c001a24",
			830 => x"0900211c",
			831 => x"0200ca14",
			832 => x"0400210c",
			833 => x"09001d04",
			834 => x"ffe30dd5",
			835 => x"00009604",
			836 => x"fffb0dd5",
			837 => x"007b0dd5",
			838 => x"0000ca04",
			839 => x"ffba0dd5",
			840 => x"001a0dd5",
			841 => x"05003a04",
			842 => x"ff850dd5",
			843 => x"00160dd5",
			844 => x"06006b04",
			845 => x"ffee0dd5",
			846 => x"00870dd5",
			847 => x"05003a04",
			848 => x"ff5c0dd5",
			849 => x"0a003b04",
			850 => x"004c0dd5",
			851 => x"07003904",
			852 => x"ffaf0dd5",
			853 => x"00150dd5",
			854 => x"0400211c",
			855 => x"08002408",
			856 => x"07003204",
			857 => x"fff50dd5",
			858 => x"00550dd5",
			859 => x"08002a10",
			860 => x"04001a08",
			861 => x"04001804",
			862 => x"fffb0dd5",
			863 => x"001b0dd5",
			864 => x"0e008604",
			865 => x"00070dd5",
			866 => x"ff490dd5",
			867 => x"003f0dd5",
			868 => x"0a00431c",
			869 => x"0d00200c",
			870 => x"00014c08",
			871 => x"0e008004",
			872 => x"00150dd5",
			873 => x"00cd0dd5",
			874 => x"ffeb0dd5",
			875 => x"09002b08",
			876 => x"05003804",
			877 => x"ffa50dd5",
			878 => x"002a0dd5",
			879 => x"00012804",
			880 => x"00000dd5",
			881 => x"00500dd5",
			882 => x"03004504",
			883 => x"00030dd5",
			884 => x"ffb20dd5",
			885 => x"0d001708",
			886 => x"08002204",
			887 => x"fe6f0e49",
			888 => x"ff6b0e49",
			889 => x"03004530",
			890 => x"05003920",
			891 => x"0400291c",
			892 => x"0d001f10",
			893 => x"0f00ae08",
			894 => x"06005e04",
			895 => x"fea30e49",
			896 => x"01650e49",
			897 => x"07003304",
			898 => x"fe460e49",
			899 => x"ffdf0e49",
			900 => x"0e009508",
			901 => x"08002a04",
			902 => x"01100e49",
			903 => x"ff4a0e49",
			904 => x"01930e49",
			905 => x"feee0e49",
			906 => x"08002204",
			907 => x"fead0e49",
			908 => x"0b001b04",
			909 => x"00720e49",
			910 => x"02010b04",
			911 => x"009f0e49",
			912 => x"01960e49",
			913 => x"fe7a0e49",
			914 => x"0d001714",
			915 => x"0500240c",
			916 => x"09001d04",
			917 => x"ffe40ef5",
			918 => x"0a002504",
			919 => x"fffb0ef5",
			920 => x"00520ef5",
			921 => x"09002304",
			922 => x"ff4b0ef5",
			923 => x"00050ef5",
			924 => x"0300403c",
			925 => x"05003928",
			926 => x"04002820",
			927 => x"04002110",
			928 => x"0e008608",
			929 => x"05002904",
			930 => x"ffcb0ef5",
			931 => x"00b40ef5",
			932 => x"04002004",
			933 => x"ffee0ef5",
			934 => x"ff300ef5",
			935 => x"01001408",
			936 => x"0d001904",
			937 => x"001f0ef5",
			938 => x"ff8a0ef5",
			939 => x"08002b04",
			940 => x"00cf0ef5",
			941 => x"ffb70ef5",
			942 => x"01001704",
			943 => x"ff5c0ef5",
			944 => x"00410ef5",
			945 => x"0f00b808",
			946 => x"09002504",
			947 => x"ffa90ef5",
			948 => x"00370ef5",
			949 => x"03003b08",
			950 => x"03002f04",
			951 => x"00120ef5",
			952 => x"00e90ef5",
			953 => x"fff30ef5",
			954 => x"04003604",
			955 => x"00060ef5",
			956 => x"ff7b0ef5",
			957 => x"0d002130",
			958 => x"09001d04",
			959 => x"fecf0f61",
			960 => x"0e00a428",
			961 => x"0201371c",
			962 => x"0f00c710",
			963 => x"0c001808",
			964 => x"04001f04",
			965 => x"ff7e0f61",
			966 => x"01000f61",
			967 => x"08002204",
			968 => x"feda0f61",
			969 => x"ffea0f61",
			970 => x"01001404",
			971 => x"ff630f61",
			972 => x"0f00cf04",
			973 => x"015c0f61",
			974 => x"00510f61",
			975 => x"05003908",
			976 => x"05002f04",
			977 => x"ff9c0f61",
			978 => x"fea90f61",
			979 => x"ffe30f61",
			980 => x"00ed0f61",
			981 => x"06009804",
			982 => x"ff9f0f61",
			983 => x"01560f61",
			984 => x"0d001f50",
			985 => x"0201262c",
			986 => x"0f00b820",
			987 => x"0f00aa1c",
			988 => x"0d001810",
			989 => x"05002408",
			990 => x"03002404",
			991 => x"ffe9103d",
			992 => x"003a103d",
			993 => x"0e007704",
			994 => x"ff9a103d",
			995 => x"0001103d",
			996 => x"0f006504",
			997 => x"ffcc103d",
			998 => x"0c001e04",
			999 => x"00b0103d",
			1000 => x"ffed103d",
			1001 => x"ff6e103d",
			1002 => x"05002e04",
			1003 => x"ffa8103d",
			1004 => x"04002704",
			1005 => x"00b6103d",
			1006 => x"fff5103d",
			1007 => x"04002718",
			1008 => x"0a002c08",
			1009 => x"05002804",
			1010 => x"fff0103d",
			1011 => x"0049103d",
			1012 => x"0500380c",
			1013 => x"05003308",
			1014 => x"05003204",
			1015 => x"ff82103d",
			1016 => x"0029103d",
			1017 => x"ff21103d",
			1018 => x"fff7103d",
			1019 => x"03003508",
			1020 => x"0d001804",
			1021 => x"fff4103d",
			1022 => x"0085103d",
			1023 => x"ffdb103d",
			1024 => x"04002b10",
			1025 => x"08002d08",
			1026 => x"0000f404",
			1027 => x"ffed103d",
			1028 => x"00c7103d",
			1029 => x"0600bc04",
			1030 => x"ffbe103d",
			1031 => x"0037103d",
			1032 => x"0d002004",
			1033 => x"0040103d",
			1034 => x"01001704",
			1035 => x"ff82103d",
			1036 => x"00011604",
			1037 => x"fffb103d",
			1038 => x"001f103d",
			1039 => x"08002750",
			1040 => x"0f00c138",
			1041 => x"07002a10",
			1042 => x"0d001904",
			1043 => x"ff761121",
			1044 => x"03002408",
			1045 => x"0a001e04",
			1046 => x"fffb1121",
			1047 => x"002c1121",
			1048 => x"ffdb1121",
			1049 => x"03003514",
			1050 => x"04002910",
			1051 => x"0a003108",
			1052 => x"0d001504",
			1053 => x"ffdc1121",
			1054 => x"00801121",
			1055 => x"03003104",
			1056 => x"ff901121",
			1057 => x"00351121",
			1058 => x"00ab1121",
			1059 => x"0700380c",
			1060 => x"07003308",
			1061 => x"07003004",
			1062 => x"ffe41121",
			1063 => x"00171121",
			1064 => x"ff861121",
			1065 => x"0b002104",
			1066 => x"00151121",
			1067 => x"fffa1121",
			1068 => x"0a00360c",
			1069 => x"04001b08",
			1070 => x"04001a04",
			1071 => x"ffe61121",
			1072 => x"00211121",
			1073 => x"ff241121",
			1074 => x"07003b08",
			1075 => x"03003104",
			1076 => x"003a1121",
			1077 => x"ff961121",
			1078 => x"005a1121",
			1079 => x"0e008a0c",
			1080 => x"0a003104",
			1081 => x"ffad1121",
			1082 => x"06009504",
			1083 => x"ffec1121",
			1084 => x"00461121",
			1085 => x"02013708",
			1086 => x"0600bd04",
			1087 => x"00f61121",
			1088 => x"fff81121",
			1089 => x"02013c04",
			1090 => x"ffc51121",
			1091 => x"0600c204",
			1092 => x"007a1121",
			1093 => x"0f00e204",
			1094 => x"ffed1121",
			1095 => x"ffff1121",
			1096 => x"08002324",
			1097 => x"0600951c",
			1098 => x"06008010",
			1099 => x"0d001804",
			1100 => x"ff9911dd",
			1101 => x"00009604",
			1102 => x"ffe711dd",
			1103 => x"0d001a04",
			1104 => x"002e11dd",
			1105 => x"fffb11dd",
			1106 => x"05004a08",
			1107 => x"03002404",
			1108 => x"fff611dd",
			1109 => x"006811dd",
			1110 => x"fff511dd",
			1111 => x"04002a04",
			1112 => x"ff6011dd",
			1113 => x"002b11dd",
			1114 => x"07004034",
			1115 => x"0201372c",
			1116 => x"03003118",
			1117 => x"0d001d0c",
			1118 => x"0f00bc08",
			1119 => x"00010404",
			1120 => x"004f11dd",
			1121 => x"ffd511dd",
			1122 => x"00b511dd",
			1123 => x"09002804",
			1124 => x"ffb011dd",
			1125 => x"0000f504",
			1126 => x"fff411dd",
			1127 => x"006811dd",
			1128 => x"05003804",
			1129 => x"ffa411dd",
			1130 => x"03003508",
			1131 => x"0a003804",
			1132 => x"fff011dd",
			1133 => x"007511dd",
			1134 => x"07003804",
			1135 => x"ffb411dd",
			1136 => x"001111dd",
			1137 => x"05003604",
			1138 => x"ffa611dd",
			1139 => x"fff211dd",
			1140 => x"0600a004",
			1141 => x"fff011dd",
			1142 => x"009e11dd",
			1143 => x"07003f50",
			1144 => x"02013744",
			1145 => x"08002218",
			1146 => x"0000d114",
			1147 => x"0200b00c",
			1148 => x"0a002a08",
			1149 => x"0a002804",
			1150 => x"ffdb12a9",
			1151 => x"003212a9",
			1152 => x"ff9b12a9",
			1153 => x"0f008204",
			1154 => x"ffe612a9",
			1155 => x"006412a9",
			1156 => x"ff4312a9",
			1157 => x"09002514",
			1158 => x"04002008",
			1159 => x"07002c04",
			1160 => x"ffef12a9",
			1161 => x"00cf12a9",
			1162 => x"0e008808",
			1163 => x"0000be04",
			1164 => x"fffc12a9",
			1165 => x"ff5512a9",
			1166 => x"005112a9",
			1167 => x"05003810",
			1168 => x"03002708",
			1169 => x"0c002104",
			1170 => x"006c12a9",
			1171 => x"ffe812a9",
			1172 => x"0e008604",
			1173 => x"003312a9",
			1174 => x"ff6b12a9",
			1175 => x"03004604",
			1176 => x"00bd12a9",
			1177 => x"ff9e12a9",
			1178 => x"0e009904",
			1179 => x"ff2412a9",
			1180 => x"03002d04",
			1181 => x"ffab12a9",
			1182 => x"006212a9",
			1183 => x"0c002108",
			1184 => x"0a003b04",
			1185 => x"00bf12a9",
			1186 => x"fffc12a9",
			1187 => x"0d002108",
			1188 => x"03003304",
			1189 => x"ffba12a9",
			1190 => x"000912a9",
			1191 => x"02010a04",
			1192 => x"ffe512a9",
			1193 => x"006812a9",
			1194 => x"0d001708",
			1195 => x"08002204",
			1196 => x"fe73135d",
			1197 => x"ff62135d",
			1198 => x"0900252c",
			1199 => x"03002f18",
			1200 => x"01001414",
			1201 => x"0e00800c",
			1202 => x"09001e04",
			1203 => x"feb2135d",
			1204 => x"06006504",
			1205 => x"fef7135d",
			1206 => x"0192135d",
			1207 => x"04002004",
			1208 => x"00b3135d",
			1209 => x"fe65135d",
			1210 => x"01b5135d",
			1211 => x"0b001b10",
			1212 => x"05003904",
			1213 => x"feea135d",
			1214 => x"0a003b04",
			1215 => x"013b135d",
			1216 => x"09002204",
			1217 => x"ffe4135d",
			1218 => x"fe58135d",
			1219 => x"013c135d",
			1220 => x"0500381c",
			1221 => x"01001710",
			1222 => x"0500330c",
			1223 => x"03002a08",
			1224 => x"08002604",
			1225 => x"fe88135d",
			1226 => x"0042135d",
			1227 => x"014e135d",
			1228 => x"fe3f135d",
			1229 => x"03002e08",
			1230 => x"0d002204",
			1231 => x"fefb135d",
			1232 => x"00fc135d",
			1233 => x"0188135d",
			1234 => x"03004608",
			1235 => x"08002404",
			1236 => x"ffc1135d",
			1237 => x"018a135d",
			1238 => x"fe8c135d",
			1239 => x"07003f58",
			1240 => x"08002644",
			1241 => x"03002f28",
			1242 => x"0f00bc14",
			1243 => x"0f00aa10",
			1244 => x"09001e08",
			1245 => x"05002204",
			1246 => x"00331439",
			1247 => x"ff731439",
			1248 => x"0f006504",
			1249 => x"ffb11439",
			1250 => x"00aa1439",
			1251 => x"ff491439",
			1252 => x"0f00ce08",
			1253 => x"07003304",
			1254 => x"ffcc1439",
			1255 => x"00be1439",
			1256 => x"00014008",
			1257 => x"03002a04",
			1258 => x"fff41439",
			1259 => x"001b1439",
			1260 => x"ff871439",
			1261 => x"0a00380c",
			1262 => x"00012308",
			1263 => x"0f009904",
			1264 => x"ffad1439",
			1265 => x"00401439",
			1266 => x"fef11439",
			1267 => x"05003d04",
			1268 => x"007d1439",
			1269 => x"0b001c04",
			1270 => x"ff461439",
			1271 => x"09002804",
			1272 => x"00351439",
			1273 => x"ffef1439",
			1274 => x"0d001c04",
			1275 => x"00ce1439",
			1276 => x"0a002d04",
			1277 => x"ff391439",
			1278 => x"00013d08",
			1279 => x"0c002204",
			1280 => x"00d71439",
			1281 => x"ffd61439",
			1282 => x"ffd11439",
			1283 => x"0c002108",
			1284 => x"0f00d004",
			1285 => x"000c1439",
			1286 => x"00d71439",
			1287 => x"0d002108",
			1288 => x"09002c04",
			1289 => x"ffc21439",
			1290 => x"000e1439",
			1291 => x"02010a04",
			1292 => x"ffe41439",
			1293 => x"006b1439",
			1294 => x"0700405c",
			1295 => x"03002f28",
			1296 => x"03002a18",
			1297 => x"01001610",
			1298 => x"09001d04",
			1299 => x"ff22150d",
			1300 => x"00012d08",
			1301 => x"0200b004",
			1302 => x"ffdd150d",
			1303 => x"00e6150d",
			1304 => x"ff78150d",
			1305 => x"04001d04",
			1306 => x"006c150d",
			1307 => x"feb7150d",
			1308 => x"09002104",
			1309 => x"ff38150d",
			1310 => x"04001e04",
			1311 => x"ff70150d",
			1312 => x"05003604",
			1313 => x"0129150d",
			1314 => x"0020150d",
			1315 => x"05003914",
			1316 => x"08002610",
			1317 => x"0e00890c",
			1318 => x"0f009904",
			1319 => x"ff8a150d",
			1320 => x"00012d04",
			1321 => x"007a150d",
			1322 => x"ffd2150d",
			1323 => x"feba150d",
			1324 => x"ffda150d",
			1325 => x"03003508",
			1326 => x"09002004",
			1327 => x"ff82150d",
			1328 => x"0113150d",
			1329 => x"0c001f0c",
			1330 => x"00012808",
			1331 => x"00010404",
			1332 => x"ff72150d",
			1333 => x"005d150d",
			1334 => x"ff1a150d",
			1335 => x"05005308",
			1336 => x"0e008504",
			1337 => x"fff2150d",
			1338 => x"00b9150d",
			1339 => x"ff96150d",
			1340 => x"0c002104",
			1341 => x"0127150d",
			1342 => x"05003504",
			1343 => x"ff86150d",
			1344 => x"03005604",
			1345 => x"00a9150d",
			1346 => x"ffea150d",
			1347 => x"07004050",
			1348 => x"0f00ae24",
			1349 => x"07002904",
			1350 => x"fefc15d1",
			1351 => x"04001e0c",
			1352 => x"09001e04",
			1353 => x"ff5615d1",
			1354 => x"0c001b04",
			1355 => x"008215d1",
			1356 => x"ffbb15d1",
			1357 => x"0400360c",
			1358 => x"01000c04",
			1359 => x"ffc015d1",
			1360 => x"06005e04",
			1361 => x"fff315d1",
			1362 => x"014315d1",
			1363 => x"0f009c04",
			1364 => x"ff7415d1",
			1365 => x"000b15d1",
			1366 => x"07003304",
			1367 => x"fed115d1",
			1368 => x"04002110",
			1369 => x"0400200c",
			1370 => x"0a003108",
			1371 => x"04001804",
			1372 => x"ffd115d1",
			1373 => x"013515d1",
			1374 => x"ff7f15d1",
			1375 => x"fea515d1",
			1376 => x"04002608",
			1377 => x"02013704",
			1378 => x"013b15d1",
			1379 => x"fff715d1",
			1380 => x"08002608",
			1381 => x"05003904",
			1382 => x"fedd15d1",
			1383 => x"002b15d1",
			1384 => x"0d002004",
			1385 => x"012315d1",
			1386 => x"ff5415d1",
			1387 => x"0c002104",
			1388 => x"013f15d1",
			1389 => x"0d002108",
			1390 => x"05004104",
			1391 => x"ff6c15d1",
			1392 => x"001115d1",
			1393 => x"02010a04",
			1394 => x"ffd115d1",
			1395 => x"00ca15d1",
			1396 => x"07003f58",
			1397 => x"0201374c",
			1398 => x"08002220",
			1399 => x"0000d114",
			1400 => x"0200b00c",
			1401 => x"0a002a08",
			1402 => x"0a002804",
			1403 => x"ffdc16ad",
			1404 => x"003116ad",
			1405 => x"ff9f16ad",
			1406 => x"0f008204",
			1407 => x"ffe716ad",
			1408 => x"006216ad",
			1409 => x"06009008",
			1410 => x"06008a04",
			1411 => x"ffa216ad",
			1412 => x"003d16ad",
			1413 => x"ff3b16ad",
			1414 => x"0d001d1c",
			1415 => x"0f00b810",
			1416 => x"0a002d08",
			1417 => x"07002c04",
			1418 => x"ffed16ad",
			1419 => x"007216ad",
			1420 => x"0d001c04",
			1421 => x"ff5716ad",
			1422 => x"003816ad",
			1423 => x"07003704",
			1424 => x"fffa16ad",
			1425 => x"03003104",
			1426 => x"00e716ad",
			1427 => x"002816ad",
			1428 => x"0f00c30c",
			1429 => x"03004608",
			1430 => x"06008504",
			1431 => x"ffe116ad",
			1432 => x"00b716ad",
			1433 => x"ffa916ad",
			1434 => x"ff8d16ad",
			1435 => x"0e009904",
			1436 => x"ff2e16ad",
			1437 => x"03002d04",
			1438 => x"ffac16ad",
			1439 => x"005d16ad",
			1440 => x"0c002108",
			1441 => x"0a003b04",
			1442 => x"00ba16ad",
			1443 => x"fffc16ad",
			1444 => x"0d002108",
			1445 => x"03003304",
			1446 => x"ffc016ad",
			1447 => x"000816ad",
			1448 => x"02010a04",
			1449 => x"ffe616ad",
			1450 => x"006416ad",
			1451 => x"08001f04",
			1452 => x"fed61749",
			1453 => x"00012224",
			1454 => x"07002904",
			1455 => x"feeb1749",
			1456 => x"0a003714",
			1457 => x"04001e0c",
			1458 => x"0a002708",
			1459 => x"05001f04",
			1460 => x"ffa01749",
			1461 => x"00b71749",
			1462 => x"ff631749",
			1463 => x"06008004",
			1464 => x"00801749",
			1465 => x"01621749",
			1466 => x"04002b04",
			1467 => x"ff0f1749",
			1468 => x"04003804",
			1469 => x"00d51749",
			1470 => x"ff8a1749",
			1471 => x"08002308",
			1472 => x"00014b04",
			1473 => x"fe891749",
			1474 => x"004a1749",
			1475 => x"09002b18",
			1476 => x"0500380c",
			1477 => x"05003608",
			1478 => x"0d001d04",
			1479 => x"00a81749",
			1480 => x"ff7d1749",
			1481 => x"fef51749",
			1482 => x"07003b08",
			1483 => x"05003c04",
			1484 => x"003a1749",
			1485 => x"ff8b1749",
			1486 => x"01421749",
			1487 => x"0f00bf04",
			1488 => x"ffd11749",
			1489 => x"01571749",
			1490 => x"09001d04",
			1491 => x"fe9a17e5",
			1492 => x"03002710",
			1493 => x"06006504",
			1494 => x"ff0317e5",
			1495 => x"08001f04",
			1496 => x"ff4b17e5",
			1497 => x"00012c04",
			1498 => x"016217e5",
			1499 => x"00c117e5",
			1500 => x"08002214",
			1501 => x"0b001504",
			1502 => x"00d617e5",
			1503 => x"07003c0c",
			1504 => x"0a002f08",
			1505 => x"03002a04",
			1506 => x"007f17e5",
			1507 => x"ffbc17e5",
			1508 => x"fe6e17e5",
			1509 => x"008517e5",
			1510 => x"0400210c",
			1511 => x"04002008",
			1512 => x"0a003104",
			1513 => x"017317e5",
			1514 => x"ff4e17e5",
			1515 => x"fe9f17e5",
			1516 => x"0700350c",
			1517 => x"06009908",
			1518 => x"0f006504",
			1519 => x"ff4017e5",
			1520 => x"00fa17e5",
			1521 => x"fee117e5",
			1522 => x"02013008",
			1523 => x"03003804",
			1524 => x"019417e5",
			1525 => x"ffaf17e5",
			1526 => x"01001904",
			1527 => x"ffae17e5",
			1528 => x"015017e5",
			1529 => x"0d001708",
			1530 => x"08002204",
			1531 => x"fe6d1891",
			1532 => x"ff5e1891",
			1533 => x"07003f40",
			1534 => x"02013738",
			1535 => x"09002518",
			1536 => x"03003410",
			1537 => x"09002408",
			1538 => x"06009704",
			1539 => x"01261891",
			1540 => x"ffd31891",
			1541 => x"0000d804",
			1542 => x"ff9f1891",
			1543 => x"01dd1891",
			1544 => x"03003b04",
			1545 => x"fe4f1891",
			1546 => x"ff641891",
			1547 => x"04002110",
			1548 => x"0d001f08",
			1549 => x"0c002104",
			1550 => x"fdda1891",
			1551 => x"ff5c1891",
			1552 => x"0c002404",
			1553 => x"01111891",
			1554 => x"ff101891",
			1555 => x"08002608",
			1556 => x"0c001e04",
			1557 => x"00921891",
			1558 => x"fe9b1891",
			1559 => x"0c002204",
			1560 => x"018e1891",
			1561 => x"fed91891",
			1562 => x"0600b704",
			1563 => x"fe3f1891",
			1564 => x"ffc41891",
			1565 => x"05003508",
			1566 => x"0600c104",
			1567 => x"01511891",
			1568 => x"ff891891",
			1569 => x"03005304",
			1570 => x"01961891",
			1571 => x"ff181891",
			1572 => x"0d002144",
			1573 => x"07002904",
			1574 => x"fec81925",
			1575 => x"0f00aa1c",
			1576 => x"06008110",
			1577 => x"0e00650c",
			1578 => x"03002f08",
			1579 => x"0c001b04",
			1580 => x"01441925",
			1581 => x"ffb01925",
			1582 => x"ff201925",
			1583 => x"feef1925",
			1584 => x"01000c04",
			1585 => x"ffa31925",
			1586 => x"05004c04",
			1587 => x"01561925",
			1588 => x"00191925",
			1589 => x"07003304",
			1590 => x"feb51925",
			1591 => x"03002e10",
			1592 => x"08002408",
			1593 => x"00011a04",
			1594 => x"ff551925",
			1595 => x"01131925",
			1596 => x"08002704",
			1597 => x"fee41925",
			1598 => x"ffd11925",
			1599 => x"08002608",
			1600 => x"04002604",
			1601 => x"00ac1925",
			1602 => x"ff8c1925",
			1603 => x"0a003e04",
			1604 => x"016f1925",
			1605 => x"fff21925",
			1606 => x"06009804",
			1607 => x"ff9a1925",
			1608 => x"01611925",
			1609 => x"07003f64",
			1610 => x"0800264c",
			1611 => x"03002f30",
			1612 => x"0e008b1c",
			1613 => x"0f00aa10",
			1614 => x"09001e08",
			1615 => x"05002204",
			1616 => x"00351a11",
			1617 => x"ff6d1a11",
			1618 => x"0f006504",
			1619 => x"ffae1a11",
			1620 => x"00b11a11",
			1621 => x"01001008",
			1622 => x"01000c04",
			1623 => x"ffdf1a11",
			1624 => x"00231a11",
			1625 => x"ff3b1a11",
			1626 => x"0f00ce08",
			1627 => x"0c001704",
			1628 => x"ffee1a11",
			1629 => x"00bb1a11",
			1630 => x"00014008",
			1631 => x"03002a04",
			1632 => x"fff41a11",
			1633 => x"001c1a11",
			1634 => x"ff851a11",
			1635 => x"0a00380c",
			1636 => x"00012308",
			1637 => x"0f009904",
			1638 => x"ffaa1a11",
			1639 => x"003f1a11",
			1640 => x"fee91a11",
			1641 => x"05003d04",
			1642 => x"00841a11",
			1643 => x"0b001c04",
			1644 => x"ff3a1a11",
			1645 => x"09002804",
			1646 => x"00371a11",
			1647 => x"ffef1a11",
			1648 => x"0d001c04",
			1649 => x"00d41a11",
			1650 => x"0a002d04",
			1651 => x"ff321a11",
			1652 => x"07003e0c",
			1653 => x"0a004808",
			1654 => x"04002704",
			1655 => x"00291a11",
			1656 => x"00d61a11",
			1657 => x"ffc21a11",
			1658 => x"ff9d1a11",
			1659 => x"0c002104",
			1660 => x"00db1a11",
			1661 => x"0d002108",
			1662 => x"09002c04",
			1663 => x"ffbe1a11",
			1664 => x"000e1a11",
			1665 => x"02010a04",
			1666 => x"ffe41a11",
			1667 => x"006f1a11",
			1668 => x"09001d04",
			1669 => x"fea01acf",
			1670 => x"0300270c",
			1671 => x"06006504",
			1672 => x"ff0f1acf",
			1673 => x"08001f04",
			1674 => x"ff551acf",
			1675 => x"012b1acf",
			1676 => x"05003a2c",
			1677 => x"02012118",
			1678 => x"05002d08",
			1679 => x"0b001b04",
			1680 => x"00151acf",
			1681 => x"feab1acf",
			1682 => x"0e008808",
			1683 => x"05002f04",
			1684 => x"01341acf",
			1685 => x"ff6c1acf",
			1686 => x"05003504",
			1687 => x"018f1acf",
			1688 => x"00881acf",
			1689 => x"0d001b04",
			1690 => x"fe811acf",
			1691 => x"03002e08",
			1692 => x"0d002104",
			1693 => x"fefa1acf",
			1694 => x"01041acf",
			1695 => x"03003104",
			1696 => x"016e1acf",
			1697 => x"ff8c1acf",
			1698 => x"0300350c",
			1699 => x"09002004",
			1700 => x"ff5a1acf",
			1701 => x"08002304",
			1702 => x"00921acf",
			1703 => x"017a1acf",
			1704 => x"07003b10",
			1705 => x"0b001b08",
			1706 => x"07003304",
			1707 => x"ff7c1acf",
			1708 => x"feaa1acf",
			1709 => x"0f009f04",
			1710 => x"ff651acf",
			1711 => x"00da1acf",
			1712 => x"03004b04",
			1713 => x"013f1acf",
			1714 => x"ff8e1acf",
			1715 => x"01001220",
			1716 => x"08002210",
			1717 => x"01000e04",
			1718 => x"fe431b51",
			1719 => x"0b001508",
			1720 => x"0b001404",
			1721 => x"fe4b1b51",
			1722 => x"ffe31b51",
			1723 => x"fe3f1b51",
			1724 => x"0c001b08",
			1725 => x"0f00bd04",
			1726 => x"04151b51",
			1727 => x"ffe51b51",
			1728 => x"0c001d04",
			1729 => x"ffe61b51",
			1730 => x"fe421b51",
			1731 => x"0f008908",
			1732 => x"09002304",
			1733 => x"01051b51",
			1734 => x"fe441b51",
			1735 => x"0d001904",
			1736 => x"ff7b1b51",
			1737 => x"0a004314",
			1738 => x"0500390c",
			1739 => x"00012204",
			1740 => x"03a61b51",
			1741 => x"08002604",
			1742 => x"00331b51",
			1743 => x"02891b51",
			1744 => x"08002604",
			1745 => x"03741b51",
			1746 => x"02f11b51",
			1747 => x"01341b51",
			1748 => x"01000e08",
			1749 => x"08002304",
			1750 => x"fe651bc5",
			1751 => x"010a1bc5",
			1752 => x"07003f24",
			1753 => x"02013718",
			1754 => x"06005e04",
			1755 => x"fe711bc5",
			1756 => x"0000d304",
			1757 => x"01841bc5",
			1758 => x"08002608",
			1759 => x"04002004",
			1760 => x"00751bc5",
			1761 => x"ff3a1bc5",
			1762 => x"0c002204",
			1763 => x"01041bc5",
			1764 => x"feab1bc5",
			1765 => x"00015108",
			1766 => x"0f00cf04",
			1767 => x"fec31bc5",
			1768 => x"fe0f1bc5",
			1769 => x"00161bc5",
			1770 => x"05003508",
			1771 => x"07004404",
			1772 => x"ff6d1bc5",
			1773 => x"01871bc5",
			1774 => x"03005304",
			1775 => x"01b51bc5",
			1776 => x"feb61bc5",
			1777 => x"01001430",
			1778 => x"01001220",
			1779 => x"01001014",
			1780 => x"01000e08",
			1781 => x"08002304",
			1782 => x"fe2e1c69",
			1783 => x"feb11c69",
			1784 => x"0f008c04",
			1785 => x"fe2f1c69",
			1786 => x"0600ab04",
			1787 => x"01441c69",
			1788 => x"fe351c69",
			1789 => x"0f008204",
			1790 => x"fe2f1c69",
			1791 => x"00012e04",
			1792 => x"02771c69",
			1793 => x"ff261c69",
			1794 => x"0f008208",
			1795 => x"06006504",
			1796 => x"fe2f1c69",
			1797 => x"ff181c69",
			1798 => x"05003804",
			1799 => x"00b71c69",
			1800 => x"04b01c69",
			1801 => x"0f009308",
			1802 => x"09002c04",
			1803 => x"ff101c69",
			1804 => x"fe2f1c69",
			1805 => x"0b001a04",
			1806 => x"01b31c69",
			1807 => x"03002a08",
			1808 => x"0d001f04",
			1809 => x"012a1c69",
			1810 => x"061c1c69",
			1811 => x"00013d04",
			1812 => x"06071c69",
			1813 => x"0e009904",
			1814 => x"03081c69",
			1815 => x"03002f04",
			1816 => x"04c31c69",
			1817 => x"05fb1c69",
			1818 => x"08002634",
			1819 => x"02011c24",
			1820 => x"02010d18",
			1821 => x"0f00ae14",
			1822 => x"07002904",
			1823 => x"fee91d15",
			1824 => x"03002f08",
			1825 => x"04001e04",
			1826 => x"00031d15",
			1827 => x"011b1d15",
			1828 => x"0f009904",
			1829 => x"ff281d15",
			1830 => x"00711d15",
			1831 => x"feac1d15",
			1832 => x"0600af08",
			1833 => x"07003204",
			1834 => x"ff9a1d15",
			1835 => x"012d1d15",
			1836 => x"fefd1d15",
			1837 => x"0d001b08",
			1838 => x"05003a04",
			1839 => x"fe881d15",
			1840 => x"002a1d15",
			1841 => x"0c001d04",
			1842 => x"007b1d15",
			1843 => x"ff6e1d15",
			1844 => x"0a003b18",
			1845 => x"02013710",
			1846 => x"0e007e08",
			1847 => x"07003504",
			1848 => x"ff6f1d15",
			1849 => x"ffff1d15",
			1850 => x"0600bc04",
			1851 => x"017f1d15",
			1852 => x"00101d15",
			1853 => x"03002e04",
			1854 => x"ff221d15",
			1855 => x"01141d15",
			1856 => x"05003e04",
			1857 => x"fecf1d15",
			1858 => x"03004604",
			1859 => x"00e91d15",
			1860 => x"ff691d15",
			1861 => x"0a003120",
			1862 => x"09001e0c",
			1863 => x"0000b808",
			1864 => x"06008004",
			1865 => x"fff41dd1",
			1866 => x"001f1dd1",
			1867 => x"ffba1dd1",
			1868 => x"06006504",
			1869 => x"ffda1dd1",
			1870 => x"0d001704",
			1871 => x"ffeb1dd1",
			1872 => x"05003308",
			1873 => x"02013504",
			1874 => x"00911dd1",
			1875 => x"000e1dd1",
			1876 => x"fff61dd1",
			1877 => x"0500381c",
			1878 => x"02011a10",
			1879 => x"06009e08",
			1880 => x"07002d04",
			1881 => x"000b1dd1",
			1882 => x"ffba1dd1",
			1883 => x"08002004",
			1884 => x"fff71dd1",
			1885 => x"00701dd1",
			1886 => x"09002b08",
			1887 => x"0e00a304",
			1888 => x"ff721dd1",
			1889 => x"fffa1dd1",
			1890 => x"002e1dd1",
			1891 => x"03003510",
			1892 => x"09002208",
			1893 => x"0f00ba04",
			1894 => x"ffe01dd1",
			1895 => x"00031dd1",
			1896 => x"00014f04",
			1897 => x"00871dd1",
			1898 => x"00071dd1",
			1899 => x"0600b710",
			1900 => x"01001608",
			1901 => x"0a003904",
			1902 => x"00021dd1",
			1903 => x"ffa01dd1",
			1904 => x"0a004704",
			1905 => x"00191dd1",
			1906 => x"ffee1dd1",
			1907 => x"00281dd1",
			1908 => x"0d00170c",
			1909 => x"08001f04",
			1910 => x"fe621e3d",
			1911 => x"05002204",
			1912 => x"013c1e3d",
			1913 => x"fe6b1e3d",
			1914 => x"0f006504",
			1915 => x"fe681e3d",
			1916 => x"03004624",
			1917 => x"07003f14",
			1918 => x"0201370c",
			1919 => x"0000d304",
			1920 => x"021d1e3d",
			1921 => x"09002004",
			1922 => x"fe281e3d",
			1923 => x"00b41e3d",
			1924 => x"0600b704",
			1925 => x"fe181e3d",
			1926 => x"ffe91e3d",
			1927 => x"0f00db08",
			1928 => x"0b001e04",
			1929 => x"02101e3d",
			1930 => x"01aa1e3d",
			1931 => x"04002b04",
			1932 => x"019d1e3d",
			1933 => x"00101e3d",
			1934 => x"fe521e3d",
			1935 => x"0d001710",
			1936 => x"09002308",
			1937 => x"08002204",
			1938 => x"fe781ed1",
			1939 => x"ff371ed1",
			1940 => x"05004404",
			1941 => x"00821ed1",
			1942 => x"ffa61ed1",
			1943 => x"0a003b28",
			1944 => x"05003a20",
			1945 => x"0d002118",
			1946 => x"02013510",
			1947 => x"08002708",
			1948 => x"0c001e04",
			1949 => x"00451ed1",
			1950 => x"fedd1ed1",
			1951 => x"0e008a04",
			1952 => x"00331ed1",
			1953 => x"01961ed1",
			1954 => x"07003e04",
			1955 => x"fe751ed1",
			1956 => x"ffd91ed1",
			1957 => x"00011404",
			1958 => x"ff591ed1",
			1959 => x"017d1ed1",
			1960 => x"0f00ad04",
			1961 => x"00591ed1",
			1962 => x"01921ed1",
			1963 => x"0e009910",
			1964 => x"0001380c",
			1965 => x"0d001b04",
			1966 => x"fe6d1ed1",
			1967 => x"03004604",
			1968 => x"01491ed1",
			1969 => x"fed81ed1",
			1970 => x"fe5e1ed1",
			1971 => x"01521ed1",
			1972 => x"0d001710",
			1973 => x"08001f04",
			1974 => x"fe681f45",
			1975 => x"05002404",
			1976 => x"013f1f45",
			1977 => x"05003604",
			1978 => x"fe6b1f45",
			1979 => x"ff151f45",
			1980 => x"0f006504",
			1981 => x"fe7a1f45",
			1982 => x"05005624",
			1983 => x"05003810",
			1984 => x"0f00ae04",
			1985 => x"017d1f45",
			1986 => x"09002104",
			1987 => x"fe471f45",
			1988 => x"05003604",
			1989 => x"00641f45",
			1990 => x"feec1f45",
			1991 => x"0700380c",
			1992 => x"03003404",
			1993 => x"00e71f45",
			1994 => x"03003b04",
			1995 => x"fe0b1f45",
			1996 => x"ff381f45",
			1997 => x"0a004304",
			1998 => x"01ab1f45",
			1999 => x"00921f45",
			2000 => x"fe781f45",
			2001 => x"01001220",
			2002 => x"08002210",
			2003 => x"01000e04",
			2004 => x"fe501fd9",
			2005 => x"0b001708",
			2006 => x"09001d04",
			2007 => x"fe511fd9",
			2008 => x"012f1fd9",
			2009 => x"fe511fd9",
			2010 => x"0c001d0c",
			2011 => x"07002c04",
			2012 => x"fe551fd9",
			2013 => x"02012904",
			2014 => x"02e81fd9",
			2015 => x"00681fd9",
			2016 => x"fe521fd9",
			2017 => x"0f008708",
			2018 => x"0b001c04",
			2019 => x"ff5d1fd9",
			2020 => x"fe531fd9",
			2021 => x"0d001904",
			2022 => x"ffbb1fd9",
			2023 => x"0400381c",
			2024 => x"05003810",
			2025 => x"02013708",
			2026 => x"03002f04",
			2027 => x"02391fd9",
			2028 => x"00f81fd9",
			2029 => x"0d001f04",
			2030 => x"fe861fd9",
			2031 => x"01d61fd9",
			2032 => x"0c001c04",
			2033 => x"01941fd9",
			2034 => x"01001704",
			2035 => x"025c1fd9",
			2036 => x"022e1fd9",
			2037 => x"006c1fd9",
			2038 => x"0a003120",
			2039 => x"09001e0c",
			2040 => x"0000b808",
			2041 => x"06008004",
			2042 => x"fff420a5",
			2043 => x"001e20a5",
			2044 => x"ffbc20a5",
			2045 => x"06006504",
			2046 => x"ffdb20a5",
			2047 => x"0d001704",
			2048 => x"ffec20a5",
			2049 => x"05003308",
			2050 => x"02013504",
			2051 => x"008b20a5",
			2052 => x"000d20a5",
			2053 => x"fff820a5",
			2054 => x"05003820",
			2055 => x"02011a10",
			2056 => x"06009e08",
			2057 => x"07002d04",
			2058 => x"000b20a5",
			2059 => x"ffbd20a5",
			2060 => x"05003004",
			2061 => x"fff720a5",
			2062 => x"006b20a5",
			2063 => x"09002b0c",
			2064 => x"05003308",
			2065 => x"05003004",
			2066 => x"ffd220a5",
			2067 => x"001f20a5",
			2068 => x"ff7120a5",
			2069 => x"002d20a5",
			2070 => x"03003514",
			2071 => x"09002208",
			2072 => x"0f00ba04",
			2073 => x"ffe120a5",
			2074 => x"000320a5",
			2075 => x"01001804",
			2076 => x"008120a5",
			2077 => x"00014d04",
			2078 => x"001620a5",
			2079 => x"ffee20a5",
			2080 => x"0600b710",
			2081 => x"01001608",
			2082 => x"0a003904",
			2083 => x"000220a5",
			2084 => x"ffa320a5",
			2085 => x"0a004704",
			2086 => x"001820a5",
			2087 => x"ffef20a5",
			2088 => x"002720a5",
			2089 => x"0d001710",
			2090 => x"05002208",
			2091 => x"0a002704",
			2092 => x"fff32151",
			2093 => x"001e2151",
			2094 => x"09002304",
			2095 => x"ff9c2151",
			2096 => x"00032151",
			2097 => x"04002b2c",
			2098 => x"0d001f24",
			2099 => x"0c001e14",
			2100 => x"02013710",
			2101 => x"08002308",
			2102 => x"0c001904",
			2103 => x"00462151",
			2104 => x"ffab2151",
			2105 => x"0e008804",
			2106 => x"fff12151",
			2107 => x"00bd2151",
			2108 => x"ffbe2151",
			2109 => x"0a002c08",
			2110 => x"07003304",
			2111 => x"fff92151",
			2112 => x"00232151",
			2113 => x"0f00c304",
			2114 => x"001e2151",
			2115 => x"ff7a2151",
			2116 => x"0000f404",
			2117 => x"ffeb2151",
			2118 => x"00972151",
			2119 => x"04002e0c",
			2120 => x"01001908",
			2121 => x"00012904",
			2122 => x"ffff2151",
			2123 => x"ff9e2151",
			2124 => x"000f2151",
			2125 => x"03004008",
			2126 => x"00010404",
			2127 => x"fff52151",
			2128 => x"006b2151",
			2129 => x"01001704",
			2130 => x"ffc72151",
			2131 => x"00012151",
			2132 => x"0d001714",
			2133 => x"0500240c",
			2134 => x"09001d04",
			2135 => x"ffe521ed",
			2136 => x"0a002504",
			2137 => x"fffb21ed",
			2138 => x"004e21ed",
			2139 => x"09002304",
			2140 => x"ff5121ed",
			2141 => x"000521ed",
			2142 => x"0a004334",
			2143 => x"05003924",
			2144 => x"0400281c",
			2145 => x"0d001f10",
			2146 => x"02012608",
			2147 => x"0f00b804",
			2148 => x"ffdd21ed",
			2149 => x"008221ed",
			2150 => x"05003304",
			2151 => x"001621ed",
			2152 => x"ff4e21ed",
			2153 => x"08002d08",
			2154 => x"0000f404",
			2155 => x"ffef21ed",
			2156 => x"00d421ed",
			2157 => x"ffc421ed",
			2158 => x"01001704",
			2159 => x"ff6921ed",
			2160 => x"003e21ed",
			2161 => x"0f00b808",
			2162 => x"0d001b04",
			2163 => x"ffa921ed",
			2164 => x"002f21ed",
			2165 => x"0600c604",
			2166 => x"00dd21ed",
			2167 => x"000121ed",
			2168 => x"07004104",
			2169 => x"ff8a21ed",
			2170 => x"000821ed",
			2171 => x"07004038",
			2172 => x"0201372c",
			2173 => x"0f00cd24",
			2174 => x"00013c20",
			2175 => x"07003a10",
			2176 => x"02011c08",
			2177 => x"0f00b804",
			2178 => x"ffde2279",
			2179 => x"006d2279",
			2180 => x"0a003804",
			2181 => x"ff642279",
			2182 => x"001f2279",
			2183 => x"00012508",
			2184 => x"00011a04",
			2185 => x"00212279",
			2186 => x"ffa02279",
			2187 => x"09002904",
			2188 => x"00af2279",
			2189 => x"fffa2279",
			2190 => x"ff762279",
			2191 => x"0c001704",
			2192 => x"fff42279",
			2193 => x"007c2279",
			2194 => x"03002e04",
			2195 => x"ff672279",
			2196 => x"0600b704",
			2197 => x"ffa12279",
			2198 => x"005c2279",
			2199 => x"0600a304",
			2200 => x"ffed2279",
			2201 => x"01001a04",
			2202 => x"00922279",
			2203 => x"01001c04",
			2204 => x"ffe82279",
			2205 => x"00282279",
			2206 => x"0d001708",
			2207 => x"08002204",
			2208 => x"fe7a22f5",
			2209 => x"ff7e22f5",
			2210 => x"08002b30",
			2211 => x"0c002118",
			2212 => x"07003e14",
			2213 => x"02013710",
			2214 => x"03003508",
			2215 => x"0a003804",
			2216 => x"001b22f5",
			2217 => x"014a22f5",
			2218 => x"0d001b04",
			2219 => x"fe9e22f5",
			2220 => x"003822f5",
			2221 => x"fe7e22f5",
			2222 => x"016322f5",
			2223 => x"01001710",
			2224 => x"0b00200c",
			2225 => x"04003b08",
			2226 => x"07002e04",
			2227 => x"ffbe22f5",
			2228 => x"00f122f5",
			2229 => x"ff6022f5",
			2230 => x"fe2b22f5",
			2231 => x"0e009d04",
			2232 => x"013222f5",
			2233 => x"ff4e22f5",
			2234 => x"00011604",
			2235 => x"ff9722f5",
			2236 => x"017422f5",
			2237 => x"08002320",
			2238 => x"01000e04",
			2239 => x"fe632391",
			2240 => x"0f00ba14",
			2241 => x"0f006c04",
			2242 => x"fe712391",
			2243 => x"03003408",
			2244 => x"0d001704",
			2245 => x"ffa02391",
			2246 => x"01bd2391",
			2247 => x"08002204",
			2248 => x"fe7a2391",
			2249 => x"ffdc2391",
			2250 => x"0e00a004",
			2251 => x"fe292391",
			2252 => x"00612391",
			2253 => x"0300452c",
			2254 => x"0500381c",
			2255 => x"0c001e08",
			2256 => x"0b001a04",
			2257 => x"00452391",
			2258 => x"01c02391",
			2259 => x"0100170c",
			2260 => x"01001608",
			2261 => x"01001404",
			2262 => x"fe1a2391",
			2263 => x"013c2391",
			2264 => x"fd7c2391",
			2265 => x"09002a04",
			2266 => x"fff82391",
			2267 => x"01a42391",
			2268 => x"0c001c04",
			2269 => x"00402391",
			2270 => x"00014f08",
			2271 => x"02010b04",
			2272 => x"00ef2391",
			2273 => x"01ad2391",
			2274 => x"00f82391",
			2275 => x"fe522391",
			2276 => x"08001f10",
			2277 => x"01000e04",
			2278 => x"fe8a2425",
			2279 => x"03002904",
			2280 => x"feed2425",
			2281 => x"03002f04",
			2282 => x"008c2425",
			2283 => x"ff612425",
			2284 => x"0300270c",
			2285 => x"06006504",
			2286 => x"ff0e2425",
			2287 => x"0a002a04",
			2288 => x"016b2425",
			2289 => x"00a62425",
			2290 => x"05002d08",
			2291 => x"0b001e04",
			2292 => x"fea32425",
			2293 => x"00482425",
			2294 => x"0a003108",
			2295 => x"04002304",
			2296 => x"014b2425",
			2297 => x"ffe82425",
			2298 => x"05003810",
			2299 => x"03002f08",
			2300 => x"0f00cb04",
			2301 => x"00b52425",
			2302 => x"ff152425",
			2303 => x"01001704",
			2304 => x"fea32425",
			2305 => x"01312425",
			2306 => x"0a004308",
			2307 => x"08002404",
			2308 => x"fffa2425",
			2309 => x"015a2425",
			2310 => x"08002604",
			2311 => x"feab2425",
			2312 => x"ffca2425",
			2313 => x"08002010",
			2314 => x"01000e04",
			2315 => x"fe672499",
			2316 => x"0000f308",
			2317 => x"06006d04",
			2318 => x"fe862499",
			2319 => x"018f2499",
			2320 => x"fe752499",
			2321 => x"0f006504",
			2322 => x"fe7b2499",
			2323 => x"01001b24",
			2324 => x"03004620",
			2325 => x"05003810",
			2326 => x"0f00c008",
			2327 => x"01001404",
			2328 => x"00602499",
			2329 => x"01d32499",
			2330 => x"0c001d04",
			2331 => x"00812499",
			2332 => x"fee72499",
			2333 => x"07003808",
			2334 => x"0a003b04",
			2335 => x"00d42499",
			2336 => x"fe5a2499",
			2337 => x"03003b04",
			2338 => x"01b22499",
			2339 => x"00be2499",
			2340 => x"fe722499",
			2341 => x"01982499",
			2342 => x"01000e08",
			2343 => x"08002304",
			2344 => x"fe852535",
			2345 => x"00bc2535",
			2346 => x"02013734",
			2347 => x"0a003b20",
			2348 => x"08002714",
			2349 => x"01001810",
			2350 => x"07003508",
			2351 => x"0f00aa04",
			2352 => x"00c22535",
			2353 => x"ff272535",
			2354 => x"09002504",
			2355 => x"01512535",
			2356 => x"ffd82535",
			2357 => x"fee42535",
			2358 => x"0600bd08",
			2359 => x"06008504",
			2360 => x"ff7b2535",
			2361 => x"018f2535",
			2362 => x"fff22535",
			2363 => x"05003f04",
			2364 => x"feb72535",
			2365 => x"03004108",
			2366 => x"04003504",
			2367 => x"01362535",
			2368 => x"00392535",
			2369 => x"01001704",
			2370 => x"fed22535",
			2371 => x"00352535",
			2372 => x"0e00a40c",
			2373 => x"0c002208",
			2374 => x"03003104",
			2375 => x"fe9c2535",
			2376 => x"ff9c2535",
			2377 => x"010f2535",
			2378 => x"02014704",
			2379 => x"015f2535",
			2380 => x"ff8d2535",
			2381 => x"0d001708",
			2382 => x"08002204",
			2383 => x"fe7525d9",
			2384 => x"ff6e25d9",
			2385 => x"09002528",
			2386 => x"03002f14",
			2387 => x"02013710",
			2388 => x"09001e04",
			2389 => x"feb525d9",
			2390 => x"0f006504",
			2391 => x"fee125d9",
			2392 => x"09002104",
			2393 => x"00a825d9",
			2394 => x"01ae25d9",
			2395 => x"feaf25d9",
			2396 => x"0700340c",
			2397 => x"0c001b04",
			2398 => x"fe6a25d9",
			2399 => x"0c001c04",
			2400 => x"006325d9",
			2401 => x"ffe025d9",
			2402 => x"01001204",
			2403 => x"00f325d9",
			2404 => x"ffa425d9",
			2405 => x"05003818",
			2406 => x"07004414",
			2407 => x"0a003108",
			2408 => x"07003a04",
			2409 => x"fe8425d9",
			2410 => x"007e25d9",
			2411 => x"0e008604",
			2412 => x"00e825d9",
			2413 => x"01001704",
			2414 => x"fe7525d9",
			2415 => x"ff7625d9",
			2416 => x"013525d9",
			2417 => x"03004608",
			2418 => x"08002404",
			2419 => x"ffcc25d9",
			2420 => x"018525d9",
			2421 => x"fe9725d9",
			2422 => x"07004050",
			2423 => x"0f00ae1c",
			2424 => x"06008010",
			2425 => x"0d001704",
			2426 => x"fed5269d",
			2427 => x"0c001904",
			2428 => x"0095269d",
			2429 => x"0f008204",
			2430 => x"ff0c269d",
			2431 => x"001f269d",
			2432 => x"01000c04",
			2433 => x"ff9f269d",
			2434 => x"04003604",
			2435 => x"0146269d",
			2436 => x"0005269d",
			2437 => x"05003a24",
			2438 => x"0800261c",
			2439 => x"0400200c",
			2440 => x"00011904",
			2441 => x"fec4269d",
			2442 => x"0f00ce04",
			2443 => x"00ea269d",
			2444 => x"feed269d",
			2445 => x"0b001808",
			2446 => x"07003404",
			2447 => x"ff24269d",
			2448 => x"00b1269d",
			2449 => x"05003304",
			2450 => x"ff8d269d",
			2451 => x"fe9d269d",
			2452 => x"0f00c304",
			2453 => x"00db269d",
			2454 => x"ffbe269d",
			2455 => x"03003508",
			2456 => x"0d001a04",
			2457 => x"007a269d",
			2458 => x"014c269d",
			2459 => x"0c001f04",
			2460 => x"ff12269d",
			2461 => x"0069269d",
			2462 => x"0c002104",
			2463 => x"0159269d",
			2464 => x"0d002108",
			2465 => x"03003304",
			2466 => x"ff48269d",
			2467 => x"0022269d",
			2468 => x"00011404",
			2469 => x"ffcc269d",
			2470 => x"00de269d",
			2471 => x"0d001b34",
			2472 => x"0c001a24",
			2473 => x"0900211c",
			2474 => x"0200ca14",
			2475 => x"0400210c",
			2476 => x"09001d04",
			2477 => x"ffe42781",
			2478 => x"00009604",
			2479 => x"fffb2781",
			2480 => x"00782781",
			2481 => x"0000ca04",
			2482 => x"ffbc2781",
			2483 => x"00192781",
			2484 => x"05003a04",
			2485 => x"ff8a2781",
			2486 => x"00152781",
			2487 => x"07002c04",
			2488 => x"ffee2781",
			2489 => x"00812781",
			2490 => x"05003a04",
			2491 => x"ff632781",
			2492 => x"0a003b04",
			2493 => x"004b2781",
			2494 => x"07003904",
			2495 => x"ffb12781",
			2496 => x"00152781",
			2497 => x"0400211c",
			2498 => x"08002408",
			2499 => x"07003204",
			2500 => x"fff62781",
			2501 => x"00532781",
			2502 => x"08002a10",
			2503 => x"04001a08",
			2504 => x"04001804",
			2505 => x"fffb2781",
			2506 => x"001b2781",
			2507 => x"0e008604",
			2508 => x"00072781",
			2509 => x"ff502781",
			2510 => x"003c2781",
			2511 => x"0a00431c",
			2512 => x"0d00200c",
			2513 => x"00014c08",
			2514 => x"07003704",
			2515 => x"001b2781",
			2516 => x"00d02781",
			2517 => x"ffed2781",
			2518 => x"09002b08",
			2519 => x"05003804",
			2520 => x"ffab2781",
			2521 => x"00292781",
			2522 => x"00012804",
			2523 => x"00002781",
			2524 => x"004d2781",
			2525 => x"03004504",
			2526 => x"00032781",
			2527 => x"ffb32781",
			2528 => x"08002640",
			2529 => x"02011c30",
			2530 => x"07002904",
			2531 => x"fef2284d",
			2532 => x"09002518",
			2533 => x"01000e0c",
			2534 => x"0a002d08",
			2535 => x"03002704",
			2536 => x"ffaf284d",
			2537 => x"0076284d",
			2538 => x"ff10284d",
			2539 => x"09002108",
			2540 => x"0a002d04",
			2541 => x"00c0284d",
			2542 => x"ff7a284d",
			2543 => x"0162284d",
			2544 => x"0a003108",
			2545 => x"03001a04",
			2546 => x"ffe0284d",
			2547 => x"00e3284d",
			2548 => x"09002704",
			2549 => x"fee3284d",
			2550 => x"09002904",
			2551 => x"0056284d",
			2552 => x"ffda284d",
			2553 => x"0b001b0c",
			2554 => x"05003904",
			2555 => x"fe8f284d",
			2556 => x"0a003b04",
			2557 => x"00a3284d",
			2558 => x"ff0c284d",
			2559 => x"0023284d",
			2560 => x"0201371c",
			2561 => x"0c00220c",
			2562 => x"06009c04",
			2563 => x"ffd7284d",
			2564 => x"0e009d04",
			2565 => x"0179284d",
			2566 => x"000a284d",
			2567 => x"01001708",
			2568 => x"07004004",
			2569 => x"fed0284d",
			2570 => x"0010284d",
			2571 => x"00010c04",
			2572 => x"ffca284d",
			2573 => x"00c2284d",
			2574 => x"03002e04",
			2575 => x"ff2b284d",
			2576 => x"0a003d04",
			2577 => x"010a284d",
			2578 => x"000a284d",
			2579 => x"01000e08",
			2580 => x"08002304",
			2581 => x"fe8a28d9",
			2582 => x"00af28d9",
			2583 => x"07004438",
			2584 => x"02013728",
			2585 => x"0c002214",
			2586 => x"0800270c",
			2587 => x"01001808",
			2588 => x"05002404",
			2589 => x"016928d9",
			2590 => x"002128d9",
			2591 => x"fefe28d9",
			2592 => x"0e009804",
			2593 => x"017428d9",
			2594 => x"006a28d9",
			2595 => x"0100170c",
			2596 => x"07004008",
			2597 => x"09002a04",
			2598 => x"ffe628d9",
			2599 => x"fe6d28d9",
			2600 => x"fffd28d9",
			2601 => x"0c002704",
			2602 => x"00e528d9",
			2603 => x"ffcb28d9",
			2604 => x"0e00a40c",
			2605 => x"02014108",
			2606 => x"0a003604",
			2607 => x"fe7228d9",
			2608 => x"ff8e28d9",
			2609 => x"003628d9",
			2610 => x"00b728d9",
			2611 => x"00011e04",
			2612 => x"ffdf28d9",
			2613 => x"015a28d9",
			2614 => x"07004040",
			2615 => x"01000e08",
			2616 => x"08002304",
			2617 => x"fef0297d",
			2618 => x"0040297d",
			2619 => x"0600a418",
			2620 => x"0f00b514",
			2621 => x"0f00ae10",
			2622 => x"0f008208",
			2623 => x"0d001904",
			2624 => x"ff22297d",
			2625 => x"003c297d",
			2626 => x"06008004",
			2627 => x"0028297d",
			2628 => x"00ec297d",
			2629 => x"ff45297d",
			2630 => x"00ff297d",
			2631 => x"07003708",
			2632 => x"0d001804",
			2633 => x"ffe7297d",
			2634 => x"fed0297d",
			2635 => x"0d001d0c",
			2636 => x"00014308",
			2637 => x"0f00c404",
			2638 => x"0042297d",
			2639 => x"0149297d",
			2640 => x"ff72297d",
			2641 => x"0f00cd08",
			2642 => x"0f00c304",
			2643 => x"fff3297d",
			2644 => x"fef7297d",
			2645 => x"0026297d",
			2646 => x"0c002104",
			2647 => x"011b297d",
			2648 => x"0d002108",
			2649 => x"03003304",
			2650 => x"ff7c297d",
			2651 => x"001a297d",
			2652 => x"02010a04",
			2653 => x"ffec297d",
			2654 => x"00a1297d",
			2655 => x"08001f10",
			2656 => x"01000e04",
			2657 => x"feb42a19",
			2658 => x"09001e04",
			2659 => x"ff4e2a19",
			2660 => x"09002004",
			2661 => x"00392a19",
			2662 => x"ff932a19",
			2663 => x"0a002a08",
			2664 => x"06006504",
			2665 => x"ff572a19",
			2666 => x"01192a19",
			2667 => x"0900210c",
			2668 => x"01001008",
			2669 => x"0d001704",
			2670 => x"ff072a19",
			2671 => x"008d2a19",
			2672 => x"fec42a19",
			2673 => x"04002110",
			2674 => x"04001f0c",
			2675 => x"0a003108",
			2676 => x"04001a04",
			2677 => x"ffad2a19",
			2678 => x"016c2a19",
			2679 => x"ff4f2a19",
			2680 => x"fefe2a19",
			2681 => x"0a003b10",
			2682 => x"0c001e08",
			2683 => x"02013904",
			2684 => x"01292a19",
			2685 => x"002f2a19",
			2686 => x"09002804",
			2687 => x"fef02a19",
			2688 => x"00a42a19",
			2689 => x"0e009908",
			2690 => x"01001704",
			2691 => x"ff1f2a19",
			2692 => x"008c2a19",
			2693 => x"01132a19",
			2694 => x"0d001714",
			2695 => x"08001f04",
			2696 => x"fe642aad",
			2697 => x"05002408",
			2698 => x"01000c04",
			2699 => x"fefb2aad",
			2700 => x"01cd2aad",
			2701 => x"04002804",
			2702 => x"fe5f2aad",
			2703 => x"ff072aad",
			2704 => x"0f006504",
			2705 => x"fe6e2aad",
			2706 => x"0300412c",
			2707 => x"0500391c",
			2708 => x"0a00310c",
			2709 => x"09001e04",
			2710 => x"fe7a2aad",
			2711 => x"06009704",
			2712 => x"02322aad",
			2713 => x"00ea2aad",
			2714 => x"08002608",
			2715 => x"00012404",
			2716 => x"00ae2aad",
			2717 => x"fe3c2aad",
			2718 => x"00014304",
			2719 => x"012d2aad",
			2720 => x"ff532aad",
			2721 => x"08002004",
			2722 => x"fe972aad",
			2723 => x"07003b08",
			2724 => x"03003404",
			2725 => x"017c2aad",
			2726 => x"fff22aad",
			2727 => x"01ac2aad",
			2728 => x"0d002104",
			2729 => x"fe592aad",
			2730 => x"ff6b2aad",
			2731 => x"08002320",
			2732 => x"01000e04",
			2733 => x"fe602b41",
			2734 => x"0f006c04",
			2735 => x"fe672b41",
			2736 => x"0f00bb10",
			2737 => x"0c001704",
			2738 => x"ff562b41",
			2739 => x"03003404",
			2740 => x"025b2b41",
			2741 => x"08002204",
			2742 => x"fe6b2b41",
			2743 => x"ff8f2b41",
			2744 => x"0600c404",
			2745 => x"fe302b41",
			2746 => x"00e22b41",
			2747 => x"0f007504",
			2748 => x"fe672b41",
			2749 => x"03004624",
			2750 => x"05003814",
			2751 => x"03002704",
			2752 => x"01cc2b41",
			2753 => x"02012708",
			2754 => x"08002704",
			2755 => x"00642b41",
			2756 => x"01c72b41",
			2757 => x"03002e04",
			2758 => x"fea02b41",
			2759 => x"00c12b41",
			2760 => x"07003b08",
			2761 => x"09002604",
			2762 => x"00492b41",
			2763 => x"01b72b41",
			2764 => x"0c001e04",
			2765 => x"02232b41",
			2766 => x"01b42b41",
			2767 => x"fe322b41",
			2768 => x"0e009448",
			2769 => x"0001313c",
			2770 => x"0e009134",
			2771 => x"01001420",
			2772 => x"04002110",
			2773 => x"04001d08",
			2774 => x"01001004",
			2775 => x"ff732c1d",
			2776 => x"00132c1d",
			2777 => x"01000e04",
			2778 => x"ffdf2c1d",
			2779 => x"00fa2c1d",
			2780 => x"03002d08",
			2781 => x"05003304",
			2782 => x"ff782c1d",
			2783 => x"007f2c1d",
			2784 => x"08002304",
			2785 => x"ffc62c1d",
			2786 => x"ff0d2c1d",
			2787 => x"0200fd10",
			2788 => x"0a003408",
			2789 => x"0d001f04",
			2790 => x"ff612c1d",
			2791 => x"00122c1d",
			2792 => x"0f006504",
			2793 => x"ffd72c1d",
			2794 => x"00552c1d",
			2795 => x"01352c1d",
			2796 => x"05003804",
			2797 => x"ff092c1d",
			2798 => x"002b2c1d",
			2799 => x"09002608",
			2800 => x"04002904",
			2801 => x"feb82c1d",
			2802 => x"fffe2c1d",
			2803 => x"004c2c1d",
			2804 => x"03002e18",
			2805 => x"0a002f08",
			2806 => x"04001804",
			2807 => x"ffe32c1d",
			2808 => x"00e82c1d",
			2809 => x"02013308",
			2810 => x"01001204",
			2811 => x"ffef2c1d",
			2812 => x"00c02c1d",
			2813 => x"0f00dc04",
			2814 => x"fef32c1d",
			2815 => x"ffd82c1d",
			2816 => x"0a003b08",
			2817 => x"0b001804",
			2818 => x"ffb52c1d",
			2819 => x"01262c1d",
			2820 => x"04002c04",
			2821 => x"ff4c2c1d",
			2822 => x"00912c1d",
			2823 => x"0d001920",
			2824 => x"07002a04",
			2825 => x"ff3d2cc9",
			2826 => x"0200e910",
			2827 => x"0b001404",
			2828 => x"ffc92cc9",
			2829 => x"05003908",
			2830 => x"01000c04",
			2831 => x"ffed2cc9",
			2832 => x"00d02cc9",
			2833 => x"ffcd2cc9",
			2834 => x"03003304",
			2835 => x"ff412cc9",
			2836 => x"0c001a04",
			2837 => x"005b2cc9",
			2838 => x"ffb02cc9",
			2839 => x"03004534",
			2840 => x"0500392c",
			2841 => x"01001410",
			2842 => x"0a00340c",
			2843 => x"0b001c08",
			2844 => x"08002004",
			2845 => x"ffd42cc9",
			2846 => x"00c02cc9",
			2847 => x"ffa62cc9",
			2848 => x"ff232cc9",
			2849 => x"04002110",
			2850 => x"04001d08",
			2851 => x"0c002604",
			2852 => x"00aa2cc9",
			2853 => x"ffe62cc9",
			2854 => x"0e009304",
			2855 => x"ff622cc9",
			2856 => x"ffe72cc9",
			2857 => x"02013708",
			2858 => x"0a003204",
			2859 => x"001b2cc9",
			2860 => x"01332cc9",
			2861 => x"ffc62cc9",
			2862 => x"01001204",
			2863 => x"fffd2cc9",
			2864 => x"01042cc9",
			2865 => x"ff582cc9",
			2866 => x"0d001f64",
			2867 => x"05003438",
			2868 => x"0000c714",
			2869 => x"0200b00c",
			2870 => x"0d001704",
			2871 => x"ff3a2dd5",
			2872 => x"0e004304",
			2873 => x"ffba2dd5",
			2874 => x"00a72dd5",
			2875 => x"0b001704",
			2876 => x"01002dd5",
			2877 => x"fff82dd5",
			2878 => x"0e009410",
			2879 => x"0201210c",
			2880 => x"00012808",
			2881 => x"03002904",
			2882 => x"ff042dd5",
			2883 => x"ffd22dd5",
			2884 => x"00f02dd5",
			2885 => x"fea42dd5",
			2886 => x"0a002f08",
			2887 => x"0f00e004",
			2888 => x"00ee2dd5",
			2889 => x"ffd32dd5",
			2890 => x"02013308",
			2891 => x"00012804",
			2892 => x"ffdd2dd5",
			2893 => x"00922dd5",
			2894 => x"fefe2dd5",
			2895 => x"0d001b1c",
			2896 => x"0c001b10",
			2897 => x"0700330c",
			2898 => x"03002e08",
			2899 => x"07002a04",
			2900 => x"ffb62dd5",
			2901 => x"00942dd5",
			2902 => x"ff112dd5",
			2903 => x"00e52dd5",
			2904 => x"0c001d04",
			2905 => x"fee32dd5",
			2906 => x"0c001e04",
			2907 => x"005a2dd5",
			2908 => x"ff782dd5",
			2909 => x"0001430c",
			2910 => x"03004408",
			2911 => x"07003604",
			2912 => x"00672dd5",
			2913 => x"01532dd5",
			2914 => x"ff6b2dd5",
			2915 => x"ff662dd5",
			2916 => x"04002b10",
			2917 => x"08002d08",
			2918 => x"0000f404",
			2919 => x"ffd02dd5",
			2920 => x"015d2dd5",
			2921 => x"05003604",
			2922 => x"00752dd5",
			2923 => x"ff552dd5",
			2924 => x"0d002004",
			2925 => x"00c42dd5",
			2926 => x"01001708",
			2927 => x"08002704",
			2928 => x"00182dd5",
			2929 => x"feeb2dd5",
			2930 => x"00011604",
			2931 => x"ffee2dd5",
			2932 => x"007c2dd5",
			2933 => x"08002750",
			2934 => x"0f00c138",
			2935 => x"0600a934",
			2936 => x"03002d1c",
			2937 => x"09001e0c",
			2938 => x"05002208",
			2939 => x"0a002704",
			2940 => x"ffe92eb9",
			2941 => x"003c2eb9",
			2942 => x"ff8c2eb9",
			2943 => x"09002508",
			2944 => x"06006504",
			2945 => x"ffd62eb9",
			2946 => x"00b12eb9",
			2947 => x"0d001d04",
			2948 => x"ffb42eb9",
			2949 => x"001c2eb9",
			2950 => x"0400260c",
			2951 => x"0f00b908",
			2952 => x"0d001a04",
			2953 => x"00052eb9",
			2954 => x"ff8e2eb9",
			2955 => x"007d2eb9",
			2956 => x"08002608",
			2957 => x"07003a04",
			2958 => x"ff4b2eb9",
			2959 => x"00102eb9",
			2960 => x"00442eb9",
			2961 => x"00872eb9",
			2962 => x"0a00360c",
			2963 => x"04001b08",
			2964 => x"04001a04",
			2965 => x"ffe72eb9",
			2966 => x"00212eb9",
			2967 => x"ff342eb9",
			2968 => x"07003b08",
			2969 => x"03003104",
			2970 => x"00372eb9",
			2971 => x"ff9a2eb9",
			2972 => x"00562eb9",
			2973 => x"0e008a0c",
			2974 => x"0a003104",
			2975 => x"ffae2eb9",
			2976 => x"06009504",
			2977 => x"ffec2eb9",
			2978 => x"00432eb9",
			2979 => x"02013708",
			2980 => x"0600bd04",
			2981 => x"00ec2eb9",
			2982 => x"fff72eb9",
			2983 => x"02013c04",
			2984 => x"ffc82eb9",
			2985 => x"0600c204",
			2986 => x"00772eb9",
			2987 => x"0f00e204",
			2988 => x"ffee2eb9",
			2989 => x"00002eb9",
			2990 => x"0700405c",
			2991 => x"05003a40",
			2992 => x"0a003120",
			2993 => x"04002010",
			2994 => x"09001e04",
			2995 => x"ff9f2f7d",
			2996 => x"04001804",
			2997 => x"ffdc2f7d",
			2998 => x"06007004",
			2999 => x"fff62f7d",
			3000 => x"00bd2f7d",
			3001 => x"07002c08",
			3002 => x"09001d04",
			3003 => x"ffe42f7d",
			3004 => x"005a2f7d",
			3005 => x"04002304",
			3006 => x"ff6c2f7d",
			3007 => x"00122f7d",
			3008 => x"02011a10",
			3009 => x"05003204",
			3010 => x"ffa42f7d",
			3011 => x"03002f04",
			3012 => x"00822f7d",
			3013 => x"0d001904",
			3014 => x"00112f7d",
			3015 => x"ffbc2f7d",
			3016 => x"0800260c",
			3017 => x"0b001808",
			3018 => x"05003604",
			3019 => x"ffdf2f7d",
			3020 => x"00122f7d",
			3021 => x"ff322f7d",
			3022 => x"ffeb2f7d",
			3023 => x"03003508",
			3024 => x"08002004",
			3025 => x"ffef2f7d",
			3026 => x"009f2f7d",
			3027 => x"0100160c",
			3028 => x"07003e08",
			3029 => x"0a003904",
			3030 => x"00042f7d",
			3031 => x"ff942f7d",
			3032 => x"000a2f7d",
			3033 => x"03003a04",
			3034 => x"00342f7d",
			3035 => x"ffe22f7d",
			3036 => x"0600a304",
			3037 => x"ffec2f7d",
			3038 => x"008e2f7d",
			3039 => x"0700404c",
			3040 => x"0f00ae20",
			3041 => x"07002904",
			3042 => x"ff063039",
			3043 => x"0d001504",
			3044 => x"ff7a3039",
			3045 => x"04003610",
			3046 => x"04001e08",
			3047 => x"0000c704",
			3048 => x"006c3039",
			3049 => x"ff9b3039",
			3050 => x"06005e04",
			3051 => x"fff23039",
			3052 => x"01313039",
			3053 => x"06008b04",
			3054 => x"ff8d3039",
			3055 => x"000b3039",
			3056 => x"07003304",
			3057 => x"fedc3039",
			3058 => x"04002110",
			3059 => x"0400200c",
			3060 => x"0a003108",
			3061 => x"04001804",
			3062 => x"ffd23039",
			3063 => x"01283039",
			3064 => x"ff893039",
			3065 => x"febb3039",
			3066 => x"04002608",
			3067 => x"02013704",
			3068 => x"012e3039",
			3069 => x"fff53039",
			3070 => x"08002608",
			3071 => x"05003904",
			3072 => x"feeb3039",
			3073 => x"00213039",
			3074 => x"0d002004",
			3075 => x"01183039",
			3076 => x"ff683039",
			3077 => x"0c002104",
			3078 => x"01383039",
			3079 => x"0d002108",
			3080 => x"05004104",
			3081 => x"ff783039",
			3082 => x"00113039",
			3083 => x"02010a04",
			3084 => x"ffd33039",
			3085 => x"00c43039",
			3086 => x"08002328",
			3087 => x"03003320",
			3088 => x"0600901c",
			3089 => x"06008014",
			3090 => x"0500360c",
			3091 => x"02009008",
			3092 => x"00009204",
			3093 => x"ffec311d",
			3094 => x"0013311d",
			3095 => x"ffb7311d",
			3096 => x"0000aa04",
			3097 => x"fff2311d",
			3098 => x"0015311d",
			3099 => x"03002404",
			3100 => x"fff7311d",
			3101 => x"004c311d",
			3102 => x"ff6f311d",
			3103 => x"0a003704",
			3104 => x"0045311d",
			3105 => x"ffdb311d",
			3106 => x"0201373c",
			3107 => x"03003124",
			3108 => x"00012614",
			3109 => x"09002508",
			3110 => x"0f006504",
			3111 => x"fff9311d",
			3112 => x"0050311d",
			3113 => x"08002704",
			3114 => x"ff9f311d",
			3115 => x"0e007304",
			3116 => x"fff0311d",
			3117 => x"001e311d",
			3118 => x"0c001e04",
			3119 => x"00ad311d",
			3120 => x"0600b604",
			3121 => x"ffd6311d",
			3122 => x"0600bc04",
			3123 => x"0055311d",
			3124 => x"fff9311d",
			3125 => x"05003804",
			3126 => x"ffb3311d",
			3127 => x"0600a80c",
			3128 => x"07003504",
			3129 => x"0013311d",
			3130 => x"01001504",
			3131 => x"ffb7311d",
			3132 => x"0003311d",
			3133 => x"04003504",
			3134 => x"005c311d",
			3135 => x"ffff311d",
			3136 => x"0b00210c",
			3137 => x"03002e04",
			3138 => x"ff80311d",
			3139 => x"0600bc04",
			3140 => x"ffd4311d",
			3141 => x"0042311d",
			3142 => x"003f311d",
			3143 => x"07004050",
			3144 => x"01000e08",
			3145 => x"08002304",
			3146 => x"feba31e1",
			3147 => x"008f31e1",
			3148 => x"0f00ae20",
			3149 => x"0600801c",
			3150 => x"0d001910",
			3151 => x"08001d08",
			3152 => x"08001c04",
			3153 => x"ffe631e1",
			3154 => x"008031e1",
			3155 => x"03001f04",
			3156 => x"003831e1",
			3157 => x"fed831e1",
			3158 => x"06005e04",
			3159 => x"ff6031e1",
			3160 => x"0200ce04",
			3161 => x"011331e1",
			3162 => x"ffac31e1",
			3163 => x"013531e1",
			3164 => x"05003818",
			3165 => x"0400200c",
			3166 => x"0a003108",
			3167 => x"05002804",
			3168 => x"ff3d31e1",
			3169 => x"012e31e1",
			3170 => x"ff8931e1",
			3171 => x"08002608",
			3172 => x"0b001804",
			3173 => x"002b31e1",
			3174 => x"fee031e1",
			3175 => x"ffd431e1",
			3176 => x"03003508",
			3177 => x"08002404",
			3178 => x"000631e1",
			3179 => x"013f31e1",
			3180 => x"0e009204",
			3181 => x"ff5931e1",
			3182 => x"003e31e1",
			3183 => x"0c002104",
			3184 => x"014e31e1",
			3185 => x"0d002108",
			3186 => x"03003304",
			3187 => x"ff5731e1",
			3188 => x"002231e1",
			3189 => x"00011404",
			3190 => x"ffcf31e1",
			3191 => x"00d531e1",
			3192 => x"0d001708",
			3193 => x"08002204",
			3194 => x"fe6b327d",
			3195 => x"ffa0327d",
			3196 => x"03004544",
			3197 => x"0500392c",
			3198 => x"02012110",
			3199 => x"0f006504",
			3200 => x"fe8e327d",
			3201 => x"0e009108",
			3202 => x"0d001c04",
			3203 => x"0085327d",
			3204 => x"01c7327d",
			3205 => x"ff2b327d",
			3206 => x"08002610",
			3207 => x"00014208",
			3208 => x"03002d04",
			3209 => x"fe05327d",
			3210 => x"fea5327d",
			3211 => x"01001204",
			3212 => x"febb327d",
			3213 => x"004c327d",
			3214 => x"05003304",
			3215 => x"012d327d",
			3216 => x"03002e04",
			3217 => x"fee4327d",
			3218 => x"00bd327d",
			3219 => x"0f00b80c",
			3220 => x"08002408",
			3221 => x"03003804",
			3222 => x"ff27327d",
			3223 => x"fe2f327d",
			3224 => x"015e327d",
			3225 => x"00013f04",
			3226 => x"01aa327d",
			3227 => x"0f00d304",
			3228 => x"ff73327d",
			3229 => x"017f327d",
			3230 => x"fe75327d",
			3231 => x"07003f54",
			3232 => x"0201374c",
			3233 => x"03002f28",
			3234 => x"03002a14",
			3235 => x"01001610",
			3236 => x"0c001708",
			3237 => x"05002404",
			3238 => x"003b3349",
			3239 => x"ff883349",
			3240 => x"06006504",
			3241 => x"ffd23349",
			3242 => x"00a23349",
			3243 => x"ff5b3349",
			3244 => x"07003510",
			3245 => x"06008d08",
			3246 => x"02009204",
			3247 => x"ffd73349",
			3248 => x"00613349",
			3249 => x"04002004",
			3250 => x"00293349",
			3251 => x"ff6e3349",
			3252 => x"00c93349",
			3253 => x"08002414",
			3254 => x"0b001708",
			3255 => x"02011604",
			3256 => x"ffcb3349",
			3257 => x"003a3349",
			3258 => x"0d001c04",
			3259 => x"ff203349",
			3260 => x"0d001d04",
			3261 => x"00053349",
			3262 => x"fffa3349",
			3263 => x"07003d0c",
			3264 => x"03004508",
			3265 => x"0e007f04",
			3266 => x"ffcb3349",
			3267 => x"00a73349",
			3268 => x"ffb63349",
			3269 => x"ff8b3349",
			3270 => x"00015504",
			3271 => x"ff403349",
			3272 => x"000c3349",
			3273 => x"03005310",
			3274 => x"01001a04",
			3275 => x"00c63349",
			3276 => x"0e00a108",
			3277 => x"01001d04",
			3278 => x"ffd33349",
			3279 => x"00093349",
			3280 => x"002d3349",
			3281 => x"ffe13349",
			3282 => x"01000e08",
			3283 => x"08002304",
			3284 => x"fe6a33e7",
			3285 => x"005633e7",
			3286 => x"09001e04",
			3287 => x"fe7633e7",
			3288 => x"02012524",
			3289 => x"0f006504",
			3290 => x"fe8c33e7",
			3291 => x"0a003710",
			3292 => x"09002508",
			3293 => x"04002304",
			3294 => x"01ad33e7",
			3295 => x"013733e7",
			3296 => x"00012704",
			3297 => x"ff6333e7",
			3298 => x"01ab33e7",
			3299 => x"08002408",
			3300 => x"07003c04",
			3301 => x"fe2833e7",
			3302 => x"ffc633e7",
			3303 => x"0e007f04",
			3304 => x"ff4e33e7",
			3305 => x"016b33e7",
			3306 => x"07003f14",
			3307 => x"0800260c",
			3308 => x"03002d04",
			3309 => x"fdfb33e7",
			3310 => x"0d001b04",
			3311 => x"fea833e7",
			3312 => x"002133e7",
			3313 => x"0a003904",
			3314 => x"007933e7",
			3315 => x"ff3433e7",
			3316 => x"03002e08",
			3317 => x"07004504",
			3318 => x"ff5f33e7",
			3319 => x"017533e7",
			3320 => x"019f33e7",
			3321 => x"0100121c",
			3322 => x"08002210",
			3323 => x"01000e04",
			3324 => x"fe563459",
			3325 => x"0b001708",
			3326 => x"09001d04",
			3327 => x"fe583459",
			3328 => x"01073459",
			3329 => x"fe573459",
			3330 => x"0b001b08",
			3331 => x"0f00bd04",
			3332 => x"01973459",
			3333 => x"ffa63459",
			3334 => x"fe593459",
			3335 => x"0f006504",
			3336 => x"fe553459",
			3337 => x"0a004a18",
			3338 => x"0d001904",
			3339 => x"ffad3459",
			3340 => x"0500390c",
			3341 => x"00011f04",
			3342 => x"02953459",
			3343 => x"07004004",
			3344 => x"00533459",
			3345 => x"01cc3459",
			3346 => x"0c001c04",
			3347 => x"01913459",
			3348 => x"02053459",
			3349 => x"fe113459",
			3350 => x"08002428",
			3351 => x"0a002d10",
			3352 => x"09001d04",
			3353 => x"ffcd3515",
			3354 => x"0f00aa08",
			3355 => x"06006504",
			3356 => x"ffe53515",
			3357 => x"00793515",
			3358 => x"ffe53515",
			3359 => x"0e00960c",
			3360 => x"0b001508",
			3361 => x"03002a04",
			3362 => x"00133515",
			3363 => x"fff93515",
			3364 => x"ff843515",
			3365 => x"02013104",
			3366 => x"ffd73515",
			3367 => x"0d001804",
			3368 => x"fff33515",
			3369 => x"00463515",
			3370 => x"03002e14",
			3371 => x"03002708",
			3372 => x"00007204",
			3373 => x"fff63515",
			3374 => x"00633515",
			3375 => x"02011d04",
			3376 => x"00413515",
			3377 => x"07004404",
			3378 => x"ff673515",
			3379 => x"00293515",
			3380 => x"0a003e14",
			3381 => x"00012508",
			3382 => x"00011f04",
			3383 => x"00193515",
			3384 => x"ffbc3515",
			3385 => x"0c002204",
			3386 => x"00b63515",
			3387 => x"0d002204",
			3388 => x"ffe13515",
			3389 => x"00243515",
			3390 => x"01001708",
			3391 => x"07004004",
			3392 => x"ffb73515",
			3393 => x"00053515",
			3394 => x"00011604",
			3395 => x"fffb3515",
			3396 => x"00103515",
			3397 => x"01001434",
			3398 => x"01001224",
			3399 => x"01000e08",
			3400 => x"08002304",
			3401 => x"fe3735b9",
			3402 => x"feba35b9",
			3403 => x"0f008c0c",
			3404 => x"0c001908",
			3405 => x"05002a04",
			3406 => x"fe3e35b9",
			3407 => x"003135b9",
			3408 => x"fe3635b9",
			3409 => x"08002208",
			3410 => x"00010a04",
			3411 => x"008635b9",
			3412 => x"fe3235b9",
			3413 => x"0f00c204",
			3414 => x"03f235b9",
			3415 => x"fff335b9",
			3416 => x"0f008208",
			3417 => x"06006504",
			3418 => x"fe3935b9",
			3419 => x"ff3d35b9",
			3420 => x"05003804",
			3421 => x"006735b9",
			3422 => x"037135b9",
			3423 => x"0f009308",
			3424 => x"0c002404",
			3425 => x"ff2b35b9",
			3426 => x"fe3835b9",
			3427 => x"09002404",
			3428 => x"010c35b9",
			3429 => x"03002a08",
			3430 => x"07003e04",
			3431 => x"01f635b9",
			3432 => x"048635b9",
			3433 => x"0f00c204",
			3434 => x"047235b9",
			3435 => x"0f00c404",
			3436 => x"037935b9",
			3437 => x"044835b9",
			3438 => x"0d001910",
			3439 => x"05002208",
			3440 => x"0a002704",
			3441 => x"ffe9365d",
			3442 => x"002a365d",
			3443 => x"0e00a504",
			3444 => x"ff8f365d",
			3445 => x"0006365d",
			3446 => x"0900251c",
			3447 => x"0400200c",
			3448 => x"0b001c08",
			3449 => x"04001804",
			3450 => x"fffc365d",
			3451 => x"009c365d",
			3452 => x"fff4365d",
			3453 => x"04002508",
			3454 => x"0f00c204",
			3455 => x"fffb365d",
			3456 => x"ffa6365d",
			3457 => x"0600a704",
			3458 => x"ffe9365d",
			3459 => x"007f365d",
			3460 => x"0500381c",
			3461 => x"09002b14",
			3462 => x"0500330c",
			3463 => x"03002908",
			3464 => x"04001a04",
			3465 => x"0014365d",
			3466 => x"ff91365d",
			3467 => x"0072365d",
			3468 => x"01001904",
			3469 => x"ff3e365d",
			3470 => x"0031365d",
			3471 => x"00012804",
			3472 => x"ffea365d",
			3473 => x"0063365d",
			3474 => x"03004608",
			3475 => x"05003904",
			3476 => x"0004365d",
			3477 => x"008a365d",
			3478 => x"ffae365d",
			3479 => x"0f00bf24",
			3480 => x"0f006c0c",
			3481 => x"0000a204",
			3482 => x"ffab3721",
			3483 => x"0000a604",
			3484 => x"00143721",
			3485 => x"ffeb3721",
			3486 => x"09001e08",
			3487 => x"0000b804",
			3488 => x"00243721",
			3489 => x"ffb23721",
			3490 => x"0d001708",
			3491 => x"09002304",
			3492 => x"ffcc3721",
			3493 => x"00043721",
			3494 => x"05005304",
			3495 => x"008f3721",
			3496 => x"ffd33721",
			3497 => x"0e009414",
			3498 => x"07003a0c",
			3499 => x"0b001808",
			3500 => x"0b001704",
			3501 => x"fff13721",
			3502 => x"00133721",
			3503 => x"ff6d3721",
			3504 => x"05003904",
			3505 => x"ffeb3721",
			3506 => x"00133721",
			3507 => x"03002e14",
			3508 => x"0a002f08",
			3509 => x"04001804",
			3510 => x"fff93721",
			3511 => x"005d3721",
			3512 => x"02013308",
			3513 => x"01001204",
			3514 => x"fffc3721",
			3515 => x"003e3721",
			3516 => x"ff6f3721",
			3517 => x"0a003b0c",
			3518 => x"0d001b08",
			3519 => x"00013a04",
			3520 => x"00023721",
			3521 => x"ffe13721",
			3522 => x"00a33721",
			3523 => x"04002c04",
			3524 => x"ffc13721",
			3525 => x"00014904",
			3526 => x"00163721",
			3527 => x"00003721",
			3528 => x"01001224",
			3529 => x"08002214",
			3530 => x"01000e04",
			3531 => x"fe5c37ad",
			3532 => x"0b001508",
			3533 => x"0d001504",
			3534 => x"fe6a37ad",
			3535 => x"019637ad",
			3536 => x"0b001704",
			3537 => x"ff3c37ad",
			3538 => x"fe6037ad",
			3539 => x"0c001d0c",
			3540 => x"07002c04",
			3541 => x"fe6c37ad",
			3542 => x"0f00be04",
			3543 => x"01c637ad",
			3544 => x"002837ad",
			3545 => x"fe6137ad",
			3546 => x"06005e04",
			3547 => x"fe5e37ad",
			3548 => x"0300461c",
			3549 => x"0d001904",
			3550 => x"ff8e37ad",
			3551 => x"0201370c",
			3552 => x"0e007d04",
			3553 => x"02b037ad",
			3554 => x"07003704",
			3555 => x"005937ad",
			3556 => x"01bd37ad",
			3557 => x"0e009904",
			3558 => x"fe0637ad",
			3559 => x"03002e04",
			3560 => x"ffba37ad",
			3561 => x"01ea37ad",
			3562 => x"fdfc37ad",
			3563 => x"0900211c",
			3564 => x"0200ca10",
			3565 => x"0200ae04",
			3566 => x"ffa23859",
			3567 => x"0e006204",
			3568 => x"fff73859",
			3569 => x"03002404",
			3570 => x"00033859",
			3571 => x"007c3859",
			3572 => x"05003a04",
			3573 => x"ff5f3859",
			3574 => x"05003e04",
			3575 => x"001b3859",
			3576 => x"fffa3859",
			3577 => x"04002110",
			3578 => x"0400200c",
			3579 => x"0a003108",
			3580 => x"05002804",
			3581 => x"ffce3859",
			3582 => x"00bd3859",
			3583 => x"ff9b3859",
			3584 => x"ff6f3859",
			3585 => x"0a003b18",
			3586 => x"02013710",
			3587 => x"08002304",
			3588 => x"ffea3859",
			3589 => x"0d001e04",
			3590 => x"00cc3859",
			3591 => x"0b001f04",
			3592 => x"ffd93859",
			3593 => x"00673859",
			3594 => x"03002e04",
			3595 => x"ff823859",
			3596 => x"00663859",
			3597 => x"0600b710",
			3598 => x"0001390c",
			3599 => x"0d001b04",
			3600 => x"ffaa3859",
			3601 => x"04003e04",
			3602 => x"00673859",
			3603 => x"ffcf3859",
			3604 => x"ff7b3859",
			3605 => x"00323859",
			3606 => x"0d001714",
			3607 => x"08001f04",
			3608 => x"fe6b38e5",
			3609 => x"05002408",
			3610 => x"0e002f04",
			3611 => x"ff5638e5",
			3612 => x"015838e5",
			3613 => x"04002804",
			3614 => x"fe7338e5",
			3615 => x"ff2138e5",
			3616 => x"03004530",
			3617 => x"05003914",
			3618 => x"04002910",
			3619 => x"0700420c",
			3620 => x"0e009b08",
			3621 => x"0e009404",
			3622 => x"fff838e5",
			3623 => x"012e38e5",
			3624 => x"feb038e5",
			3625 => x"019138e5",
			3626 => x"fede38e5",
			3627 => x"0f00b80c",
			3628 => x"08002408",
			3629 => x"0b001a04",
			3630 => x"ff2a38e5",
			3631 => x"fdf338e5",
			3632 => x"015c38e5",
			3633 => x"02013a08",
			3634 => x"00013d04",
			3635 => x"01b538e5",
			3636 => x"012038e5",
			3637 => x"0e00a404",
			3638 => x"ff4538e5",
			3639 => x"019838e5",
			3640 => x"fe6d38e5",
			3641 => x"0d001714",
			3642 => x"08001f04",
			3643 => x"fe663979",
			3644 => x"05002408",
			3645 => x"07002804",
			3646 => x"ff1b3979",
			3647 => x"01a23979",
			3648 => x"0c001904",
			3649 => x"fe613979",
			3650 => x"ff133979",
			3651 => x"07003f28",
			3652 => x"0f006504",
			3653 => x"fe743979",
			3654 => x"0000d308",
			3655 => x"04003c04",
			3656 => x"01df3979",
			3657 => x"fecd3979",
			3658 => x"08002610",
			3659 => x"04002008",
			3660 => x"03002904",
			3661 => x"ffa83979",
			3662 => x"01833979",
			3663 => x"0600af04",
			3664 => x"ff833979",
			3665 => x"fdea3979",
			3666 => x"04002104",
			3667 => x"ff453979",
			3668 => x"08002a04",
			3669 => x"016d3979",
			3670 => x"ff963979",
			3671 => x"05003508",
			3672 => x"07004404",
			3673 => x"ff753979",
			3674 => x"017c3979",
			3675 => x"03005304",
			3676 => x"01b13979",
			3677 => x"febe3979",
			3678 => x"08002744",
			3679 => x"0d001b2c",
			3680 => x"0c001a20",
			3681 => x"09002118",
			3682 => x"0200ca0c",
			3683 => x"07002904",
			3684 => x"ff653a3d",
			3685 => x"0b001404",
			3686 => x"ffa73a3d",
			3687 => x"00ce3a3d",
			3688 => x"05003a04",
			3689 => x"fedf3a3d",
			3690 => x"05003e04",
			3691 => x"003e3a3d",
			3692 => x"ffef3a3d",
			3693 => x"0a003704",
			3694 => x"00d53a3d",
			3695 => x"ffc73a3d",
			3696 => x"07003a08",
			3697 => x"09002304",
			3698 => x"fec73a3d",
			3699 => x"ff9e3a3d",
			3700 => x"fff73a3d",
			3701 => x"0001260c",
			3702 => x"0f00b008",
			3703 => x"06007e04",
			3704 => x"ffa83a3d",
			3705 => x"00ac3a3d",
			3706 => x"ff413a3d",
			3707 => x"02013908",
			3708 => x"00013804",
			3709 => x"011d3a3d",
			3710 => x"00793a3d",
			3711 => x"ff673a3d",
			3712 => x"02013718",
			3713 => x"0a003b0c",
			3714 => x"06008504",
			3715 => x"ffd63a3d",
			3716 => x"0600bc04",
			3717 => x"01443a3d",
			3718 => x"00163a3d",
			3719 => x"02012c08",
			3720 => x"06009604",
			3721 => x"ffdc3a3d",
			3722 => x"00843a3d",
			3723 => x"ff453a3d",
			3724 => x"03002e04",
			3725 => x"ff6a3a3d",
			3726 => x"00db3a3d",
			3727 => x"0d001710",
			3728 => x"09002308",
			3729 => x"08002204",
			3730 => x"fe713ae1",
			3731 => x"ff173ae1",
			3732 => x"08001d04",
			3733 => x"ff773ae1",
			3734 => x"00643ae1",
			3735 => x"08002728",
			3736 => x"07003e20",
			3737 => x"0e009018",
			3738 => x"07003a10",
			3739 => x"02011c08",
			3740 => x"09002504",
			3741 => x"00ae3ae1",
			3742 => x"fec43ae1",
			3743 => x"0d001a04",
			3744 => x"fe5e3ae1",
			3745 => x"ff703ae1",
			3746 => x"01001204",
			3747 => x"ff683ae1",
			3748 => x"01b53ae1",
			3749 => x"05003804",
			3750 => x"fdf23ae1",
			3751 => x"000e3ae1",
			3752 => x"03005304",
			3753 => x"01433ae1",
			3754 => x"ff7a3ae1",
			3755 => x"03002e14",
			3756 => x"02013710",
			3757 => x"0e008a08",
			3758 => x"08002904",
			3759 => x"ff563ae1",
			3760 => x"00933ae1",
			3761 => x"0600bb04",
			3762 => x"01b13ae1",
			3763 => x"ffc13ae1",
			3764 => x"ff563ae1",
			3765 => x"03004504",
			3766 => x"018e3ae1",
			3767 => x"fed03ae1",
			3768 => x"08002320",
			3769 => x"01000e04",
			3770 => x"fe5f3b6d",
			3771 => x"0f00bb14",
			3772 => x"0f00820c",
			3773 => x"0f006c04",
			3774 => x"fe653b6d",
			3775 => x"0f007404",
			3776 => x"016d3b6d",
			3777 => x"fe533b6d",
			3778 => x"0f00a904",
			3779 => x"01ba3b6d",
			3780 => x"ffb53b6d",
			3781 => x"00014c04",
			3782 => x"fe243b6d",
			3783 => x"ffc13b6d",
			3784 => x"0f006504",
			3785 => x"fe683b6d",
			3786 => x"03004620",
			3787 => x"05003810",
			3788 => x"04002004",
			3789 => x"01b83b6d",
			3790 => x"0d001b04",
			3791 => x"fee43b6d",
			3792 => x"0f00c204",
			3793 => x"01d23b6d",
			3794 => x"00113b6d",
			3795 => x"07003b08",
			3796 => x"03003304",
			3797 => x"01ab3b6d",
			3798 => x"00023b6d",
			3799 => x"08002604",
			3800 => x"02373b6d",
			3801 => x"01bb3b6d",
			3802 => x"fe4b3b6d",
			3803 => x"0d001f48",
			3804 => x"0201262c",
			3805 => x"0f00b820",
			3806 => x"0f00aa1c",
			3807 => x"0d001810",
			3808 => x"05002408",
			3809 => x"08001f04",
			3810 => x"ffea3c39",
			3811 => x"003a3c39",
			3812 => x"0e007704",
			3813 => x"ff933c39",
			3814 => x"00013c39",
			3815 => x"0f006504",
			3816 => x"ffca3c39",
			3817 => x"0c001e04",
			3818 => x"00b73c39",
			3819 => x"ffed3c39",
			3820 => x"ff653c39",
			3821 => x"05002e04",
			3822 => x"ffa53c39",
			3823 => x"04002704",
			3824 => x"00c23c39",
			3825 => x"fff33c39",
			3826 => x"04002710",
			3827 => x"0a002c08",
			3828 => x"05002804",
			3829 => x"fff03c39",
			3830 => x"004d3c39",
			3831 => x"05003804",
			3832 => x"ff373c39",
			3833 => x"fff63c39",
			3834 => x"03003508",
			3835 => x"0d001804",
			3836 => x"fff43c39",
			3837 => x"00883c39",
			3838 => x"ffd83c39",
			3839 => x"04002b10",
			3840 => x"08002d08",
			3841 => x"0000f404",
			3842 => x"ffec3c39",
			3843 => x"00cd3c39",
			3844 => x"0600bc04",
			3845 => x"ffbc3c39",
			3846 => x"00383c39",
			3847 => x"0d002004",
			3848 => x"00413c39",
			3849 => x"01001704",
			3850 => x"ff7d3c39",
			3851 => x"00011604",
			3852 => x"fffa3c39",
			3853 => x"00203c39",
			3854 => x"0e00943c",
			3855 => x"02012430",
			3856 => x"0e00912c",
			3857 => x"0f00b81c",
			3858 => x"0a002d0c",
			3859 => x"0e005b04",
			3860 => x"ffdf3ce5",
			3861 => x"0c001704",
			3862 => x"fff03ce5",
			3863 => x"00663ce5",
			3864 => x"0d001c08",
			3865 => x"07003b04",
			3866 => x"ff833ce5",
			3867 => x"00013ce5",
			3868 => x"0b002204",
			3869 => x"00343ce5",
			3870 => x"fff13ce5",
			3871 => x"04002608",
			3872 => x"09002104",
			3873 => x"fff53ce5",
			3874 => x"008d3ce5",
			3875 => x"03003304",
			3876 => x"ffd53ce5",
			3877 => x"001b3ce5",
			3878 => x"ffb03ce5",
			3879 => x"0b001808",
			3880 => x"0b001704",
			3881 => x"fff73ce5",
			3882 => x"000d3ce5",
			3883 => x"ff8d3ce5",
			3884 => x"01001710",
			3885 => x"05003808",
			3886 => x"0600b704",
			3887 => x"001f3ce5",
			3888 => x"ff9e3ce5",
			3889 => x"0600b704",
			3890 => x"fffc3ce5",
			3891 => x"004a3ce5",
			3892 => x"01001a04",
			3893 => x"00723ce5",
			3894 => x"09002b04",
			3895 => x"ffe63ce5",
			3896 => x"001b3ce5",
			3897 => x"01000c04",
			3898 => x"fe883d49",
			3899 => x"0a002808",
			3900 => x"06007104",
			3901 => x"fef83d49",
			3902 => x"01993d49",
			3903 => x"09001e04",
			3904 => x"fe973d49",
			3905 => x"0f00ae10",
			3906 => x"0f006504",
			3907 => x"feeb3d49",
			3908 => x"04003608",
			3909 => x"0c001f04",
			3910 => x"015e3d49",
			3911 => x"00693d49",
			3912 => x"ff003d49",
			3913 => x"07003308",
			3914 => x"05003004",
			3915 => x"ff833d49",
			3916 => x"fe703d49",
			3917 => x"03002904",
			3918 => x"ff4f3d49",
			3919 => x"0d001b04",
			3920 => x"ff863d49",
			3921 => x"00893d49",
			3922 => x"0d001714",
			3923 => x"08001f04",
			3924 => x"fe6a3df5",
			3925 => x"05002408",
			3926 => x"00006104",
			3927 => x"ff493df5",
			3928 => x"016e3df5",
			3929 => x"04002804",
			3930 => x"fe6e3df5",
			3931 => x"ff143df5",
			3932 => x"07003f34",
			3933 => x"0201372c",
			3934 => x"0c002218",
			3935 => x"08002710",
			3936 => x"03002f08",
			3937 => x"05002e04",
			3938 => x"ff5a3df5",
			3939 => x"011d3df5",
			3940 => x"08002404",
			3941 => x"fef33df5",
			3942 => x"00693df5",
			3943 => x"04002604",
			3944 => x"00923df5",
			3945 => x"019d3df5",
			3946 => x"0a003b08",
			3947 => x"04001b04",
			3948 => x"feb03df5",
			3949 => x"00bf3df5",
			3950 => x"07003c08",
			3951 => x"07003a04",
			3952 => x"fedf3df5",
			3953 => x"00013df5",
			3954 => x"fdd63df5",
			3955 => x"0600b704",
			3956 => x"fe663df5",
			3957 => x"ff7a3df5",
			3958 => x"05003508",
			3959 => x"0a003104",
			3960 => x"017d3df5",
			3961 => x"ff763df5",
			3962 => x"03005304",
			3963 => x"01a73df5",
			3964 => x"fee33df5",
			3965 => x"01001220",
			3966 => x"08002210",
			3967 => x"01000e04",
			3968 => x"fe583e91",
			3969 => x"0c001808",
			3970 => x"09001d04",
			3971 => x"fe5d3e91",
			3972 => x"00ee3e91",
			3973 => x"fe5a3e91",
			3974 => x"0c001d0c",
			3975 => x"07002c04",
			3976 => x"fe623e91",
			3977 => x"05003404",
			3978 => x"00863e91",
			3979 => x"02433e91",
			3980 => x"fe5b3e91",
			3981 => x"0f006504",
			3982 => x"fe593e91",
			3983 => x"0a004a28",
			3984 => x"0d001f14",
			3985 => x"0f00aa04",
			3986 => x"029e3e91",
			3987 => x"07003708",
			3988 => x"0f00bf04",
			3989 => x"ff5c3e91",
			3990 => x"fe193e91",
			3991 => x"03002a04",
			3992 => x"ffcd3e91",
			3993 => x"019c3e91",
			3994 => x"01001708",
			3995 => x"05003904",
			3996 => x"00b53e91",
			3997 => x"01ed3e91",
			3998 => x"03002e08",
			3999 => x"0c002204",
			4000 => x"015e3e91",
			4001 => x"01ec3e91",
			4002 => x"01f63e91",
			4003 => x"fe1a3e91",
			4004 => x"08002320",
			4005 => x"01000e04",
			4006 => x"fe5e3f25",
			4007 => x"0f00bb14",
			4008 => x"0f00820c",
			4009 => x"01001204",
			4010 => x"fe623f25",
			4011 => x"07002b04",
			4012 => x"002b3f25",
			4013 => x"fe823f25",
			4014 => x"0000f304",
			4015 => x"020d3f25",
			4016 => x"ffe63f25",
			4017 => x"0e00a004",
			4018 => x"fe1b3f25",
			4019 => x"ffb43f25",
			4020 => x"0f006504",
			4021 => x"fe653f25",
			4022 => x"03004624",
			4023 => x"07003f14",
			4024 => x"02013710",
			4025 => x"0f00af08",
			4026 => x"0b001e04",
			4027 => x"02653f25",
			4028 => x"01513f25",
			4029 => x"07003704",
			4030 => x"ffd03f25",
			4031 => x"01433f25",
			4032 => x"fef83f25",
			4033 => x"05003508",
			4034 => x"00014104",
			4035 => x"01bd3f25",
			4036 => x"00313f25",
			4037 => x"0c001f04",
			4038 => x"025c3f25",
			4039 => x"01be3f25",
			4040 => x"fe473f25",
			4041 => x"08002324",
			4042 => x"0f00a81c",
			4043 => x"06008014",
			4044 => x"01001004",
			4045 => x"ff3a3fc9",
			4046 => x"07002a08",
			4047 => x"03002404",
			4048 => x"00453fc9",
			4049 => x"ff703fc9",
			4050 => x"06006e04",
			4051 => x"ffea3fc9",
			4052 => x"00743fc9",
			4053 => x"01000c04",
			4054 => x"ffd83fc9",
			4055 => x"00a63fc9",
			4056 => x"04002a04",
			4057 => x"fedd3fc9",
			4058 => x"00673fc9",
			4059 => x"0300452c",
			4060 => x"05003920",
			4061 => x"0a00371c",
			4062 => x"0b001f10",
			4063 => x"0f00c008",
			4064 => x"0200fd04",
			4065 => x"fff83fc9",
			4066 => x"00c13fc9",
			4067 => x"0c001d04",
			4068 => x"00393fc9",
			4069 => x"ff3d3fc9",
			4070 => x"0000f404",
			4071 => x"ffc43fc9",
			4072 => x"0e00a204",
			4073 => x"01113fc9",
			4074 => x"00163fc9",
			4075 => x"ff653fc9",
			4076 => x"0c001c04",
			4077 => x"00243fc9",
			4078 => x"0e008404",
			4079 => x"00033fc9",
			4080 => x"010b3fc9",
			4081 => x"ff403fc9",
			4082 => x"08002224",
			4083 => x"0b00150c",
			4084 => x"04001e04",
			4085 => x"ffb8408d",
			4086 => x"01000e04",
			4087 => x"ffeb408d",
			4088 => x"0067408d",
			4089 => x"02009008",
			4090 => x"02008c04",
			4091 => x"ffec408d",
			4092 => x"0028408d",
			4093 => x"07003c0c",
			4094 => x"04001908",
			4095 => x"04001804",
			4096 => x"fffa408d",
			4097 => x"000e408d",
			4098 => x"ff4a408d",
			4099 => x"0011408d",
			4100 => x"0a004334",
			4101 => x"05003928",
			4102 => x"02013720",
			4103 => x"08002610",
			4104 => x"0a002d08",
			4105 => x"07002c04",
			4106 => x"ffe2408d",
			4107 => x"0089408d",
			4108 => x"09002204",
			4109 => x"0022408d",
			4110 => x"ff95408d",
			4111 => x"0c002208",
			4112 => x"00012704",
			4113 => x"fffc408d",
			4114 => x"00cc408d",
			4115 => x"0600b604",
			4116 => x"ff98408d",
			4117 => x"0047408d",
			4118 => x"07004004",
			4119 => x"ff63408d",
			4120 => x"0060408d",
			4121 => x"0f00b808",
			4122 => x"00011b04",
			4123 => x"0034408d",
			4124 => x"ffc0408d",
			4125 => x"00b6408d",
			4126 => x"01001808",
			4127 => x"07004104",
			4128 => x"ffa0408d",
			4129 => x"0003408d",
			4130 => x"0007408d",
			4131 => x"08002648",
			4132 => x"0a002d10",
			4133 => x"09001d04",
			4134 => x"ffd14169",
			4135 => x"06006504",
			4136 => x"ffe74169",
			4137 => x"08001f04",
			4138 => x"fffc4169",
			4139 => x"00714169",
			4140 => x"05003a1c",
			4141 => x"0000d108",
			4142 => x"0000a104",
			4143 => x"ffee4169",
			4144 => x"00284169",
			4145 => x"02014110",
			4146 => x"04001b08",
			4147 => x"00012604",
			4148 => x"fffe4169",
			4149 => x"00114169",
			4150 => x"00014204",
			4151 => x"ff724169",
			4152 => x"fff54169",
			4153 => x"000f4169",
			4154 => x"0a004014",
			4155 => x"0f00b80c",
			4156 => x"0a003d08",
			4157 => x"05003e04",
			4158 => x"00054169",
			4159 => x"ffcf4169",
			4160 => x"00104169",
			4161 => x"0d001904",
			4162 => x"00004169",
			4163 => x"00744169",
			4164 => x"07003f04",
			4165 => x"ffba4169",
			4166 => x"00024169",
			4167 => x"04002110",
			4168 => x"0300270c",
			4169 => x"08002704",
			4170 => x"fff84169",
			4171 => x"0b002504",
			4172 => x"00344169",
			4173 => x"fffa4169",
			4174 => x"ffc64169",
			4175 => x"01001408",
			4176 => x"0200e304",
			4177 => x"00024169",
			4178 => x"ffec4169",
			4179 => x"08002d08",
			4180 => x"03004404",
			4181 => x"00ca4169",
			4182 => x"fffd4169",
			4183 => x"0e009504",
			4184 => x"ffdc4169",
			4185 => x"00234169",
			4186 => x"07003f40",
			4187 => x"02013734",
			4188 => x"01000c04",
			4189 => x"feaa4215",
			4190 => x"09002518",
			4191 => x"09002410",
			4192 => x"02011c08",
			4193 => x"07002904",
			4194 => x"fed24215",
			4195 => x"00a64215",
			4196 => x"0600ad04",
			4197 => x"fea74215",
			4198 => x"00b64215",
			4199 => x"0f009304",
			4200 => x"ffc94215",
			4201 => x"01684215",
			4202 => x"03002a0c",
			4203 => x"01001608",
			4204 => x"0c002004",
			4205 => x"010a4215",
			4206 => x"ff914215",
			4207 => x"fe934215",
			4208 => x"05003304",
			4209 => x"01574215",
			4210 => x"01001704",
			4211 => x"ff454215",
			4212 => x"013a4215",
			4213 => x"0e009904",
			4214 => x"fea44215",
			4215 => x"03002c04",
			4216 => x"ff234215",
			4217 => x"004e4215",
			4218 => x"0c002108",
			4219 => x"02013f04",
			4220 => x"01694215",
			4221 => x"009e4215",
			4222 => x"0d002108",
			4223 => x"05004104",
			4224 => x"ff074215",
			4225 => x"00334215",
			4226 => x"02010a04",
			4227 => x"ffad4215",
			4228 => x"01344215",
			4229 => x"0700404c",
			4230 => x"0c001e38",
			4231 => x"07003728",
			4232 => x"02011814",
			4233 => x"07002904",
			4234 => x"ff3642d9",
			4235 => x"0a003708",
			4236 => x"09002104",
			4237 => x"002a42d9",
			4238 => x"010942d9",
			4239 => x"09002404",
			4240 => x"ff5542d9",
			4241 => x"004542d9",
			4242 => x"0600a208",
			4243 => x"0600a004",
			4244 => x"ffaf42d9",
			4245 => x"007842d9",
			4246 => x"01001008",
			4247 => x"05003604",
			4248 => x"ff7342d9",
			4249 => x"004842d9",
			4250 => x"fece42d9",
			4251 => x"05003004",
			4252 => x"ff7142d9",
			4253 => x"00014308",
			4254 => x"0600aa04",
			4255 => x"004442d9",
			4256 => x"012b42d9",
			4257 => x"ffd342d9",
			4258 => x"0f00c30c",
			4259 => x"06009504",
			4260 => x"ff7842d9",
			4261 => x"07003d04",
			4262 => x"00ed42d9",
			4263 => x"ffef42d9",
			4264 => x"05003804",
			4265 => x"ff0a42d9",
			4266 => x"005f42d9",
			4267 => x"0c002104",
			4268 => x"010a42d9",
			4269 => x"08002b0c",
			4270 => x"03003104",
			4271 => x"ff8142d9",
			4272 => x"03007504",
			4273 => x"005242d9",
			4274 => x"fff142d9",
			4275 => x"00011604",
			4276 => x"ffe442d9",
			4277 => x"00a042d9",
			4278 => x"08002224",
			4279 => x"0b00150c",
			4280 => x"04001e04",
			4281 => x"ffb643b5",
			4282 => x"0d001504",
			4283 => x"fff143b5",
			4284 => x"006343b5",
			4285 => x"02009008",
			4286 => x"02008c04",
			4287 => x"ffeb43b5",
			4288 => x"002943b5",
			4289 => x"07003c0c",
			4290 => x"04001908",
			4291 => x"04001804",
			4292 => x"fffa43b5",
			4293 => x"000f43b5",
			4294 => x"ff4243b5",
			4295 => x"001243b5",
			4296 => x"0a003b38",
			4297 => x"0201372c",
			4298 => x"08002618",
			4299 => x"0c001e0c",
			4300 => x"0e008808",
			4301 => x"04002304",
			4302 => x"004543b5",
			4303 => x"ffa543b5",
			4304 => x"008543b5",
			4305 => x"09002804",
			4306 => x"ff6643b5",
			4307 => x"09002904",
			4308 => x"002543b5",
			4309 => x"fff543b5",
			4310 => x"01001a0c",
			4311 => x"0e009d08",
			4312 => x"06007504",
			4313 => x"fff143b5",
			4314 => x"010c43b5",
			4315 => x"ffef43b5",
			4316 => x"00012a04",
			4317 => x"ffb543b5",
			4318 => x"002543b5",
			4319 => x"07004004",
			4320 => x"ff7643b5",
			4321 => x"01001a04",
			4322 => x"007e43b5",
			4323 => x"fffb43b5",
			4324 => x"04002e0c",
			4325 => x"05003f04",
			4326 => x"ff6a43b5",
			4327 => x"0e009804",
			4328 => x"002343b5",
			4329 => x"ffde43b5",
			4330 => x"03004604",
			4331 => x"009343b5",
			4332 => x"ff9d43b5",
			4333 => x"08002338",
			4334 => x"0e008930",
			4335 => x"07002f20",
			4336 => x"0a002a14",
			4337 => x"0400200c",
			4338 => x"0c001704",
			4339 => x"ff8e4499",
			4340 => x"0c001904",
			4341 => x"002f4499",
			4342 => x"ffe54499",
			4343 => x"05002d04",
			4344 => x"00784499",
			4345 => x"fff14499",
			4346 => x"0b001508",
			4347 => x"0b001404",
			4348 => x"ffd14499",
			4349 => x"00104499",
			4350 => x"ff3c4499",
			4351 => x"0400360c",
			4352 => x"00012508",
			4353 => x"01000e04",
			4354 => x"fff54499",
			4355 => x"00bc4499",
			4356 => x"ffd94499",
			4357 => x"ffd04499",
			4358 => x"0e00a504",
			4359 => x"fefe4499",
			4360 => x"002a4499",
			4361 => x"0a003b24",
			4362 => x"00014618",
			4363 => x"0e008a0c",
			4364 => x"0f00b008",
			4365 => x"0f006504",
			4366 => x"ffc14499",
			4367 => x"009f4499",
			4368 => x"ffa24499",
			4369 => x"0c001e04",
			4370 => x"011f4499",
			4371 => x"08002904",
			4372 => x"ffa84499",
			4373 => x"00c84499",
			4374 => x"0d001f04",
			4375 => x"ff4c4499",
			4376 => x"04002704",
			4377 => x"00a34499",
			4378 => x"fff14499",
			4379 => x"0600b714",
			4380 => x"0100170c",
			4381 => x"00012a08",
			4382 => x"00010804",
			4383 => x"ffe24499",
			4384 => x"00174499",
			4385 => x"ff364499",
			4386 => x"00011604",
			4387 => x"fff54499",
			4388 => x"002c4499",
			4389 => x"006e4499",
			4390 => x"08002324",
			4391 => x"0f00a81c",
			4392 => x"06008014",
			4393 => x"01001004",
			4394 => x"ff434555",
			4395 => x"07002a08",
			4396 => x"03002404",
			4397 => x"00404555",
			4398 => x"ff784555",
			4399 => x"06006e04",
			4400 => x"ffeb4555",
			4401 => x"00704555",
			4402 => x"01000c04",
			4403 => x"ffd94555",
			4404 => x"009d4555",
			4405 => x"04002a04",
			4406 => x"fee84555",
			4407 => x"00634555",
			4408 => x"03004538",
			4409 => x"0500391c",
			4410 => x"03003114",
			4411 => x"03002e0c",
			4412 => x"0c001b04",
			4413 => x"009a4555",
			4414 => x"0d001f04",
			4415 => x"ff754555",
			4416 => x"00904555",
			4417 => x"02011e04",
			4418 => x"ffbe4555",
			4419 => x"01084555",
			4420 => x"0a003604",
			4421 => x"00394555",
			4422 => x"ff5b4555",
			4423 => x"03003510",
			4424 => x"0a00380c",
			4425 => x"0a003604",
			4426 => x"005a4555",
			4427 => x"0600ad04",
			4428 => x"ffb34555",
			4429 => x"00234555",
			4430 => x"01134555",
			4431 => x"05004104",
			4432 => x"ff644555",
			4433 => x"0600a604",
			4434 => x"00094555",
			4435 => x"00b04555",
			4436 => x"ff464555",
			4437 => x"08002328",
			4438 => x"03003320",
			4439 => x"0600901c",
			4440 => x"06008014",
			4441 => x"0500360c",
			4442 => x"02009008",
			4443 => x"00009204",
			4444 => x"ffeb4629",
			4445 => x"00144629",
			4446 => x"ffb44629",
			4447 => x"0000aa04",
			4448 => x"fff24629",
			4449 => x"00154629",
			4450 => x"03002404",
			4451 => x"fff74629",
			4452 => x"004e4629",
			4453 => x"ff6a4629",
			4454 => x"0a003704",
			4455 => x"00484629",
			4456 => x"ffda4629",
			4457 => x"02013734",
			4458 => x"0300311c",
			4459 => x"09002508",
			4460 => x"0f006504",
			4461 => x"fff94629",
			4462 => x"009f4629",
			4463 => x"0400210c",
			4464 => x"08002a08",
			4465 => x"04001a04",
			4466 => x"000e4629",
			4467 => x"ff8d4629",
			4468 => x"000e4629",
			4469 => x"0c001f04",
			4470 => x"00024629",
			4471 => x"007b4629",
			4472 => x"05003804",
			4473 => x"ffae4629",
			4474 => x"03003808",
			4475 => x"0a003804",
			4476 => x"fff24629",
			4477 => x"00684629",
			4478 => x"07003904",
			4479 => x"ffba4629",
			4480 => x"03004604",
			4481 => x"00304629",
			4482 => x"ffde4629",
			4483 => x"0b00210c",
			4484 => x"03002e04",
			4485 => x"ff7c4629",
			4486 => x"0600bc04",
			4487 => x"ffd34629",
			4488 => x"00434629",
			4489 => x"00414629",
			4490 => x"0e009448",
			4491 => x"0001313c",
			4492 => x"0e009134",
			4493 => x"01001420",
			4494 => x"04002110",
			4495 => x"04001d08",
			4496 => x"01001204",
			4497 => x"ff834705",
			4498 => x"001b4705",
			4499 => x"01000e04",
			4500 => x"ffe74705",
			4501 => x"00f04705",
			4502 => x"03002d08",
			4503 => x"05003304",
			4504 => x"ff804705",
			4505 => x"007a4705",
			4506 => x"08002304",
			4507 => x"ffca4705",
			4508 => x"ff194705",
			4509 => x"0200fd10",
			4510 => x"01001508",
			4511 => x"07003404",
			4512 => x"00324705",
			4513 => x"fffa4705",
			4514 => x"03002704",
			4515 => x"001e4705",
			4516 => x"ff6a4705",
			4517 => x"012d4705",
			4518 => x"05003804",
			4519 => x"ff134705",
			4520 => x"002a4705",
			4521 => x"0b001c08",
			4522 => x"04002904",
			4523 => x"fec34705",
			4524 => x"fff24705",
			4525 => x"003a4705",
			4526 => x"03002e18",
			4527 => x"0a002f08",
			4528 => x"04001804",
			4529 => x"ffe44705",
			4530 => x"00e24705",
			4531 => x"02013308",
			4532 => x"01001204",
			4533 => x"fff04705",
			4534 => x"00b94705",
			4535 => x"0f00dc04",
			4536 => x"fefb4705",
			4537 => x"ffd64705",
			4538 => x"0a003b08",
			4539 => x"0b001804",
			4540 => x"ffb74705",
			4541 => x"011e4705",
			4542 => x"0e009904",
			4543 => x"ff544705",
			4544 => x"008e4705",
			4545 => x"08002760",
			4546 => x"0d001b38",
			4547 => x"0c001a20",
			4548 => x"09002118",
			4549 => x"0200ca0c",
			4550 => x"07002904",
			4551 => x"ff5d4819",
			4552 => x"0b001404",
			4553 => x"ffa64819",
			4554 => x"00da4819",
			4555 => x"05003a04",
			4556 => x"fed54819",
			4557 => x"05003e04",
			4558 => x"00424819",
			4559 => x"ffef4819",
			4560 => x"0a003704",
			4561 => x"00da4819",
			4562 => x"ffc24819",
			4563 => x"05003a0c",
			4564 => x"06009608",
			4565 => x"0000c204",
			4566 => x"ffd04819",
			4567 => x"00084819",
			4568 => x"fec24819",
			4569 => x"0a003b04",
			4570 => x"007a4819",
			4571 => x"07003904",
			4572 => x"ff204819",
			4573 => x"003f4819",
			4574 => x"0001261c",
			4575 => x"09002508",
			4576 => x"0000b004",
			4577 => x"ffdf4819",
			4578 => x"00514819",
			4579 => x"0500380c",
			4580 => x"09002804",
			4581 => x"fecc4819",
			4582 => x"0c002104",
			4583 => x"00544819",
			4584 => x"ffe04819",
			4585 => x"00010404",
			4586 => x"ffde4819",
			4587 => x"00764819",
			4588 => x"02013004",
			4589 => x"011c4819",
			4590 => x"0c001d04",
			4591 => x"00154819",
			4592 => x"ff504819",
			4593 => x"07003e10",
			4594 => x"03002a08",
			4595 => x"0b002404",
			4596 => x"00064819",
			4597 => x"fff34819",
			4598 => x"03003a04",
			4599 => x"01214819",
			4600 => x"fffd4819",
			4601 => x"0600b60c",
			4602 => x"00013608",
			4603 => x"06009e04",
			4604 => x"ffd64819",
			4605 => x"00624819",
			4606 => x"ff114819",
			4607 => x"01001804",
			4608 => x"ffe74819",
			4609 => x"01001a04",
			4610 => x"00f14819",
			4611 => x"01001d04",
			4612 => x"ffc14819",
			4613 => x"006f4819",
			4614 => x"08001f04",
			4615 => x"fecc48bd",
			4616 => x"00012228",
			4617 => x"0600801c",
			4618 => x"0d001914",
			4619 => x"01000e0c",
			4620 => x"04002008",
			4621 => x"07002904",
			4622 => x"ffee48bd",
			4623 => x"008c48bd",
			4624 => x"ffc548bd",
			4625 => x"05002704",
			4626 => x"004048bd",
			4627 => x"febb48bd",
			4628 => x"0b001b04",
			4629 => x"00ec48bd",
			4630 => x"ff2848bd",
			4631 => x"0a003704",
			4632 => x"015548bd",
			4633 => x"05004504",
			4634 => x"ff2248bd",
			4635 => x"008d48bd",
			4636 => x"09002b20",
			4637 => x"08002308",
			4638 => x"00014b04",
			4639 => x"fe7e48bd",
			4640 => x"004f48bd",
			4641 => x"0500380c",
			4642 => x"05003608",
			4643 => x"02013504",
			4644 => x"007948bd",
			4645 => x"ff1548bd",
			4646 => x"fed248bd",
			4647 => x"07003b08",
			4648 => x"05003c04",
			4649 => x"004148bd",
			4650 => x"ff8048bd",
			4651 => x"014d48bd",
			4652 => x"0f00bf04",
			4653 => x"ffcc48bd",
			4654 => x"016248bd",
			4655 => x"08001f0c",
			4656 => x"01000e04",
			4657 => x"fead4969",
			4658 => x"05002e04",
			4659 => x"ff224969",
			4660 => x"00334969",
			4661 => x"0a003b34",
			4662 => x"05003a30",
			4663 => x"0f00c018",
			4664 => x"06009e10",
			4665 => x"0a002d08",
			4666 => x"06006504",
			4667 => x"ff3e4969",
			4668 => x"01324969",
			4669 => x"06009704",
			4670 => x"002b4969",
			4671 => x"fee34969",
			4672 => x"09002104",
			4673 => x"ff194969",
			4674 => x"016f4969",
			4675 => x"0e00940c",
			4676 => x"05003004",
			4677 => x"fe7e4969",
			4678 => x"03002f04",
			4679 => x"004d4969",
			4680 => x"feed4969",
			4681 => x"0a003104",
			4682 => x"01324969",
			4683 => x"04002704",
			4684 => x"ff504969",
			4685 => x"00df4969",
			4686 => x"01544969",
			4687 => x"0e009914",
			4688 => x"0100170c",
			4689 => x"04002e04",
			4690 => x"feba4969",
			4691 => x"05004e04",
			4692 => x"00834969",
			4693 => x"ff154969",
			4694 => x"0a004a04",
			4695 => x"00ae4969",
			4696 => x"ffdd4969",
			4697 => x"011f4969",
			4698 => x"01000c04",
			4699 => x"fe8049ed",
			4700 => x"0a003118",
			4701 => x"06006504",
			4702 => x"fec449ed",
			4703 => x"09001d04",
			4704 => x"fed549ed",
			4705 => x"0f00aa04",
			4706 => x"01a349ed",
			4707 => x"09002104",
			4708 => x"fe8449ed",
			4709 => x"0c001f04",
			4710 => x"015249ed",
			4711 => x"007e49ed",
			4712 => x"05003004",
			4713 => x"fe4f49ed",
			4714 => x"08002208",
			4715 => x"07003b04",
			4716 => x"fe5549ed",
			4717 => x"009649ed",
			4718 => x"02011a10",
			4719 => x"0a003708",
			4720 => x"00010c04",
			4721 => x"006649ed",
			4722 => x"017249ed",
			4723 => x"04002904",
			4724 => x"fec549ed",
			4725 => x"009e49ed",
			4726 => x"07003704",
			4727 => x"ff0b49ed",
			4728 => x"0600af04",
			4729 => x"014049ed",
			4730 => x"ffca49ed",
			4731 => x"0d001920",
			4732 => x"07002a04",
			4733 => x"ff344a99",
			4734 => x"02011c14",
			4735 => x"0a003710",
			4736 => x"09001d04",
			4737 => x"ffaf4a99",
			4738 => x"0d001504",
			4739 => x"ffce4a99",
			4740 => x"01000c04",
			4741 => x"ffeb4a99",
			4742 => x"00d24a99",
			4743 => x"ff874a99",
			4744 => x"0e00a404",
			4745 => x"ff2c4a99",
			4746 => x"001d4a99",
			4747 => x"03004534",
			4748 => x"0500392c",
			4749 => x"01001410",
			4750 => x"0a00340c",
			4751 => x"0b001c08",
			4752 => x"08002004",
			4753 => x"ffd54a99",
			4754 => x"00c84a99",
			4755 => x"ffa44a99",
			4756 => x"ff1b4a99",
			4757 => x"04002110",
			4758 => x"04001d08",
			4759 => x"0c002604",
			4760 => x"00b34a99",
			4761 => x"ffe54a99",
			4762 => x"0e009304",
			4763 => x"ff564a99",
			4764 => x"ffe64a99",
			4765 => x"02013708",
			4766 => x"0a003204",
			4767 => x"00204a99",
			4768 => x"013b4a99",
			4769 => x"ffc14a99",
			4770 => x"01001204",
			4771 => x"fffe4a99",
			4772 => x"01114a99",
			4773 => x"ff4f4a99",
			4774 => x"09001d04",
			4775 => x"fea94b2d",
			4776 => x"0b001508",
			4777 => x"0000b704",
			4778 => x"ffff4b2d",
			4779 => x"016b4b2d",
			4780 => x"07003f28",
			4781 => x"08002214",
			4782 => x"0a002c0c",
			4783 => x"0d001704",
			4784 => x"ff484b2d",
			4785 => x"07002e04",
			4786 => x"00bf4b2d",
			4787 => x"ffb94b2d",
			4788 => x"04001b04",
			4789 => x"00024b2d",
			4790 => x"fe844b2d",
			4791 => x"02013710",
			4792 => x"09002508",
			4793 => x"07003704",
			4794 => x"00014b2d",
			4795 => x"01624b2d",
			4796 => x"03002a04",
			4797 => x"ff044b2d",
			4798 => x"001a4b2d",
			4799 => x"ff004b2d",
			4800 => x"0c002108",
			4801 => x"02013f04",
			4802 => x"01634b2d",
			4803 => x"00914b2d",
			4804 => x"0d002108",
			4805 => x"05004104",
			4806 => x"ff1a4b2d",
			4807 => x"002f4b2d",
			4808 => x"02010a04",
			4809 => x"ffb34b2d",
			4810 => x"012b4b2d",
			4811 => x"0700405c",
			4812 => x"0f00c13c",
			4813 => x"01001430",
			4814 => x"04002114",
			4815 => x"01000e08",
			4816 => x"08002304",
			4817 => x"ff554c11",
			4818 => x"00594c11",
			4819 => x"06008108",
			4820 => x"09001e04",
			4821 => x"ff824c11",
			4822 => x"00564c11",
			4823 => x"00e44c11",
			4824 => x"07003510",
			4825 => x"0b001508",
			4826 => x"03002904",
			4827 => x"ffbd4c11",
			4828 => x"00404c11",
			4829 => x"09002404",
			4830 => x"fef34c11",
			4831 => x"00044c11",
			4832 => x"07003604",
			4833 => x"008a4c11",
			4834 => x"0d001c04",
			4835 => x"ff4d4c11",
			4836 => x"00344c11",
			4837 => x"0b001a04",
			4838 => x"ffc04c11",
			4839 => x"09002c04",
			4840 => x"012e4c11",
			4841 => x"ffac4c11",
			4842 => x"05003818",
			4843 => x"03002f14",
			4844 => x"03002e10",
			4845 => x"04001b08",
			4846 => x"0600b704",
			4847 => x"009f4c11",
			4848 => x"ffc54c11",
			4849 => x"04002304",
			4850 => x"feda4c11",
			4851 => x"ffb84c11",
			4852 => x"00f34c11",
			4853 => x"fed84c11",
			4854 => x"07003904",
			4855 => x"ffbd4c11",
			4856 => x"00d24c11",
			4857 => x"0c002104",
			4858 => x"00fe4c11",
			4859 => x"08002b0c",
			4860 => x"03003104",
			4861 => x"ff884c11",
			4862 => x"03007504",
			4863 => x"00504c11",
			4864 => x"fff14c11",
			4865 => x"00011604",
			4866 => x"ffe54c11",
			4867 => x"009a4c11",
			4868 => x"01000c04",
			4869 => x"fe844ca5",
			4870 => x"0a003118",
			4871 => x"06006504",
			4872 => x"fecf4ca5",
			4873 => x"09001d04",
			4874 => x"fede4ca5",
			4875 => x"05002f0c",
			4876 => x"0a002d08",
			4877 => x"06009b04",
			4878 => x"01bc4ca5",
			4879 => x"00e44ca5",
			4880 => x"00a44ca5",
			4881 => x"005e4ca5",
			4882 => x"05003004",
			4883 => x"fe5a4ca5",
			4884 => x"09002310",
			4885 => x"0b001808",
			4886 => x"0600a204",
			4887 => x"fec34ca5",
			4888 => x"01184ca5",
			4889 => x"04002d04",
			4890 => x"fe7c4ca5",
			4891 => x"00a24ca5",
			4892 => x"00013e0c",
			4893 => x"03002f04",
			4894 => x"01a74ca5",
			4895 => x"02011e04",
			4896 => x"ff6f4ca5",
			4897 => x"00e54ca5",
			4898 => x"04002708",
			4899 => x"07004304",
			4900 => x"febe4ca5",
			4901 => x"012d4ca5",
			4902 => x"04002b04",
			4903 => x"01914ca5",
			4904 => x"ff364ca5",
			4905 => x"0d001f78",
			4906 => x"05003444",
			4907 => x"0f00aa20",
			4908 => x"07002b0c",
			4909 => x"0d001904",
			4910 => x"ff1a4dd9",
			4911 => x"0c001c04",
			4912 => x"00714dd9",
			4913 => x"ffe74dd9",
			4914 => x"0000b70c",
			4915 => x"08002304",
			4916 => x"ff644dd9",
			4917 => x"0e002104",
			4918 => x"fffa4dd9",
			4919 => x"00584dd9",
			4920 => x"01000c04",
			4921 => x"ffce4dd9",
			4922 => x"01214dd9",
			4923 => x"0e008a10",
			4924 => x"04001e08",
			4925 => x"04001d04",
			4926 => x"ff784dd9",
			4927 => x"00444dd9",
			4928 => x"05002a04",
			4929 => x"ffda4dd9",
			4930 => x"feb14dd9",
			4931 => x"0f00c408",
			4932 => x"07003404",
			4933 => x"ff974dd9",
			4934 => x"01034dd9",
			4935 => x"0e009404",
			4936 => x"febc4dd9",
			4937 => x"0a002f04",
			4938 => x"00c54dd9",
			4939 => x"ff734dd9",
			4940 => x"0d001b24",
			4941 => x"0c001b10",
			4942 => x"0700330c",
			4943 => x"03002e08",
			4944 => x"07002a04",
			4945 => x"ffb94dd9",
			4946 => x"008c4dd9",
			4947 => x"ff1b4dd9",
			4948 => x"00dc4dd9",
			4949 => x"0c001d0c",
			4950 => x"07003308",
			4951 => x"07002e04",
			4952 => x"ffe44dd9",
			4953 => x"001d4dd9",
			4954 => x"fede4dd9",
			4955 => x"0c001e04",
			4956 => x"00544dd9",
			4957 => x"ff7d4dd9",
			4958 => x"0001430c",
			4959 => x"03004408",
			4960 => x"07003604",
			4961 => x"005f4dd9",
			4962 => x"014a4dd9",
			4963 => x"ff704dd9",
			4964 => x"ff694dd9",
			4965 => x"04002b10",
			4966 => x"08002d08",
			4967 => x"0000f404",
			4968 => x"ffd24dd9",
			4969 => x"01564dd9",
			4970 => x"0f00d404",
			4971 => x"ff654dd9",
			4972 => x"007f4dd9",
			4973 => x"0d002004",
			4974 => x"00b84dd9",
			4975 => x"01001708",
			4976 => x"08002704",
			4977 => x"00164dd9",
			4978 => x"fef64dd9",
			4979 => x"00011604",
			4980 => x"ffef4dd9",
			4981 => x"00754dd9",
			4982 => x"07003f70",
			4983 => x"08002650",
			4984 => x"0a00312c",
			4985 => x"09001e0c",
			4986 => x"05002208",
			4987 => x"0a002704",
			4988 => x"ffe54edf",
			4989 => x"00434edf",
			4990 => x"ff684edf",
			4991 => x"03002710",
			4992 => x"0a002708",
			4993 => x"0000b404",
			4994 => x"ffe34edf",
			4995 => x"004f4edf",
			4996 => x"0000a904",
			4997 => x"00324edf",
			4998 => x"ff8c4edf",
			4999 => x"04002008",
			5000 => x"05002a04",
			5001 => x"fff14edf",
			5002 => x"00bd4edf",
			5003 => x"03002c04",
			5004 => x"00514edf",
			5005 => x"ffae4edf",
			5006 => x"02011a14",
			5007 => x"05003408",
			5008 => x"0f00c104",
			5009 => x"ff5c4edf",
			5010 => x"00064edf",
			5011 => x"05003704",
			5012 => x"009c4edf",
			5013 => x"09002304",
			5014 => x"ff924edf",
			5015 => x"000b4edf",
			5016 => x"05003a0c",
			5017 => x"05003308",
			5018 => x"05003104",
			5019 => x"ff984edf",
			5020 => x"003c4edf",
			5021 => x"fee84edf",
			5022 => x"ffda4edf",
			5023 => x"03002a0c",
			5024 => x"01001608",
			5025 => x"04001804",
			5026 => x"fffb4edf",
			5027 => x"003f4edf",
			5028 => x"ff6d4edf",
			5029 => x"08002a0c",
			5030 => x"01001404",
			5031 => x"ffdd4edf",
			5032 => x"02010d04",
			5033 => x"00044edf",
			5034 => x"00ea4edf",
			5035 => x"0b001f04",
			5036 => x"003b4edf",
			5037 => x"ff5d4edf",
			5038 => x"03005310",
			5039 => x"01001a04",
			5040 => x"00ce4edf",
			5041 => x"0e00a108",
			5042 => x"01001d04",
			5043 => x"ffd24edf",
			5044 => x"00094edf",
			5045 => x"002e4edf",
			5046 => x"ffe14edf",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1715, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3321, initial_addr_3'length));
	end generate gen_rom_0;

	gen_rom_1: if SELECT_ROM = 1 generate
		bank <= (
			0 => x"0e008514",
			1 => x"01000810",
			2 => x"07002904",
			3 => x"ffda004d",
			4 => x"0000d508",
			5 => x"04002004",
			6 => x"0033004d",
			7 => x"fffd004d",
			8 => x"ffef004d",
			9 => x"ffb2004d",
			10 => x"02011308",
			11 => x"01001204",
			12 => x"005b004d",
			13 => x"fff5004d",
			14 => x"0600c904",
			15 => x"ff99004d",
			16 => x"03002d04",
			17 => x"0056004d",
			18 => x"ffe6004d",
			19 => x"0e009424",
			20 => x"0000f310",
			21 => x"0f007404",
			22 => x"ffc600b1",
			23 => x"05002a08",
			24 => x"01000b04",
			25 => x"007d00b1",
			26 => x"fffc00b1",
			27 => x"ffe600b1",
			28 => x"0400250c",
			29 => x"07003604",
			30 => x"ff8000b1",
			31 => x"07003a04",
			32 => x"000400b1",
			33 => x"fff900b1",
			34 => x"0600ab04",
			35 => x"ffe500b1",
			36 => x"001d00b1",
			37 => x"0001320c",
			38 => x"08001f08",
			39 => x"03002a04",
			40 => x"008400b1",
			41 => x"001600b1",
			42 => x"ffe100b1",
			43 => x"ffcf00b1",
			44 => x"03002a24",
			45 => x"07002e14",
			46 => x"0000b70c",
			47 => x"06006b04",
			48 => x"ffcb011d",
			49 => x"04001704",
			50 => x"004e011d",
			51 => x"0003011d",
			52 => x"0b001604",
			53 => x"ffab011d",
			54 => x"0000011d",
			55 => x"0001340c",
			56 => x"09001f08",
			57 => x"09001a04",
			58 => x"0026011d",
			59 => x"0094011d",
			60 => x"ffec011d",
			61 => x"ffdc011d",
			62 => x"0200f608",
			63 => x"0e007a04",
			64 => x"ffd8011d",
			65 => x"005d011d",
			66 => x"04002304",
			67 => x"ff36011d",
			68 => x"09002004",
			69 => x"003c011d",
			70 => x"ffdd011d",
			71 => x"0200f720",
			72 => x"0e006f14",
			73 => x"09001808",
			74 => x"00008904",
			75 => x"ffeb0199",
			76 => x"00230199",
			77 => x"0e006a04",
			78 => x"ffb80199",
			79 => x"08001d04",
			80 => x"000b0199",
			81 => x"fff70199",
			82 => x"05002a04",
			83 => x"009a0199",
			84 => x"01000904",
			85 => x"00080199",
			86 => x"fff00199",
			87 => x"0600bd10",
			88 => x"0c001704",
			89 => x"ff760199",
			90 => x"0e009104",
			91 => x"ffe00199",
			92 => x"09002104",
			93 => x"00480199",
			94 => x"fff80199",
			95 => x"03002a08",
			96 => x"00014004",
			97 => x"00650199",
			98 => x"ffe60199",
			99 => x"04002304",
			100 => x"ffa80199",
			101 => x"001b0199",
			102 => x"00010320",
			103 => x"0e007b18",
			104 => x"0400190c",
			105 => x"06006b04",
			106 => x"ffe8020d",
			107 => x"0000b504",
			108 => x"0030020d",
			109 => x"fffa020d",
			110 => x"03002108",
			111 => x"03001f04",
			112 => x"fffe020d",
			113 => x"0004020d",
			114 => x"ffca020d",
			115 => x"01000904",
			116 => x"fffe020d",
			117 => x"0064020d",
			118 => x"0e00a514",
			119 => x"03002f0c",
			120 => x"04002508",
			121 => x"07003904",
			122 => x"ff80020d",
			123 => x"0002020d",
			124 => x"0004020d",
			125 => x"09002004",
			126 => x"0042020d",
			127 => x"ffef020d",
			128 => x"03002d04",
			129 => x"0038020d",
			130 => x"ffdd020d",
			131 => x"0e009420",
			132 => x"0000f810",
			133 => x"0e006b04",
			134 => x"ffb80279",
			135 => x"05002d08",
			136 => x"01000b04",
			137 => x"00560279",
			138 => x"00070279",
			139 => x"fff20279",
			140 => x"0100060c",
			141 => x"04001d04",
			142 => x"fff40279",
			143 => x"01000504",
			144 => x"fffb0279",
			145 => x"00110279",
			146 => x"ff9c0279",
			147 => x"00011e04",
			148 => x"00700279",
			149 => x"0600ca0c",
			150 => x"0f00c804",
			151 => x"001a0279",
			152 => x"0a002d04",
			153 => x"ffff0279",
			154 => x"ff980279",
			155 => x"0600ce04",
			156 => x"004d0279",
			157 => x"ffe60279",
			158 => x"09001f28",
			159 => x"07002e10",
			160 => x"0000b70c",
			161 => x"06006b04",
			162 => x"fe9802e5",
			163 => x"0f008a04",
			164 => x"00c502e5",
			165 => x"015702e5",
			166 => x"fe8902e5",
			167 => x"00011e10",
			168 => x"04001804",
			169 => x"01d102e5",
			170 => x"0d001508",
			171 => x"01000a04",
			172 => x"018d02e5",
			173 => x"ff5f02e5",
			174 => x"014c02e5",
			175 => x"0600c904",
			176 => x"fe5f02e5",
			177 => x"007e02e5",
			178 => x"0100060c",
			179 => x"04002608",
			180 => x"00001304",
			181 => x"ffc102e5",
			182 => x"011f02e5",
			183 => x"feee02e5",
			184 => x"fe7502e5",
			185 => x"0e008528",
			186 => x"04001910",
			187 => x"06007004",
			188 => x"ff3e0369",
			189 => x"0000e908",
			190 => x"09001a04",
			191 => x"00e30369",
			192 => x"00240369",
			193 => x"ff730369",
			194 => x"07003010",
			195 => x"0300210c",
			196 => x"05002308",
			197 => x"03001a04",
			198 => x"ffe60369",
			199 => x"001b0369",
			200 => x"ffdd0369",
			201 => x"fed00369",
			202 => x"05002904",
			203 => x"00570369",
			204 => x"ff7a0369",
			205 => x"0201130c",
			206 => x"0a003408",
			207 => x"05002704",
			208 => x"01460369",
			209 => x"006e0369",
			210 => x"00170369",
			211 => x"0f00e308",
			212 => x"0d001104",
			213 => x"00b20369",
			214 => x"feb60369",
			215 => x"03002d04",
			216 => x"01040369",
			217 => x"ff5f0369",
			218 => x"0e006f14",
			219 => x"0b001308",
			220 => x"07002104",
			221 => x"fe9003cd",
			222 => x"012d03cd",
			223 => x"0e006c04",
			224 => x"fe5f03cd",
			225 => x"01000b04",
			226 => x"00a903cd",
			227 => x"fe7603cd",
			228 => x"0001321c",
			229 => x"09002218",
			230 => x"0200f70c",
			231 => x"0e007c08",
			232 => x"04001904",
			233 => x"01a203cd",
			234 => x"ff3a03cd",
			235 => x"01d003cd",
			236 => x"0e009104",
			237 => x"fe6c03cd",
			238 => x"03002a04",
			239 => x"01a603cd",
			240 => x"007903cd",
			241 => x"fe7b03cd",
			242 => x"fe6d03cd",
			243 => x"0600b02c",
			244 => x"0500200c",
			245 => x"06006b04",
			246 => x"ffe60449",
			247 => x"0000fc04",
			248 => x"003b0449",
			249 => x"fffb0449",
			250 => x"08001b10",
			251 => x"0700300c",
			252 => x"0200b508",
			253 => x"07002a04",
			254 => x"fff60449",
			255 => x"00150449",
			256 => x"ffd50449",
			257 => x"00200449",
			258 => x"01000808",
			259 => x"04001e04",
			260 => x"00100449",
			261 => x"fff10449",
			262 => x"04001604",
			263 => x"fff90449",
			264 => x"ff930449",
			265 => x"00011e04",
			266 => x"00620449",
			267 => x"04001708",
			268 => x"03002704",
			269 => x"00010449",
			270 => x"ffa70449",
			271 => x"04001b04",
			272 => x"004a0449",
			273 => x"ffe20449",
			274 => x"0e008528",
			275 => x"04001910",
			276 => x"06006b04",
			277 => x"ff2104cd",
			278 => x"0000b704",
			279 => x"011e04cd",
			280 => x"07002c04",
			281 => x"ff0b04cd",
			282 => x"008304cd",
			283 => x"0300210c",
			284 => x"07002b04",
			285 => x"ff8e04cd",
			286 => x"05001c04",
			287 => x"fff804cd",
			288 => x"006004cd",
			289 => x"07003004",
			290 => x"fe9404cd",
			291 => x"0e008004",
			292 => x"ff7504cd",
			293 => x"001304cd",
			294 => x"00013218",
			295 => x"03002a0c",
			296 => x"0d001408",
			297 => x"0e009204",
			298 => x"00e804cd",
			299 => x"003404cd",
			300 => x"016704cd",
			301 => x"05002d04",
			302 => x"ff7a04cd",
			303 => x"01001004",
			304 => x"013704cd",
			305 => x"ff5104cd",
			306 => x"fed604cd",
			307 => x"0e008524",
			308 => x"04001918",
			309 => x"0700290c",
			310 => x"09001708",
			311 => x"01000504",
			312 => x"00440561",
			313 => x"ffe00561",
			314 => x"ff8c0561",
			315 => x"00010408",
			316 => x"09001f04",
			317 => x"007e0561",
			318 => x"fff50561",
			319 => x"ffd40561",
			320 => x"03002108",
			321 => x"03001f04",
			322 => x"fff60561",
			323 => x"00070561",
			324 => x"ff530561",
			325 => x"02011314",
			326 => x"0a003410",
			327 => x"05002708",
			328 => x"05002404",
			329 => x"00330561",
			330 => x"00cb0561",
			331 => x"05002a04",
			332 => x"ffcc0561",
			333 => x"00640561",
			334 => x"ffca0561",
			335 => x"0600ca0c",
			336 => x"0d001104",
			337 => x"00330561",
			338 => x"03002404",
			339 => x"fff80561",
			340 => x"ff190561",
			341 => x"03002d04",
			342 => x"009c0561",
			343 => x"ffb70561",
			344 => x"0e009328",
			345 => x"0400160c",
			346 => x"06006b04",
			347 => x"ffda05cd",
			348 => x"0000fc04",
			349 => x"006905cd",
			350 => x"ffe805cd",
			351 => x"08001d18",
			352 => x"07003010",
			353 => x"03001d04",
			354 => x"000905cd",
			355 => x"05002204",
			356 => x"fffe05cd",
			357 => x"0600ad04",
			358 => x"ffb305cd",
			359 => x"fffe05cd",
			360 => x"05002f04",
			361 => x"004205cd",
			362 => x"fff605cd",
			363 => x"ff7c05cd",
			364 => x"0001320c",
			365 => x"01001008",
			366 => x"04001a04",
			367 => x"009205cd",
			368 => x"000e05cd",
			369 => x"ffeb05cd",
			370 => x"ffc705cd",
			371 => x"04001920",
			372 => x"02011210",
			373 => x"06006b04",
			374 => x"ff8b0661",
			375 => x"04001704",
			376 => x"01320661",
			377 => x"05002404",
			378 => x"ff790661",
			379 => x"00d40661",
			380 => x"0600ca0c",
			381 => x"08001804",
			382 => x"005a0661",
			383 => x"05002304",
			384 => x"ffed0661",
			385 => x"feed0661",
			386 => x"00900661",
			387 => x"0e008518",
			388 => x"07003410",
			389 => x"0300210c",
			390 => x"03001f08",
			391 => x"05002204",
			392 => x"ffe80661",
			393 => x"00040661",
			394 => x"00130661",
			395 => x"ff0a0661",
			396 => x"05002904",
			397 => x"002d0661",
			398 => x"ffcd0661",
			399 => x"0f00c408",
			400 => x"00011404",
			401 => x"00fa0661",
			402 => x"ff9c0661",
			403 => x"0d001504",
			404 => x"fefc0661",
			405 => x"00012d04",
			406 => x"008f0661",
			407 => x"ffa30661",
			408 => x"07003028",
			409 => x"09001b18",
			410 => x"00010314",
			411 => x"0700290c",
			412 => x"05001a08",
			413 => x"02006b04",
			414 => x"ff6106ed",
			415 => x"011706ed",
			416 => x"fe9c06ed",
			417 => x"07002c04",
			418 => x"00a906ed",
			419 => x"016a06ed",
			420 => x"fe9806ed",
			421 => x"0500220c",
			422 => x"05001e04",
			423 => x"ff1f06ed",
			424 => x"05001f04",
			425 => x"004806ed",
			426 => x"ffe906ed",
			427 => x"fe7c06ed",
			428 => x"0200f708",
			429 => x"09002204",
			430 => x"018106ed",
			431 => x"ff0806ed",
			432 => x"08001f10",
			433 => x"01000c08",
			434 => x"01000a04",
			435 => x"008806ed",
			436 => x"fe7c06ed",
			437 => x"0e009e04",
			438 => x"ffd806ed",
			439 => x"010b06ed",
			440 => x"00010e04",
			441 => x"00c706ed",
			442 => x"fe8906ed",
			443 => x"0600bd38",
			444 => x"0200eb14",
			445 => x"0e006a0c",
			446 => x"09001808",
			447 => x"0d001004",
			448 => x"fff00771",
			449 => x"00210771",
			450 => x"ffc00771",
			451 => x"05002d04",
			452 => x"004c0771",
			453 => x"fff20771",
			454 => x"0c001714",
			455 => x"04001d0c",
			456 => x"03002608",
			457 => x"03002304",
			458 => x"ffee0771",
			459 => x"00120771",
			460 => x"ff880771",
			461 => x"01000a04",
			462 => x"fff80771",
			463 => x"00130771",
			464 => x"01000b08",
			465 => x"0e008504",
			466 => x"fff60771",
			467 => x"003e0771",
			468 => x"04001e04",
			469 => x"00010771",
			470 => x"ffe70771",
			471 => x"0b001304",
			472 => x"ffe40771",
			473 => x"01001004",
			474 => x"00690771",
			475 => x"ffe10771",
			476 => x"08001c20",
			477 => x"07002b10",
			478 => x"0000a60c",
			479 => x"07002504",
			480 => x"ffe40805",
			481 => x"03001f04",
			482 => x"00290805",
			483 => x"00000805",
			484 => x"ffd00805",
			485 => x"0001320c",
			486 => x"0b001304",
			487 => x"00070805",
			488 => x"05004004",
			489 => x"00720805",
			490 => x"fff90805",
			491 => x"ffe80805",
			492 => x"0e009e20",
			493 => x"0b001308",
			494 => x"05002404",
			495 => x"fff80805",
			496 => x"00110805",
			497 => x"0200eb0c",
			498 => x"07003004",
			499 => x"ffd10805",
			500 => x"05002a04",
			501 => x"003d0805",
			502 => x"fff70805",
			503 => x"03003404",
			504 => x"ff860805",
			505 => x"05003b04",
			506 => x"00160805",
			507 => x"fff50805",
			508 => x"0a003104",
			509 => x"00470805",
			510 => x"0d001804",
			511 => x"ffb00805",
			512 => x"00280805",
			513 => x"0600b030",
			514 => x"0000f824",
			515 => x"0e007214",
			516 => x"09001808",
			517 => x"0a001c04",
			518 => x"ffcf0891",
			519 => x"00750891",
			520 => x"0e006a04",
			521 => x"ff3d0891",
			522 => x"01000804",
			523 => x"00280891",
			524 => x"ffbb0891",
			525 => x"0800220c",
			526 => x"05002a08",
			527 => x"0000bc04",
			528 => x"00130891",
			529 => x"00d50891",
			530 => x"fff50891",
			531 => x"ffe20891",
			532 => x"07003504",
			533 => x"ff180891",
			534 => x"08002004",
			535 => x"00360891",
			536 => x"ffaf0891",
			537 => x"00011e04",
			538 => x"00930891",
			539 => x"0600ca0c",
			540 => x"0f00c804",
			541 => x"00560891",
			542 => x"03002404",
			543 => x"00030891",
			544 => x"ff0a0891",
			545 => x"03002d04",
			546 => x"00a70891",
			547 => x"ff900891",
			548 => x"0600bd30",
			549 => x"0200f720",
			550 => x"0e007b18",
			551 => x"01000814",
			552 => x"0000b70c",
			553 => x"00008904",
			554 => x"fff308fd",
			555 => x"0b001504",
			556 => x"003208fd",
			557 => x"ffff08fd",
			558 => x"01000504",
			559 => x"ffe608fd",
			560 => x"000808fd",
			561 => x"ffc408fd",
			562 => x"07003304",
			563 => x"003e08fd",
			564 => x"000108fd",
			565 => x"0c001704",
			566 => x"ff9d08fd",
			567 => x"0e009104",
			568 => x"ffe608fd",
			569 => x"0b001904",
			570 => x"003008fd",
			571 => x"fffb08fd",
			572 => x"00013304",
			573 => x"003f08fd",
			574 => x"ffe208fd",
			575 => x"0e008524",
			576 => x"0900180c",
			577 => x"07002504",
			578 => x"ffdc0989",
			579 => x"0000fc04",
			580 => x"003f0989",
			581 => x"fff80989",
			582 => x"0700300c",
			583 => x"08001504",
			584 => x"00030989",
			585 => x"01000204",
			586 => x"00020989",
			587 => x"ff9e0989",
			588 => x"08001d08",
			589 => x"07003304",
			590 => x"00130989",
			591 => x"fffe0989",
			592 => x"ffee0989",
			593 => x"00013220",
			594 => x"03002a0c",
			595 => x"01000c08",
			596 => x"0200f104",
			597 => x"ffeb0989",
			598 => x"00180989",
			599 => x"008f0989",
			600 => x"0f00c810",
			601 => x"0f00c30c",
			602 => x"0f00bf08",
			603 => x"0a003604",
			604 => x"001d0989",
			605 => x"fff50989",
			606 => x"ffe50989",
			607 => x"00550989",
			608 => x"ffc80989",
			609 => x"ffbe0989",
			610 => x"07002e1c",
			611 => x"05001f10",
			612 => x"0a001c04",
			613 => x"ffd00a2d",
			614 => x"0000b708",
			615 => x"00008904",
			616 => x"fffc0a2d",
			617 => x"006c0a2d",
			618 => x"ffd50a2d",
			619 => x"03001d04",
			620 => x"00010a2d",
			621 => x"04001504",
			622 => x"fffe0a2d",
			623 => x"ff650a2d",
			624 => x"0a00311c",
			625 => x"05002910",
			626 => x"0d00180c",
			627 => x"0d001408",
			628 => x"0600b004",
			629 => x"ffce0a2d",
			630 => x"00550a2d",
			631 => x"00ec0a2d",
			632 => x"ffcb0a2d",
			633 => x"0f00c608",
			634 => x"0600a104",
			635 => x"ffee0a2d",
			636 => x"002d0a2d",
			637 => x"ffa80a2d",
			638 => x"01000a08",
			639 => x"05004104",
			640 => x"00770a2d",
			641 => x"ffec0a2d",
			642 => x"0f00e610",
			643 => x"0d001808",
			644 => x"0000f204",
			645 => x"00090a2d",
			646 => x"ff1e0a2d",
			647 => x"0600c204",
			648 => x"ffc30a2d",
			649 => x"00690a2d",
			650 => x"00560a2d",
			651 => x"0e008528",
			652 => x"04001914",
			653 => x"06006b04",
			654 => x"fe8d0ab9",
			655 => x"0000f40c",
			656 => x"0000ae04",
			657 => x"016c0ab9",
			658 => x"03002104",
			659 => x"ffb00ab9",
			660 => x"014e0ab9",
			661 => x"feb40ab9",
			662 => x"0700300c",
			663 => x"03002108",
			664 => x"0a002104",
			665 => x"ff220ab9",
			666 => x"007f0ab9",
			667 => x"fe620ab9",
			668 => x"05002d04",
			669 => x"00f30ab9",
			670 => x"fe9f0ab9",
			671 => x"0001321c",
			672 => x"0000f804",
			673 => x"019a0ab9",
			674 => x"0600b00c",
			675 => x"0f00bd08",
			676 => x"0a003604",
			677 => x"014d0ab9",
			678 => x"fee50ab9",
			679 => x"fe0a0ab9",
			680 => x"05002e08",
			681 => x"0c001504",
			682 => x"00e80ab9",
			683 => x"ff660ab9",
			684 => x"01ab0ab9",
			685 => x"fe860ab9",
			686 => x"0e009538",
			687 => x"0000f81c",
			688 => x"0e007b18",
			689 => x"01000810",
			690 => x"0f007404",
			691 => x"ff670b4d",
			692 => x"0000b704",
			693 => x"00ff0b4d",
			694 => x"0b001804",
			695 => x"ff9f0b4d",
			696 => x"00240b4d",
			697 => x"08001804",
			698 => x"fffa0b4d",
			699 => x"fef60b4d",
			700 => x"010a0b4d",
			701 => x"07003414",
			702 => x"03002408",
			703 => x"08001c04",
			704 => x"ff8b0b4d",
			705 => x"007d0b4d",
			706 => x"08001808",
			707 => x"04002504",
			708 => x"ffc30b4d",
			709 => x"004c0b4d",
			710 => x"fea80b4d",
			711 => x"01000b04",
			712 => x"009e0b4d",
			713 => x"ff7a0b4d",
			714 => x"08001f0c",
			715 => x"00012b04",
			716 => x"00ea0b4d",
			717 => x"0f00e704",
			718 => x"ff5b0b4d",
			719 => x"00920b4d",
			720 => x"0f00c404",
			721 => x"00030b4d",
			722 => x"ff210b4d",
			723 => x"03002a30",
			724 => x"0e009324",
			725 => x"00010a20",
			726 => x"08001c10",
			727 => x"07002504",
			728 => x"ffa70be9",
			729 => x"0d001608",
			730 => x"07002904",
			731 => x"001e0be9",
			732 => x"00cb0be9",
			733 => x"ffec0be9",
			734 => x"0b001408",
			735 => x"0c001304",
			736 => x"fffe0be9",
			737 => x"ff5c0be9",
			738 => x"0e006f04",
			739 => x"ffb60be9",
			740 => x"00480be9",
			741 => x"ff560be9",
			742 => x"08001f08",
			743 => x"00013404",
			744 => x"00c30be9",
			745 => x"ffcf0be9",
			746 => x"ffc80be9",
			747 => x"09001c10",
			748 => x"00013108",
			749 => x"0000e704",
			750 => x"00030be9",
			751 => x"fef50be9",
			752 => x"00013904",
			753 => x"005d0be9",
			754 => x"ffeb0be9",
			755 => x"0e009308",
			756 => x"05002e04",
			757 => x"002e0be9",
			758 => x"ff640be9",
			759 => x"00012a04",
			760 => x"00c40be9",
			761 => x"ffd10be9",
			762 => x"0e00852c",
			763 => x"04001914",
			764 => x"01000a10",
			765 => x"06006b04",
			766 => x"ff660c75",
			767 => x"0000b704",
			768 => x"01430c75",
			769 => x"07002c04",
			770 => x"ff260c75",
			771 => x"00a70c75",
			772 => x"ff2f0c75",
			773 => x"0300210c",
			774 => x"07002b04",
			775 => x"ff950c75",
			776 => x"05001c04",
			777 => x"fff80c75",
			778 => x"005c0c75",
			779 => x"07003004",
			780 => x"fe9a0c75",
			781 => x"0e008004",
			782 => x"ff810c75",
			783 => x"000f0c75",
			784 => x"00013218",
			785 => x"05002304",
			786 => x"01420c75",
			787 => x"05002504",
			788 => x"ff3d0c75",
			789 => x"0200f704",
			790 => x"01650c75",
			791 => x"0600c108",
			792 => x"0c001704",
			793 => x"feab0c75",
			794 => x"00c80c75",
			795 => x"00ac0c75",
			796 => x"fedf0c75",
			797 => x"0600770c",
			798 => x"09001708",
			799 => x"0d001004",
			800 => x"ff330ce1",
			801 => x"00ea0ce1",
			802 => x"fe760ce1",
			803 => x"0c001204",
			804 => x"01a60ce1",
			805 => x"05002108",
			806 => x"0b001304",
			807 => x"003b0ce1",
			808 => x"01720ce1",
			809 => x"0700300c",
			810 => x"00010108",
			811 => x"09001b04",
			812 => x"01000ce1",
			813 => x"fe920ce1",
			814 => x"fe800ce1",
			815 => x"0200ec08",
			816 => x"05002e04",
			817 => x"01750ce1",
			818 => x"ff650ce1",
			819 => x"01000a04",
			820 => x"00ea0ce1",
			821 => x"0a002d04",
			822 => x"01290ce1",
			823 => x"ff6c0ce1",
			824 => x"0600bd40",
			825 => x"00010328",
			826 => x"0e00721c",
			827 => x"0900180c",
			828 => x"0b001104",
			829 => x"ff8b0d75",
			830 => x"0e004704",
			831 => x"ffdd0d75",
			832 => x"00af0d75",
			833 => x"0d001108",
			834 => x"08001804",
			835 => x"00230d75",
			836 => x"ffe00d75",
			837 => x"08001604",
			838 => x"00030d75",
			839 => x"fed10d75",
			840 => x"0b001404",
			841 => x"ffd30d75",
			842 => x"05002e04",
			843 => x"01300d75",
			844 => x"ffc60d75",
			845 => x"03003810",
			846 => x"0e009e0c",
			847 => x"01000608",
			848 => x"04002204",
			849 => x"ff6d0d75",
			850 => x"00470d75",
			851 => x"fea00d75",
			852 => x"00050d75",
			853 => x"03003a04",
			854 => x"00a80d75",
			855 => x"ffac0d75",
			856 => x"0b001304",
			857 => x"ffdf0d75",
			858 => x"01001004",
			859 => x"01250d75",
			860 => x"ff3c0d75",
			861 => x"0600b03c",
			862 => x"0000f828",
			863 => x"0e007218",
			864 => x"09001808",
			865 => x"0a001c04",
			866 => x"ffcd0e19",
			867 => x"007d0e19",
			868 => x"0e006f0c",
			869 => x"01000204",
			870 => x"00010e19",
			871 => x"08001604",
			872 => x"00030e19",
			873 => x"ff360e19",
			874 => x"fff90e19",
			875 => x"0800220c",
			876 => x"05002a08",
			877 => x"0000bc04",
			878 => x"00130e19",
			879 => x"00de0e19",
			880 => x"fff50e19",
			881 => x"ffe00e19",
			882 => x"01000608",
			883 => x"0e008504",
			884 => x"ffb50e19",
			885 => x"002e0e19",
			886 => x"08001b08",
			887 => x"07002c04",
			888 => x"ffd00e19",
			889 => x"001f0e19",
			890 => x"fefd0e19",
			891 => x"00011e04",
			892 => x"00980e19",
			893 => x"0600ca0c",
			894 => x"0f00c804",
			895 => x"005a0e19",
			896 => x"03002404",
			897 => x"00030e19",
			898 => x"ff000e19",
			899 => x"03002d04",
			900 => x"00af0e19",
			901 => x"ff890e19",
			902 => x"0600770c",
			903 => x"09001808",
			904 => x"06004904",
			905 => x"fe8b0e9d",
			906 => x"016d0e9d",
			907 => x"fe5d0e9d",
			908 => x"00011e24",
			909 => x"09002220",
			910 => x"0e008010",
			911 => x"01000b0c",
			912 => x"0000e508",
			913 => x"0000c804",
			914 => x"01fb0e9d",
			915 => x"015c0e9d",
			916 => x"fe700e9d",
			917 => x"fe180e9d",
			918 => x"0c00170c",
			919 => x"0200f708",
			920 => x"07003204",
			921 => x"023a0e9d",
			922 => x"019e0e9d",
			923 => x"00640e9d",
			924 => x"02c00e9d",
			925 => x"fe700e9d",
			926 => x"0600c90c",
			927 => x"0d001108",
			928 => x"03002d04",
			929 => x"fe830e9d",
			930 => x"01c30e9d",
			931 => x"fe540e9d",
			932 => x"09001b04",
			933 => x"02300e9d",
			934 => x"fe610e9d",
			935 => x"0e009540",
			936 => x"0200ea24",
			937 => x"0e007218",
			938 => x"0900180c",
			939 => x"0d001004",
			940 => x"ffdb0f41",
			941 => x"03001504",
			942 => x"fff70f41",
			943 => x"005c0f41",
			944 => x"0d001104",
			945 => x"00090f41",
			946 => x"08001604",
			947 => x"00050f41",
			948 => x"ff6b0f41",
			949 => x"05002e08",
			950 => x"06008604",
			951 => x"00140f41",
			952 => x"00ae0f41",
			953 => x"fff10f41",
			954 => x"04001d04",
			955 => x"ff240f41",
			956 => x"0600ab10",
			957 => x"08001c0c",
			958 => x"04002208",
			959 => x"08001804",
			960 => x"fff70f41",
			961 => x"00250f41",
			962 => x"ffed0f41",
			963 => x"ff9d0f41",
			964 => x"09001f04",
			965 => x"00600f41",
			966 => x"ffe50f41",
			967 => x"08001f0c",
			968 => x"00011f04",
			969 => x"00ca0f41",
			970 => x"0f00e304",
			971 => x"ff7d0f41",
			972 => x"00690f41",
			973 => x"0f00c504",
			974 => x"00030f41",
			975 => x"ff900f41",
			976 => x"0e008b30",
			977 => x"05001a08",
			978 => x"00008904",
			979 => x"ffe40fe5",
			980 => x"003f0fe5",
			981 => x"07003120",
			982 => x"0e008618",
			983 => x"05001f10",
			984 => x"05001c08",
			985 => x"04001304",
			986 => x"00000fe5",
			987 => x"ffe20fe5",
			988 => x"04001304",
			989 => x"fffc0fe5",
			990 => x"001b0fe5",
			991 => x"04001604",
			992 => x"000a0fe5",
			993 => x"ff7a0fe5",
			994 => x"04002004",
			995 => x"fff10fe5",
			996 => x"000f0fe5",
			997 => x"04001e04",
			998 => x"00260fe5",
			999 => x"ffd50fe5",
			1000 => x"00011e0c",
			1001 => x"05002704",
			1002 => x"00bd0fe5",
			1003 => x"05002c04",
			1004 => x"fff00fe5",
			1005 => x"00500fe5",
			1006 => x"0600ca10",
			1007 => x"03003108",
			1008 => x"03002404",
			1009 => x"00010fe5",
			1010 => x"ff670fe5",
			1011 => x"0a003704",
			1012 => x"002a0fe5",
			1013 => x"fff80fe5",
			1014 => x"03002d04",
			1015 => x"00670fe5",
			1016 => x"ffc50fe5",
			1017 => x"0e008520",
			1018 => x"01000b1c",
			1019 => x"05002918",
			1020 => x"0700290c",
			1021 => x"05001a08",
			1022 => x"0a001b04",
			1023 => x"ff881061",
			1024 => x"00cc1061",
			1025 => x"ff031061",
			1026 => x"00010408",
			1027 => x"06007704",
			1028 => x"ffde1061",
			1029 => x"012a1061",
			1030 => x"ff7a1061",
			1031 => x"ff071061",
			1032 => x"febb1061",
			1033 => x"0001321c",
			1034 => x"03002604",
			1035 => x"011a1061",
			1036 => x"08001c08",
			1037 => x"0f00ca04",
			1038 => x"01361061",
			1039 => x"00441061",
			1040 => x"0d001504",
			1041 => x"ff7f1061",
			1042 => x"02011308",
			1043 => x"0a003204",
			1044 => x"01441061",
			1045 => x"00171061",
			1046 => x"ff1a1061",
			1047 => x"ff071061",
			1048 => x"09001f3c",
			1049 => x"0700290c",
			1050 => x"09001808",
			1051 => x"07002504",
			1052 => x"fe6e10ed",
			1053 => x"01b310ed",
			1054 => x"fe5710ed",
			1055 => x"0200f710",
			1056 => x"0e006a04",
			1057 => x"ff2510ed",
			1058 => x"08001d08",
			1059 => x"08001b04",
			1060 => x"025910ed",
			1061 => x"02d610ed",
			1062 => x"015a10ed",
			1063 => x"0600bd18",
			1064 => x"09001d10",
			1065 => x"03002408",
			1066 => x"0c001504",
			1067 => x"006810ed",
			1068 => x"fe7b10ed",
			1069 => x"0600ae04",
			1070 => x"fe6310ed",
			1071 => x"fdf510ed",
			1072 => x"0600a604",
			1073 => x"fe6f10ed",
			1074 => x"021910ed",
			1075 => x"07003304",
			1076 => x"041710ed",
			1077 => x"010810ed",
			1078 => x"08001d08",
			1079 => x"0e007a04",
			1080 => x"fe6210ed",
			1081 => x"027610ed",
			1082 => x"fe6010ed",
			1083 => x"08001c24",
			1084 => x"06006b04",
			1085 => x"ffe01181",
			1086 => x"0001321c",
			1087 => x"01000a10",
			1088 => x"0500400c",
			1089 => x"08001608",
			1090 => x"0d001104",
			1091 => x"fffa1181",
			1092 => x"00031181",
			1093 => x"006c1181",
			1094 => x"fffb1181",
			1095 => x"08001904",
			1096 => x"ffdf1181",
			1097 => x"05002704",
			1098 => x"003d1181",
			1099 => x"ffe81181",
			1100 => x"ffe61181",
			1101 => x"03002608",
			1102 => x"0e008604",
			1103 => x"ffd11181",
			1104 => x"00471181",
			1105 => x"0000f708",
			1106 => x"05002a04",
			1107 => x"00251181",
			1108 => x"fff01181",
			1109 => x"0400230c",
			1110 => x"07003808",
			1111 => x"0d001804",
			1112 => x"ff771181",
			1113 => x"00011181",
			1114 => x"00151181",
			1115 => x"0d001908",
			1116 => x"04002904",
			1117 => x"00261181",
			1118 => x"fff81181",
			1119 => x"fff01181",
			1120 => x"0e008628",
			1121 => x"01000b24",
			1122 => x"04001f1c",
			1123 => x"07002910",
			1124 => x"05001a0c",
			1125 => x"07002504",
			1126 => x"ffc71215",
			1127 => x"05001304",
			1128 => x"fffb1215",
			1129 => x"008c1215",
			1130 => x"ff651215",
			1131 => x"00010c08",
			1132 => x"06007704",
			1133 => x"fff51215",
			1134 => x"00c31215",
			1135 => x"ffbd1215",
			1136 => x"05002b04",
			1137 => x"00011215",
			1138 => x"ff7a1215",
			1139 => x"ff241215",
			1140 => x"00013220",
			1141 => x"0a003110",
			1142 => x"0500290c",
			1143 => x"05002508",
			1144 => x"0200ed04",
			1145 => x"00781215",
			1146 => x"fff81215",
			1147 => x"01181215",
			1148 => x"ffc31215",
			1149 => x"05002e04",
			1150 => x"ffba1215",
			1151 => x"0e009104",
			1152 => x"ffbe1215",
			1153 => x"07004004",
			1154 => x"00d91215",
			1155 => x"fff91215",
			1156 => x"ff651215",
			1157 => x"0e009338",
			1158 => x"0f00bd30",
			1159 => x"0e008528",
			1160 => x"04001910",
			1161 => x"06006b04",
			1162 => x"feec12b1",
			1163 => x"0000ae04",
			1164 => x"012e12b1",
			1165 => x"07002a04",
			1166 => x"fed212b1",
			1167 => x"00b612b1",
			1168 => x"07003110",
			1169 => x"05002208",
			1170 => x"03001a04",
			1171 => x"ffaa12b1",
			1172 => x"004c12b1",
			1173 => x"03001e04",
			1174 => x"fff912b1",
			1175 => x"fe8e12b1",
			1176 => x"05002e04",
			1177 => x"00b312b1",
			1178 => x"ff1c12b1",
			1179 => x"05002f04",
			1180 => x"016812b1",
			1181 => x"ff3712b1",
			1182 => x"05002204",
			1183 => x"ffe012b1",
			1184 => x"fe6d12b1",
			1185 => x"01001010",
			1186 => x"0f00e30c",
			1187 => x"00011f04",
			1188 => x"00e612b1",
			1189 => x"0e009904",
			1190 => x"00ca12b1",
			1191 => x"feb812b1",
			1192 => x"013212b1",
			1193 => x"03002904",
			1194 => x"005c12b1",
			1195 => x"fec612b1",
			1196 => x"0600b044",
			1197 => x"0000f82c",
			1198 => x"0e007220",
			1199 => x"09001808",
			1200 => x"0a001c04",
			1201 => x"ffce1375",
			1202 => x"00581375",
			1203 => x"07003110",
			1204 => x"08001608",
			1205 => x"01000404",
			1206 => x"00041375",
			1207 => x"fffd1375",
			1208 => x"0d001104",
			1209 => x"ffff1375",
			1210 => x"ff531375",
			1211 => x"0e006f04",
			1212 => x"fff11375",
			1213 => x"00111375",
			1214 => x"09001e04",
			1215 => x"00b11375",
			1216 => x"08002204",
			1217 => x"00071375",
			1218 => x"ffe91375",
			1219 => x"01000608",
			1220 => x"0e008504",
			1221 => x"ffcb1375",
			1222 => x"00251375",
			1223 => x"0e00940c",
			1224 => x"08001908",
			1225 => x"08001804",
			1226 => x"ffe21375",
			1227 => x"00131375",
			1228 => x"ff201375",
			1229 => x"00061375",
			1230 => x"0f00c804",
			1231 => x"00bd1375",
			1232 => x"0600bd0c",
			1233 => x"07003804",
			1234 => x"ff421375",
			1235 => x"0e009f04",
			1236 => x"fff01375",
			1237 => x"001c1375",
			1238 => x"07003408",
			1239 => x"00013404",
			1240 => x"00b01375",
			1241 => x"ffda1375",
			1242 => x"03002a04",
			1243 => x"003b1375",
			1244 => x"ff5b1375",
			1245 => x"0e00933c",
			1246 => x"00010a38",
			1247 => x"08001d1c",
			1248 => x"0e006b10",
			1249 => x"09001808",
			1250 => x"00008604",
			1251 => x"ff551441",
			1252 => x"00be1441",
			1253 => x"0d001104",
			1254 => x"000f1441",
			1255 => x"fea41441",
			1256 => x"03003108",
			1257 => x"07002c04",
			1258 => x"007e1441",
			1259 => x"016a1441",
			1260 => x"ff7a1441",
			1261 => x"04001608",
			1262 => x"0200ac04",
			1263 => x"ff7d1441",
			1264 => x"00ed1441",
			1265 => x"0400200c",
			1266 => x"05002108",
			1267 => x"05001d04",
			1268 => x"ffe51441",
			1269 => x"002e1441",
			1270 => x"fe8c1441",
			1271 => x"04002304",
			1272 => x"007b1441",
			1273 => x"ff261441",
			1274 => x"fe8f1441",
			1275 => x"03002a10",
			1276 => x"08001f08",
			1277 => x"00013404",
			1278 => x"01211441",
			1279 => x"ff6c1441",
			1280 => x"0e009b04",
			1281 => x"00831441",
			1282 => x"ff071441",
			1283 => x"0e00a618",
			1284 => x"03002f0c",
			1285 => x"03002d08",
			1286 => x"0e009b04",
			1287 => x"00021441",
			1288 => x"00e91441",
			1289 => x"fea51441",
			1290 => x"0e00a008",
			1291 => x"02011f04",
			1292 => x"01881441",
			1293 => x"ff911441",
			1294 => x"ff5e1441",
			1295 => x"fea81441",
			1296 => x"0600bd40",
			1297 => x"0f00c834",
			1298 => x"0600b030",
			1299 => x"0000f81c",
			1300 => x"0e006f10",
			1301 => x"09001808",
			1302 => x"0a001c04",
			1303 => x"ffde14cf",
			1304 => x"003d14cf",
			1305 => x"01000204",
			1306 => x"000314cf",
			1307 => x"ff8c14cf",
			1308 => x"05002a04",
			1309 => x"008014cf",
			1310 => x"08002004",
			1311 => x"000214cf",
			1312 => x"fff114cf",
			1313 => x"01000608",
			1314 => x"0e008304",
			1315 => x"ffe214cf",
			1316 => x"001c14cf",
			1317 => x"08001b08",
			1318 => x"0e008304",
			1319 => x"fff214cf",
			1320 => x"000d14cf",
			1321 => x"ff6514cf",
			1322 => x"008d14cf",
			1323 => x"07003804",
			1324 => x"ff7214cf",
			1325 => x"0e009f04",
			1326 => x"fff614cf",
			1327 => x"000f14cf",
			1328 => x"00013304",
			1329 => x"008814cf",
			1330 => x"ffc414cf",
			1331 => x"0e008514",
			1332 => x"04001910",
			1333 => x"07002904",
			1334 => x"ffd71519",
			1335 => x"00010408",
			1336 => x"01000a04",
			1337 => x"00301519",
			1338 => x"ffff1519",
			1339 => x"fff71519",
			1340 => x"ffb51519",
			1341 => x"02011308",
			1342 => x"01001204",
			1343 => x"00561519",
			1344 => x"fff51519",
			1345 => x"0600c904",
			1346 => x"ff9c1519",
			1347 => x"03002d04",
			1348 => x"00521519",
			1349 => x"ffe61519",
			1350 => x"0e00941c",
			1351 => x"0000f810",
			1352 => x"06007704",
			1353 => x"ffb6157d",
			1354 => x"05002d08",
			1355 => x"01000b04",
			1356 => x"0059157d",
			1357 => x"0002157d",
			1358 => x"fff0157d",
			1359 => x"0f00ad08",
			1360 => x"07003504",
			1361 => x"fff4157d",
			1362 => x"000d157d",
			1363 => x"ff99157d",
			1364 => x"00011e04",
			1365 => x"0076157d",
			1366 => x"0600ca0c",
			1367 => x"0f00c804",
			1368 => x"001b157d",
			1369 => x"0a002d04",
			1370 => x"ffff157d",
			1371 => x"ff94157d",
			1372 => x"0600ce04",
			1373 => x"0050157d",
			1374 => x"ffe5157d",
			1375 => x"0e008520",
			1376 => x"04001910",
			1377 => x"06007004",
			1378 => x"ff3315f1",
			1379 => x"0000e908",
			1380 => x"08001904",
			1381 => x"00ed15f1",
			1382 => x"002215f1",
			1383 => x"ff6b15f1",
			1384 => x"07003008",
			1385 => x"05002004",
			1386 => x"fffd15f1",
			1387 => x"fecf15f1",
			1388 => x"05002904",
			1389 => x"005b15f1",
			1390 => x"ff7215f1",
			1391 => x"0201130c",
			1392 => x"0a003408",
			1393 => x"05002704",
			1394 => x"015515f1",
			1395 => x"007115f1",
			1396 => x"001515f1",
			1397 => x"0f00e308",
			1398 => x"0d001104",
			1399 => x"00b415f1",
			1400 => x"feae15f1",
			1401 => x"03002d04",
			1402 => x"010f15f1",
			1403 => x"ff5715f1",
			1404 => x"0200f720",
			1405 => x"0e006f14",
			1406 => x"09001808",
			1407 => x"00008904",
			1408 => x"ffeb166d",
			1409 => x"0022166d",
			1410 => x"0e006a04",
			1411 => x"ffbb166d",
			1412 => x"08001d04",
			1413 => x"000b166d",
			1414 => x"fff7166d",
			1415 => x"05002a04",
			1416 => x"0094166d",
			1417 => x"01000904",
			1418 => x"0008166d",
			1419 => x"fff0166d",
			1420 => x"0600bd10",
			1421 => x"0c001704",
			1422 => x"ff7c166d",
			1423 => x"0e009104",
			1424 => x"ffe0166d",
			1425 => x"09002104",
			1426 => x"0047166d",
			1427 => x"fff8166d",
			1428 => x"03002a08",
			1429 => x"00014004",
			1430 => x"0061166d",
			1431 => x"ffe6166d",
			1432 => x"04002304",
			1433 => x"ffac166d",
			1434 => x"001a166d",
			1435 => x"09001e28",
			1436 => x"07003018",
			1437 => x"07002b0c",
			1438 => x"0e006004",
			1439 => x"cd5916e1",
			1440 => x"0000d104",
			1441 => x"e26316e1",
			1442 => x"cd5c16e1",
			1443 => x"0000f304",
			1444 => x"ed2616e1",
			1445 => x"00011f04",
			1446 => x"d1a416e1",
			1447 => x"cd5b16e1",
			1448 => x"02010004",
			1449 => x"ee7116e1",
			1450 => x"00013608",
			1451 => x"04001a04",
			1452 => x"dbb016e1",
			1453 => x"d1a416e1",
			1454 => x"cd6a16e1",
			1455 => x"09001f08",
			1456 => x"07002f04",
			1457 => x"cd5d16e1",
			1458 => x"d79d16e1",
			1459 => x"08001d08",
			1460 => x"06008a04",
			1461 => x"cd5916e1",
			1462 => x"d3bc16e1",
			1463 => x"cd5816e1",
			1464 => x"05002628",
			1465 => x"02011218",
			1466 => x"0600770c",
			1467 => x"05001a08",
			1468 => x"0a001b04",
			1469 => x"ffef1765",
			1470 => x"00211765",
			1471 => x"ffd81765",
			1472 => x"07003308",
			1473 => x"07002904",
			1474 => x"fffa1765",
			1475 => x"00801765",
			1476 => x"00011765",
			1477 => x"00013108",
			1478 => x"03002604",
			1479 => x"00111765",
			1480 => x"ffb21765",
			1481 => x"00013c04",
			1482 => x"00221765",
			1483 => x"fff21765",
			1484 => x"05002e10",
			1485 => x"0f00bf08",
			1486 => x"07003104",
			1487 => x"ffea1765",
			1488 => x"00211765",
			1489 => x"09001d04",
			1490 => x"ff971765",
			1491 => x"00031765",
			1492 => x"0f00bc04",
			1493 => x"ffd71765",
			1494 => x"0c001904",
			1495 => x"00401765",
			1496 => x"fff51765",
			1497 => x"08001c18",
			1498 => x"07002e0c",
			1499 => x"0000b708",
			1500 => x"06006b04",
			1501 => x"ffbf17d1",
			1502 => x"007117d1",
			1503 => x"ff9d17d1",
			1504 => x"00013308",
			1505 => x"0a003404",
			1506 => x"00a217d1",
			1507 => x"000817d1",
			1508 => x"ffd517d1",
			1509 => x"00011e18",
			1510 => x"0600b014",
			1511 => x"0200eb10",
			1512 => x"0e007b0c",
			1513 => x"0b001804",
			1514 => x"ff9717d1",
			1515 => x"0b001904",
			1516 => x"001417d1",
			1517 => x"ffe817d1",
			1518 => x"007217d1",
			1519 => x"ff6917d1",
			1520 => x"006917d1",
			1521 => x"03002404",
			1522 => x"002817d1",
			1523 => x"ff5017d1",
			1524 => x"06007b0c",
			1525 => x"09001808",
			1526 => x"06004c04",
			1527 => x"fe701835",
			1528 => x"022d1835",
			1529 => x"fe581835",
			1530 => x"0200f714",
			1531 => x"05003010",
			1532 => x"08001d0c",
			1533 => x"08001b08",
			1534 => x"0d001304",
			1535 => x"02f11835",
			1536 => x"02861835",
			1537 => x"03da1835",
			1538 => x"01781835",
			1539 => x"fe671835",
			1540 => x"0600b004",
			1541 => x"fe551835",
			1542 => x"0001320c",
			1543 => x"08001f08",
			1544 => x"0b001304",
			1545 => x"00ec1835",
			1546 => x"03b51835",
			1547 => x"ffc11835",
			1548 => x"fe5f1835",
			1549 => x"09001f28",
			1550 => x"07002c0c",
			1551 => x"0e006004",
			1552 => x"fe5918a9",
			1553 => x"0200ae04",
			1554 => x"045618a9",
			1555 => x"fe4f18a9",
			1556 => x"00012b14",
			1557 => x"05002c10",
			1558 => x"03002a0c",
			1559 => x"00011208",
			1560 => x"08001d04",
			1561 => x"04c418a9",
			1562 => x"03bb18a9",
			1563 => x"06fa18a9",
			1564 => x"027218a9",
			1565 => x"01d718a9",
			1566 => x"0f00e204",
			1567 => x"fe5b18a9",
			1568 => x"025c18a9",
			1569 => x"01000608",
			1570 => x"0000d004",
			1571 => x"fe6018a9",
			1572 => x"02ee18a9",
			1573 => x"0b001908",
			1574 => x"07003404",
			1575 => x"fe5a18a9",
			1576 => x"025a18a9",
			1577 => x"fe5818a9",
			1578 => x"0400191c",
			1579 => x"02011210",
			1580 => x"06006b04",
			1581 => x"ff901935",
			1582 => x"04001704",
			1583 => x"01261935",
			1584 => x"05002404",
			1585 => x"ff821935",
			1586 => x"00c61935",
			1587 => x"0f00e308",
			1588 => x"08001804",
			1589 => x"00511935",
			1590 => x"ff031935",
			1591 => x"00871935",
			1592 => x"0e008518",
			1593 => x"07003110",
			1594 => x"0300210c",
			1595 => x"03001f08",
			1596 => x"05002204",
			1597 => x"ffea1935",
			1598 => x"00031935",
			1599 => x"00121935",
			1600 => x"ff0d1935",
			1601 => x"05002d04",
			1602 => x"00391935",
			1603 => x"ffb61935",
			1604 => x"0f00c408",
			1605 => x"00011404",
			1606 => x"00f21935",
			1607 => x"ffa21935",
			1608 => x"0d001504",
			1609 => x"ff071935",
			1610 => x"01001004",
			1611 => x"00841935",
			1612 => x"ffa71935",
			1613 => x"0e009530",
			1614 => x"0000f820",
			1615 => x"0e006f14",
			1616 => x"05001f0c",
			1617 => x"05001904",
			1618 => x"ffa419b9",
			1619 => x"0e004904",
			1620 => x"ffe119b9",
			1621 => x"005119b9",
			1622 => x"04001604",
			1623 => x"000119b9",
			1624 => x"ff1119b9",
			1625 => x"05002908",
			1626 => x"0b001404",
			1627 => x"003119b9",
			1628 => x"00fa19b9",
			1629 => x"ffac19b9",
			1630 => x"04001d04",
			1631 => x"fed019b9",
			1632 => x"00010e08",
			1633 => x"06009704",
			1634 => x"ffbb19b9",
			1635 => x"00c819b9",
			1636 => x"ff4719b9",
			1637 => x"08001f0c",
			1638 => x"0b001304",
			1639 => x"ffbb19b9",
			1640 => x"03002d04",
			1641 => x"013219b9",
			1642 => x"005919b9",
			1643 => x"0f00c404",
			1644 => x"000419b9",
			1645 => x"ff4219b9",
			1646 => x"0600b028",
			1647 => x"0200eb1c",
			1648 => x"0e007b18",
			1649 => x"09001808",
			1650 => x"0e005704",
			1651 => x"ff231a25",
			1652 => x"011c1a25",
			1653 => x"0e006a04",
			1654 => x"fe831a25",
			1655 => x"03002304",
			1656 => x"01061a25",
			1657 => x"01000a04",
			1658 => x"ffeb1a25",
			1659 => x"feb31a25",
			1660 => x"016b1a25",
			1661 => x"01000608",
			1662 => x"0b001504",
			1663 => x"ff061a25",
			1664 => x"004d1a25",
			1665 => x"fe571a25",
			1666 => x"0001320c",
			1667 => x"07003304",
			1668 => x"012d1a25",
			1669 => x"0600b604",
			1670 => x"017e1a25",
			1671 => x"ff991a25",
			1672 => x"fecd1a25",
			1673 => x"0e009328",
			1674 => x"0400160c",
			1675 => x"06006b04",
			1676 => x"ffdb1a91",
			1677 => x"0000fc04",
			1678 => x"00661a91",
			1679 => x"ffe91a91",
			1680 => x"08001d18",
			1681 => x"07003010",
			1682 => x"03001d04",
			1683 => x"00091a91",
			1684 => x"0600ad08",
			1685 => x"05002204",
			1686 => x"ffff1a91",
			1687 => x"ffb61a91",
			1688 => x"fffe1a91",
			1689 => x"05002f04",
			1690 => x"00401a91",
			1691 => x"fff61a91",
			1692 => x"ff811a91",
			1693 => x"0001320c",
			1694 => x"01001008",
			1695 => x"04001a04",
			1696 => x"008c1a91",
			1697 => x"000e1a91",
			1698 => x"ffeb1a91",
			1699 => x"ffc81a91",
			1700 => x"09001b28",
			1701 => x"0d001210",
			1702 => x"0000b708",
			1703 => x"06006b04",
			1704 => x"ffba1b35",
			1705 => x"00781b35",
			1706 => x"09001a04",
			1707 => x"ff441b35",
			1708 => x"000b1b35",
			1709 => x"07002c0c",
			1710 => x"01000808",
			1711 => x"06009204",
			1712 => x"00221b35",
			1713 => x"fff31b35",
			1714 => x"ffa91b35",
			1715 => x"08001904",
			1716 => x"ffd21b35",
			1717 => x"00012e04",
			1718 => x"00f61b35",
			1719 => x"00031b35",
			1720 => x"01000b18",
			1721 => x"0700300c",
			1722 => x"03002108",
			1723 => x"05001e04",
			1724 => x"fff61b35",
			1725 => x"00091b35",
			1726 => x"ff981b35",
			1727 => x"0f00c708",
			1728 => x"03003a04",
			1729 => x"00c01b35",
			1730 => x"ffe71b35",
			1731 => x"ffb21b35",
			1732 => x"05001f08",
			1733 => x"0200a104",
			1734 => x"fff61b35",
			1735 => x"00291b35",
			1736 => x"01002108",
			1737 => x"04001604",
			1738 => x"ffec1b35",
			1739 => x"ff1f1b35",
			1740 => x"00051b35",
			1741 => x"08001c20",
			1742 => x"07002b0c",
			1743 => x"0200a908",
			1744 => x"0e005a04",
			1745 => x"ffcc1bc9",
			1746 => x"00451bc9",
			1747 => x"ffbc1bc9",
			1748 => x"00013210",
			1749 => x"0a003408",
			1750 => x"05002704",
			1751 => x"009d1bc9",
			1752 => x"00051bc9",
			1753 => x"0d001404",
			1754 => x"002c1bc9",
			1755 => x"ffc61bc9",
			1756 => x"ffd21bc9",
			1757 => x"0f00d420",
			1758 => x"0200eb14",
			1759 => x"0700300c",
			1760 => x"04001408",
			1761 => x"04001304",
			1762 => x"fffa1bc9",
			1763 => x"00061bc9",
			1764 => x"ffa71bc9",
			1765 => x"09002104",
			1766 => x"00601bc9",
			1767 => x"fff31bc9",
			1768 => x"03003404",
			1769 => x"ff521bc9",
			1770 => x"04002a04",
			1771 => x"00221bc9",
			1772 => x"fff01bc9",
			1773 => x"04001804",
			1774 => x"ffb01bc9",
			1775 => x"01001004",
			1776 => x"00851bc9",
			1777 => x"ffe61bc9",
			1778 => x"09001f30",
			1779 => x"07002c10",
			1780 => x"0e006004",
			1781 => x"fe571c3d",
			1782 => x"0200ae04",
			1783 => x"06df1c3d",
			1784 => x"05001f04",
			1785 => x"00411c3d",
			1786 => x"fe4f1c3d",
			1787 => x"00011e14",
			1788 => x"0600b010",
			1789 => x"0000f80c",
			1790 => x"0f009304",
			1791 => x"04d41c3d",
			1792 => x"0f00a004",
			1793 => x"06d31c3d",
			1794 => x"05d71c3d",
			1795 => x"01551c3d",
			1796 => x"079c1c3d",
			1797 => x"0e00a508",
			1798 => x"03003104",
			1799 => x"fe581c3d",
			1800 => x"00661c3d",
			1801 => x"066a1c3d",
			1802 => x"08001d08",
			1803 => x"07003504",
			1804 => x"fe571c3d",
			1805 => x"03b91c3d",
			1806 => x"fe561c3d",
			1807 => x"0e008520",
			1808 => x"04001910",
			1809 => x"06006b04",
			1810 => x"ffc71cc1",
			1811 => x"0000f408",
			1812 => x"01000804",
			1813 => x"00641cc1",
			1814 => x"fff11cc1",
			1815 => x"ffda1cc1",
			1816 => x"0300210c",
			1817 => x"03001c04",
			1818 => x"fff81cc1",
			1819 => x"05002304",
			1820 => x"00111cc1",
			1821 => x"fff91cc1",
			1822 => x"ff811cc1",
			1823 => x"00013220",
			1824 => x"03002a0c",
			1825 => x"0e009308",
			1826 => x"0000f804",
			1827 => x"005e1cc1",
			1828 => x"ffc81cc1",
			1829 => x"00a21cc1",
			1830 => x"0e00a010",
			1831 => x"03002f08",
			1832 => x"0f00c104",
			1833 => x"00351cc1",
			1834 => x"ffbc1cc1",
			1835 => x"0600b004",
			1836 => x"ffea1cc1",
			1837 => x"00a91cc1",
			1838 => x"ffa51cc1",
			1839 => x"ff9e1cc1",
			1840 => x"0e008524",
			1841 => x"0900180c",
			1842 => x"07002504",
			1843 => x"ffdd1d4d",
			1844 => x"0000fc04",
			1845 => x"003d1d4d",
			1846 => x"fff81d4d",
			1847 => x"0700300c",
			1848 => x"08001504",
			1849 => x"00031d4d",
			1850 => x"01000204",
			1851 => x"00021d4d",
			1852 => x"ffa31d4d",
			1853 => x"08001d08",
			1854 => x"07003304",
			1855 => x"00131d4d",
			1856 => x"ffff1d4d",
			1857 => x"ffef1d4d",
			1858 => x"00013220",
			1859 => x"03002a0c",
			1860 => x"01000c08",
			1861 => x"0200f104",
			1862 => x"ffec1d4d",
			1863 => x"001a1d4d",
			1864 => x"00891d4d",
			1865 => x"08001c04",
			1866 => x"00401d4d",
			1867 => x"03002f08",
			1868 => x"0600ae04",
			1869 => x"00101d4d",
			1870 => x"ffa21d4d",
			1871 => x"00011b04",
			1872 => x"002f1d4d",
			1873 => x"ffdd1d4d",
			1874 => x"ffc11d4d",
			1875 => x"0e008524",
			1876 => x"04001910",
			1877 => x"06006b04",
			1878 => x"fea21dd1",
			1879 => x"0000e908",
			1880 => x"0b001404",
			1881 => x"01411dd1",
			1882 => x"00341dd1",
			1883 => x"fed21dd1",
			1884 => x"0700300c",
			1885 => x"03002108",
			1886 => x"0a002104",
			1887 => x"ff4b1dd1",
			1888 => x"00411dd1",
			1889 => x"fe661dd1",
			1890 => x"05002904",
			1891 => x"00e51dd1",
			1892 => x"fecd1dd1",
			1893 => x"0001321c",
			1894 => x"03002604",
			1895 => x"018f1dd1",
			1896 => x"08001c08",
			1897 => x"0b001404",
			1898 => x"01731dd1",
			1899 => x"00d31dd1",
			1900 => x"0d001504",
			1901 => x"ff2a1dd1",
			1902 => x"00011e08",
			1903 => x"0a003604",
			1904 => x"016c1dd1",
			1905 => x"fef41dd1",
			1906 => x"feb41dd1",
			1907 => x"fe911dd1",
			1908 => x"08001c1c",
			1909 => x"06006b04",
			1910 => x"ffe11e4d",
			1911 => x"00013214",
			1912 => x"05004010",
			1913 => x"0d001004",
			1914 => x"fffc1e4d",
			1915 => x"01000a04",
			1916 => x"00671e4d",
			1917 => x"01000c04",
			1918 => x"ffef1e4d",
			1919 => x"00271e4d",
			1920 => x"fffa1e4d",
			1921 => x"ffe61e4d",
			1922 => x"03002608",
			1923 => x"0e008604",
			1924 => x"ffd21e4d",
			1925 => x"00451e4d",
			1926 => x"0000f708",
			1927 => x"05002a04",
			1928 => x"00241e4d",
			1929 => x"fff01e4d",
			1930 => x"0400230c",
			1931 => x"07003808",
			1932 => x"0d001804",
			1933 => x"ff7c1e4d",
			1934 => x"00011e4d",
			1935 => x"00151e4d",
			1936 => x"0c001904",
			1937 => x"00241e4d",
			1938 => x"ffea1e4d",
			1939 => x"04001928",
			1940 => x"0700331c",
			1941 => x"0700290c",
			1942 => x"02009008",
			1943 => x"00008904",
			1944 => x"ffe31ef1",
			1945 => x"00371ef1",
			1946 => x"ffc51ef1",
			1947 => x"00011d08",
			1948 => x"09001f04",
			1949 => x"00ad1ef1",
			1950 => x"fffb1ef1",
			1951 => x"00013104",
			1952 => x"ffbf1ef1",
			1953 => x"00341ef1",
			1954 => x"07003508",
			1955 => x"08001f04",
			1956 => x"ff911ef1",
			1957 => x"00071ef1",
			1958 => x"004e1ef1",
			1959 => x"04002320",
			1960 => x"00010114",
			1961 => x"0e007d10",
			1962 => x"0b00180c",
			1963 => x"03002108",
			1964 => x"03001e04",
			1965 => x"ffff1ef1",
			1966 => x"00011ef1",
			1967 => x"ffbe1ef1",
			1968 => x"00031ef1",
			1969 => x"00571ef1",
			1970 => x"07003904",
			1971 => x"ff6a1ef1",
			1972 => x"07003b04",
			1973 => x"00031ef1",
			1974 => x"fffc1ef1",
			1975 => x"0e009104",
			1976 => x"ffbd1ef1",
			1977 => x"00012704",
			1978 => x"00531ef1",
			1979 => x"fff11ef1",
			1980 => x"09001f30",
			1981 => x"07002e14",
			1982 => x"05002410",
			1983 => x"0e006304",
			1984 => x"fe591f65",
			1985 => x"0000e908",
			1986 => x"0e007204",
			1987 => x"02841f65",
			1988 => x"031d1f65",
			1989 => x"fe6b1f65",
			1990 => x"fe561f65",
			1991 => x"00013218",
			1992 => x"0c001814",
			1993 => x"03002a0c",
			1994 => x"0f00c308",
			1995 => x"08001c04",
			1996 => x"03231f65",
			1997 => x"01f01f65",
			1998 => x"04301f65",
			1999 => x"0e00a004",
			2000 => x"02731f65",
			2001 => x"ff781f65",
			2002 => x"04381f65",
			2003 => x"fe641f65",
			2004 => x"08001d08",
			2005 => x"06008e04",
			2006 => x"fe5d1f65",
			2007 => x"044c1f65",
			2008 => x"fe5c1f65",
			2009 => x"08001c28",
			2010 => x"0d00141c",
			2011 => x"07002e10",
			2012 => x"0000b708",
			2013 => x"06006b04",
			2014 => x"ffc12019",
			2015 => x"007e2019",
			2016 => x"0b001504",
			2017 => x"ff8f2019",
			2018 => x"00052019",
			2019 => x"00013308",
			2020 => x"0d001204",
			2021 => x"00282019",
			2022 => x"00c12019",
			2023 => x"ffdc2019",
			2024 => x"00010308",
			2025 => x"0f008d04",
			2026 => x"ffe32019",
			2027 => x"00222019",
			2028 => x"ff9f2019",
			2029 => x"0e009e20",
			2030 => x"0b001308",
			2031 => x"04001804",
			2032 => x"fff72019",
			2033 => x"00362019",
			2034 => x"0200eb0c",
			2035 => x"0000bc04",
			2036 => x"ffa62019",
			2037 => x"04002304",
			2038 => x"00662019",
			2039 => x"ffeb2019",
			2040 => x"03003404",
			2041 => x"ff2c2019",
			2042 => x"04002b04",
			2043 => x"001a2019",
			2044 => x"ffe82019",
			2045 => x"0f00dd0c",
			2046 => x"0f00d404",
			2047 => x"ffe02019",
			2048 => x"0a003604",
			2049 => x"00a62019",
			2050 => x"fff62019",
			2051 => x"03002c04",
			2052 => x"fff62019",
			2053 => x"ff912019",
			2054 => x"0600770c",
			2055 => x"09001708",
			2056 => x"0d001004",
			2057 => x"fe9220a5",
			2058 => x"014e20a5",
			2059 => x"fe5f20a5",
			2060 => x"00011628",
			2061 => x"08001c14",
			2062 => x"07002904",
			2063 => x"fe9520a5",
			2064 => x"0a00340c",
			2065 => x"0e008508",
			2066 => x"0000cc04",
			2067 => x"01e320a5",
			2068 => x"00f020a5",
			2069 => x"02a320a5",
			2070 => x"ffba20a5",
			2071 => x"0e008008",
			2072 => x"01000a04",
			2073 => x"ffc220a5",
			2074 => x"fe3520a5",
			2075 => x"0200ec04",
			2076 => x"020b20a5",
			2077 => x"03002f04",
			2078 => x"feff20a5",
			2079 => x"026b20a5",
			2080 => x"0f00e30c",
			2081 => x"04001808",
			2082 => x"0b001304",
			2083 => x"fe3020a5",
			2084 => x"00ac20a5",
			2085 => x"fe6020a5",
			2086 => x"02014504",
			2087 => x"024920a5",
			2088 => x"fe8c20a5",
			2089 => x"07002e18",
			2090 => x"01000814",
			2091 => x"05002310",
			2092 => x"0a002004",
			2093 => x"ffb22131",
			2094 => x"0000ca08",
			2095 => x"02008c04",
			2096 => x"fffc2131",
			2097 => x"009c2131",
			2098 => x"fff12131",
			2099 => x"ff6e2131",
			2100 => x"ff0c2131",
			2101 => x"08001c10",
			2102 => x"00011d08",
			2103 => x"09002004",
			2104 => x"011d2131",
			2105 => x"ffe72131",
			2106 => x"03002904",
			2107 => x"ff942131",
			2108 => x"00a92131",
			2109 => x"0d001404",
			2110 => x"ff212131",
			2111 => x"03002a0c",
			2112 => x"09001e04",
			2113 => x"012a2131",
			2114 => x"01000e04",
			2115 => x"00132131",
			2116 => x"ff972131",
			2117 => x"03002f08",
			2118 => x"0f00bf04",
			2119 => x"00102131",
			2120 => x"ff0a2131",
			2121 => x"09002004",
			2122 => x"00972131",
			2123 => x"ff722131",
			2124 => x"0e00852c",
			2125 => x"04001914",
			2126 => x"0e00680c",
			2127 => x"09001808",
			2128 => x"03001504",
			2129 => x"ff4321c5",
			2130 => x"011621c5",
			2131 => x"fe7921c5",
			2132 => x"0000e904",
			2133 => x"017121c5",
			2134 => x"fedc21c5",
			2135 => x"07003010",
			2136 => x"0300210c",
			2137 => x"05002308",
			2138 => x"0a001c04",
			2139 => x"ff7021c5",
			2140 => x"00a921c5",
			2141 => x"ff5521c5",
			2142 => x"fe6b21c5",
			2143 => x"05002904",
			2144 => x"00d821c5",
			2145 => x"fed821c5",
			2146 => x"0001321c",
			2147 => x"03002604",
			2148 => x"018221c5",
			2149 => x"08001c08",
			2150 => x"0b001404",
			2151 => x"015e21c5",
			2152 => x"00c421c5",
			2153 => x"0d001504",
			2154 => x"ff3c21c5",
			2155 => x"01001004",
			2156 => x"013621c5",
			2157 => x"00011904",
			2158 => x"007121c5",
			2159 => x"feaf21c5",
			2160 => x"fe9721c5",
			2161 => x"09002028",
			2162 => x"0e006004",
			2163 => x"fe732229",
			2164 => x"00013220",
			2165 => x"05002108",
			2166 => x"0200f204",
			2167 => x"01ad2229",
			2168 => x"00d02229",
			2169 => x"07002e08",
			2170 => x"0000c704",
			2171 => x"fff92229",
			2172 => x"fe662229",
			2173 => x"08001c08",
			2174 => x"00011d04",
			2175 => x"020f2229",
			2176 => x"00de2229",
			2177 => x"0d001604",
			2178 => x"001b2229",
			2179 => x"017d2229",
			2180 => x"fe762229",
			2181 => x"01000a08",
			2182 => x"07003504",
			2183 => x"fe802229",
			2184 => x"01072229",
			2185 => x"fe6b2229",
			2186 => x"0e008520",
			2187 => x"01000b1c",
			2188 => x"05002918",
			2189 => x"0700290c",
			2190 => x"05001a08",
			2191 => x"0a001b04",
			2192 => x"feb7229d",
			2193 => x"0170229d",
			2194 => x"fe5a229d",
			2195 => x"00010408",
			2196 => x"06007704",
			2197 => x"ff11229d",
			2198 => x"019e229d",
			2199 => x"feba229d",
			2200 => x"fe7e229d",
			2201 => x"fe5c229d",
			2202 => x"00013218",
			2203 => x"03002604",
			2204 => x"01a2229d",
			2205 => x"08001c04",
			2206 => x"011c229d",
			2207 => x"0d001504",
			2208 => x"ff32229d",
			2209 => x"02011308",
			2210 => x"0a003604",
			2211 => x"01cf229d",
			2212 => x"fed5229d",
			2213 => x"fe93229d",
			2214 => x"fe7d229d",
			2215 => x"0600ca3c",
			2216 => x"00011e2c",
			2217 => x"0400160c",
			2218 => x"06006b04",
			2219 => x"ff7d2321",
			2220 => x"01000904",
			2221 => x"005a2321",
			2222 => x"012b2321",
			2223 => x"0e008314",
			2224 => x"05001f08",
			2225 => x"04001904",
			2226 => x"00572321",
			2227 => x"fff62321",
			2228 => x"07003004",
			2229 => x"fef62321",
			2230 => x"0b001904",
			2231 => x"00592321",
			2232 => x"ff9e2321",
			2233 => x"0d001504",
			2234 => x"ffbc2321",
			2235 => x"0a003604",
			2236 => x"00ed2321",
			2237 => x"ffa92321",
			2238 => x"0d001108",
			2239 => x"05002e04",
			2240 => x"ffbf2321",
			2241 => x"009f2321",
			2242 => x"05002204",
			2243 => x"ffe72321",
			2244 => x"feba2321",
			2245 => x"03002d04",
			2246 => x"00e62321",
			2247 => x"ffae2321",
			2248 => x"0e009540",
			2249 => x"0200eb24",
			2250 => x"0e007218",
			2251 => x"0900180c",
			2252 => x"0d001004",
			2253 => x"ffdc23c5",
			2254 => x"03001504",
			2255 => x"fff823c5",
			2256 => x"005823c5",
			2257 => x"0d001104",
			2258 => x"000923c5",
			2259 => x"08001604",
			2260 => x"000423c5",
			2261 => x"ff7123c5",
			2262 => x"05002d08",
			2263 => x"06008604",
			2264 => x"001223c5",
			2265 => x"00aa23c5",
			2266 => x"ffe923c5",
			2267 => x"04001d04",
			2268 => x"ff2c23c5",
			2269 => x"0600b010",
			2270 => x"08001c0c",
			2271 => x"0f00bd08",
			2272 => x"06009704",
			2273 => x"fff123c5",
			2274 => x"003a23c5",
			2275 => x"ffec23c5",
			2276 => x"ff9b23c5",
			2277 => x"0600b304",
			2278 => x"005223c5",
			2279 => x"fff723c5",
			2280 => x"08001f0c",
			2281 => x"00011f04",
			2282 => x"00bd23c5",
			2283 => x"0f00e304",
			2284 => x"ff8623c5",
			2285 => x"006323c5",
			2286 => x"0f00c504",
			2287 => x"000323c5",
			2288 => x"ff9223c5",
			2289 => x"09001f30",
			2290 => x"0700290c",
			2291 => x"09001808",
			2292 => x"07002504",
			2293 => x"fe6b2439",
			2294 => x"01f82439",
			2295 => x"fe562439",
			2296 => x"00013220",
			2297 => x"0a00361c",
			2298 => x"0400190c",
			2299 => x"0b001304",
			2300 => x"01572439",
			2301 => x"0f00c604",
			2302 => x"02632439",
			2303 => x"04062439",
			2304 => x"07003008",
			2305 => x"09001b04",
			2306 => x"00e02439",
			2307 => x"fe0b2439",
			2308 => x"0e009404",
			2309 => x"02e32439",
			2310 => x"00fd2439",
			2311 => x"fe602439",
			2312 => x"fe632439",
			2313 => x"08001d08",
			2314 => x"07003504",
			2315 => x"fe602439",
			2316 => x"030d2439",
			2317 => x"fe5f2439",
			2318 => x"09001f3c",
			2319 => x"07002c18",
			2320 => x"04001910",
			2321 => x"06006b04",
			2322 => x"fe6824c5",
			2323 => x"0000b704",
			2324 => x"024224c5",
			2325 => x"09001904",
			2326 => x"fe4f24c5",
			2327 => x"000424c5",
			2328 => x"03001d04",
			2329 => x"fff324c5",
			2330 => x"fe4a24c5",
			2331 => x"00013220",
			2332 => x"03002a14",
			2333 => x"08001d0c",
			2334 => x"0e008d08",
			2335 => x"0f00a904",
			2336 => x"023324c5",
			2337 => x"00e324c5",
			2338 => x"02ce24c5",
			2339 => x"07003004",
			2340 => x"fed224c5",
			2341 => x"01eb24c5",
			2342 => x"0d001304",
			2343 => x"fe2124c5",
			2344 => x"00011f04",
			2345 => x"01c824c5",
			2346 => x"ffa224c5",
			2347 => x"fe6824c5",
			2348 => x"09002108",
			2349 => x"07003404",
			2350 => x"fe6424c5",
			2351 => x"022d24c5",
			2352 => x"fe6124c5",
			2353 => x"0f007a0c",
			2354 => x"0b001208",
			2355 => x"0b001004",
			2356 => x"feaa2551",
			2357 => x"00d22551",
			2358 => x"fe642551",
			2359 => x"00011e28",
			2360 => x"05004024",
			2361 => x"0400170c",
			2362 => x"0c001404",
			2363 => x"02632551",
			2364 => x"0000e904",
			2365 => x"01cb2551",
			2366 => x"01242551",
			2367 => x"0700300c",
			2368 => x"0d001408",
			2369 => x"00010104",
			2370 => x"01782551",
			2371 => x"fe7b2551",
			2372 => x"fe442551",
			2373 => x"01000a04",
			2374 => x"02442551",
			2375 => x"0d001504",
			2376 => x"00082551",
			2377 => x"01ae2551",
			2378 => x"fe722551",
			2379 => x"0600c90c",
			2380 => x"0d001108",
			2381 => x"05002e04",
			2382 => x"fe942551",
			2383 => x"01972551",
			2384 => x"fe5b2551",
			2385 => x"03002a04",
			2386 => x"01bb2551",
			2387 => x"fe592551",
			2388 => x"0e009334",
			2389 => x"00010a30",
			2390 => x"08001d1c",
			2391 => x"0e006b10",
			2392 => x"09001808",
			2393 => x"0a001c04",
			2394 => x"ffb925f5",
			2395 => x"008f25f5",
			2396 => x"0d001104",
			2397 => x"000125f5",
			2398 => x"ff2d25f5",
			2399 => x"03003108",
			2400 => x"07002c04",
			2401 => x"002525f5",
			2402 => x"011925f5",
			2403 => x"ffce25f5",
			2404 => x"04001608",
			2405 => x"0200aa04",
			2406 => x"ffe125f5",
			2407 => x"007425f5",
			2408 => x"04002004",
			2409 => x"ff0025f5",
			2410 => x"04002204",
			2411 => x"001325f5",
			2412 => x"ffa625f5",
			2413 => x"fef125f5",
			2414 => x"03002f14",
			2415 => x"03002d10",
			2416 => x"0600ca0c",
			2417 => x"00011f04",
			2418 => x"00a525f5",
			2419 => x"0a002d04",
			2420 => x"fffc25f5",
			2421 => x"feee25f5",
			2422 => x"00d925f5",
			2423 => x"fefd25f5",
			2424 => x"0e00a008",
			2425 => x"00012e04",
			2426 => x"012925f5",
			2427 => x"ffe325f5",
			2428 => x"ff9d25f5",
			2429 => x"0e006a0c",
			2430 => x"09001808",
			2431 => x"00008804",
			2432 => x"feb32661",
			2433 => x"011d2661",
			2434 => x"fe642661",
			2435 => x"00013228",
			2436 => x"09002224",
			2437 => x"00011e14",
			2438 => x"0e009510",
			2439 => x"08001d08",
			2440 => x"00010a04",
			2441 => x"015c2661",
			2442 => x"fe852661",
			2443 => x"0000f504",
			2444 => x"00222661",
			2445 => x"fdc62661",
			2446 => x"018f2661",
			2447 => x"0201230c",
			2448 => x"04001704",
			2449 => x"fe492661",
			2450 => x"04001d04",
			2451 => x"01172661",
			2452 => x"fe972661",
			2453 => x"016e2661",
			2454 => x"fe822661",
			2455 => x"fe732661",
			2456 => x"0e009640",
			2457 => x"0500200c",
			2458 => x"06006b04",
			2459 => x"ffe626fd",
			2460 => x"0000fc04",
			2461 => x"003a26fd",
			2462 => x"fffb26fd",
			2463 => x"0900190c",
			2464 => x"00010308",
			2465 => x"06005d04",
			2466 => x"fffc26fd",
			2467 => x"002b26fd",
			2468 => x"ffe226fd",
			2469 => x"07003418",
			2470 => x"0800180c",
			2471 => x"08001604",
			2472 => x"fff926fd",
			2473 => x"0c001704",
			2474 => x"000026fd",
			2475 => x"000b26fd",
			2476 => x"0c001404",
			2477 => x"ffff26fd",
			2478 => x"0c001904",
			2479 => x"ff8a26fd",
			2480 => x"fffb26fd",
			2481 => x"01000b08",
			2482 => x"06009004",
			2483 => x"000026fd",
			2484 => x"002426fd",
			2485 => x"08002004",
			2486 => x"000226fd",
			2487 => x"ffe326fd",
			2488 => x"0b001304",
			2489 => x"ffdc26fd",
			2490 => x"01001008",
			2491 => x"01000c04",
			2492 => x"000a26fd",
			2493 => x"007b26fd",
			2494 => x"ffe326fd",
			2495 => x"0900204c",
			2496 => x"07002e2c",
			2497 => x"05002014",
			2498 => x"0600700c",
			2499 => x"0b001208",
			2500 => x"05001604",
			2501 => x"ff3327a9",
			2502 => x"010327a9",
			2503 => x"fe6c27a9",
			2504 => x"0000fc04",
			2505 => x"016b27a9",
			2506 => x"feeb27a9",
			2507 => x"04001608",
			2508 => x"0f00b804",
			2509 => x"00c527a9",
			2510 => x"fef827a9",
			2511 => x"07002c08",
			2512 => x"08001504",
			2513 => x"ff8627a9",
			2514 => x"fe6a27a9",
			2515 => x"05002804",
			2516 => x"000b27a9",
			2517 => x"fec627a9",
			2518 => x"0001321c",
			2519 => x"01000a08",
			2520 => x"07003304",
			2521 => x"00d627a9",
			2522 => x"01bf27a9",
			2523 => x"0d00150c",
			2524 => x"08001d08",
			2525 => x"00010604",
			2526 => x"01a927a9",
			2527 => x"003227a9",
			2528 => x"ff0a27a9",
			2529 => x"0e008604",
			2530 => x"fec127a9",
			2531 => x"015d27a9",
			2532 => x"fea827a9",
			2533 => x"01000608",
			2534 => x"04001e04",
			2535 => x"00eb27a9",
			2536 => x"fef627a9",
			2537 => x"fe7327a9",
			2538 => x"0600bd3c",
			2539 => x"0f00c830",
			2540 => x"0600b02c",
			2541 => x"0000f820",
			2542 => x"0e006f10",
			2543 => x"09001808",
			2544 => x"0a001c04",
			2545 => x"ffdf282f",
			2546 => x"003b282f",
			2547 => x"01000204",
			2548 => x"0003282f",
			2549 => x"ff90282f",
			2550 => x"05002a08",
			2551 => x"0000bc04",
			2552 => x"000b282f",
			2553 => x"0083282f",
			2554 => x"08002004",
			2555 => x"0002282f",
			2556 => x"fff1282f",
			2557 => x"07003504",
			2558 => x"ff75282f",
			2559 => x"08001f04",
			2560 => x"001f282f",
			2561 => x"ffe0282f",
			2562 => x"0087282f",
			2563 => x"07003804",
			2564 => x"ff78282f",
			2565 => x"0e009f04",
			2566 => x"fff7282f",
			2567 => x"000f282f",
			2568 => x"00013304",
			2569 => x"0080282f",
			2570 => x"ffc6282f",
			2571 => x"03002a20",
			2572 => x"0e009318",
			2573 => x"0000eb10",
			2574 => x"0e00680c",
			2575 => x"05001a08",
			2576 => x"07002504",
			2577 => x"ffe22891",
			2578 => x"00342891",
			2579 => x"ffb82891",
			2580 => x"006e2891",
			2581 => x"03002904",
			2582 => x"ff922891",
			2583 => x"00132891",
			2584 => x"00013404",
			2585 => x"007f2891",
			2586 => x"ffd82891",
			2587 => x"0200f608",
			2588 => x"0e007a04",
			2589 => x"ffd92891",
			2590 => x"005a2891",
			2591 => x"04002304",
			2592 => x"ff402891",
			2593 => x"09002004",
			2594 => x"003b2891",
			2595 => x"ffde2891",
			2596 => x"08001c14",
			2597 => x"00013210",
			2598 => x"0f007404",
			2599 => x"ffe928f5",
			2600 => x"04003108",
			2601 => x"0d001004",
			2602 => x"fffe28f5",
			2603 => x"005e28f5",
			2604 => x"fffc28f5",
			2605 => x"ffe928f5",
			2606 => x"0d001510",
			2607 => x"03002608",
			2608 => x"0a002a04",
			2609 => x"ffe128f5",
			2610 => x"002d28f5",
			2611 => x"0b001704",
			2612 => x"ff9d28f5",
			2613 => x"000928f5",
			2614 => x"00011e0c",
			2615 => x"0e008604",
			2616 => x"ffe228f5",
			2617 => x"01001204",
			2618 => x"005228f5",
			2619 => x"fff528f5",
			2620 => x"ffdb28f5",
			2621 => x"0e008524",
			2622 => x"05001f0c",
			2623 => x"0f007404",
			2624 => x"ffc82969",
			2625 => x"0000b704",
			2626 => x"006b2969",
			2627 => x"ffe32969",
			2628 => x"04001608",
			2629 => x"07002a04",
			2630 => x"fff62969",
			2631 => x"001d2969",
			2632 => x"07003008",
			2633 => x"03001d04",
			2634 => x"00012969",
			2635 => x"ff662969",
			2636 => x"0b001904",
			2637 => x"00222969",
			2638 => x"ffde2969",
			2639 => x"02011308",
			2640 => x"0d001904",
			2641 => x"00852969",
			2642 => x"ffe62969",
			2643 => x"0600ca08",
			2644 => x"08001804",
			2645 => x"002a2969",
			2646 => x"ff4e2969",
			2647 => x"03002d04",
			2648 => x"00802969",
			2649 => x"ffb82969",
			2650 => x"00010320",
			2651 => x"0e007b18",
			2652 => x"0400190c",
			2653 => x"06006b04",
			2654 => x"ffe829dd",
			2655 => x"0000b504",
			2656 => x"003129dd",
			2657 => x"fff929dd",
			2658 => x"03002108",
			2659 => x"03001f04",
			2660 => x"fffe29dd",
			2661 => x"000429dd",
			2662 => x"ffc829dd",
			2663 => x"01000904",
			2664 => x"fffe29dd",
			2665 => x"006829dd",
			2666 => x"0e00a514",
			2667 => x"03002f0c",
			2668 => x"04002508",
			2669 => x"07003904",
			2670 => x"ff7c29dd",
			2671 => x"000229dd",
			2672 => x"000529dd",
			2673 => x"09002004",
			2674 => x"004429dd",
			2675 => x"ffee29dd",
			2676 => x"03002d04",
			2677 => x"003a29dd",
			2678 => x"ffdd29dd",
			2679 => x"0e009428",
			2680 => x"0000f310",
			2681 => x"0f007404",
			2682 => x"ffc42a49",
			2683 => x"05002a08",
			2684 => x"01000b04",
			2685 => x"00812a49",
			2686 => x"fffb2a49",
			2687 => x"ffe52a49",
			2688 => x"0400250c",
			2689 => x"07003604",
			2690 => x"ff7c2a49",
			2691 => x"07003a04",
			2692 => x"00042a49",
			2693 => x"fff92a49",
			2694 => x"0c001908",
			2695 => x"04002904",
			2696 => x"001b2a49",
			2697 => x"fffb2a49",
			2698 => x"ffeb2a49",
			2699 => x"0001320c",
			2700 => x"08001f08",
			2701 => x"03002a04",
			2702 => x"00892a49",
			2703 => x"00172a49",
			2704 => x"ffe02a49",
			2705 => x"ffcd2a49",
			2706 => x"08001c1c",
			2707 => x"06006b04",
			2708 => x"ffde2abd",
			2709 => x"0d00140c",
			2710 => x"00013208",
			2711 => x"0d001004",
			2712 => x"fffb2abd",
			2713 => x"00632abd",
			2714 => x"ffe92abd",
			2715 => x"00010308",
			2716 => x"0f008d04",
			2717 => x"fff92abd",
			2718 => x"000e2abd",
			2719 => x"ffdc2abd",
			2720 => x"0d001510",
			2721 => x"03002608",
			2722 => x"0600a804",
			2723 => x"ffda2abd",
			2724 => x"00312abd",
			2725 => x"0000f804",
			2726 => x"00152abd",
			2727 => x"ff8a2abd",
			2728 => x"09001f0c",
			2729 => x"00012008",
			2730 => x"0e008604",
			2731 => x"fff32abd",
			2732 => x"005e2abd",
			2733 => x"ffe82abd",
			2734 => x"ffd62abd",
			2735 => x"08001c18",
			2736 => x"07002e0c",
			2737 => x"0000b708",
			2738 => x"06006b04",
			2739 => x"ffc22b29",
			2740 => x"006e2b29",
			2741 => x"ffa12b29",
			2742 => x"00013308",
			2743 => x"0a003404",
			2744 => x"009a2b29",
			2745 => x"00082b29",
			2746 => x"ffd62b29",
			2747 => x"00011e18",
			2748 => x"0600b014",
			2749 => x"0200eb10",
			2750 => x"0e007b0c",
			2751 => x"0b001804",
			2752 => x"ff9b2b29",
			2753 => x"0b001904",
			2754 => x"00132b29",
			2755 => x"ffe92b29",
			2756 => x"006e2b29",
			2757 => x"ff6f2b29",
			2758 => x"00632b29",
			2759 => x"03002404",
			2760 => x"00282b29",
			2761 => x"ff562b29",
			2762 => x"0e006f14",
			2763 => x"0b001308",
			2764 => x"07002104",
			2765 => x"fe8a2b8d",
			2766 => x"01462b8d",
			2767 => x"0e006c04",
			2768 => x"fe5e2b8d",
			2769 => x"01000b04",
			2770 => x"00bc2b8d",
			2771 => x"fe702b8d",
			2772 => x"0001321c",
			2773 => x"09002218",
			2774 => x"0200f70c",
			2775 => x"0e007c08",
			2776 => x"04001904",
			2777 => x"01ac2b8d",
			2778 => x"ff362b8d",
			2779 => x"01df2b8d",
			2780 => x"0e009104",
			2781 => x"fe6a2b8d",
			2782 => x"03002a04",
			2783 => x"01d92b8d",
			2784 => x"00752b8d",
			2785 => x"fe772b8d",
			2786 => x"fe6c2b8d",
			2787 => x"09001f2c",
			2788 => x"07002e14",
			2789 => x"0000b710",
			2790 => x"01000808",
			2791 => x"06006b04",
			2792 => x"fec92c01",
			2793 => x"01942c01",
			2794 => x"08001904",
			2795 => x"ffe72c01",
			2796 => x"fe922c01",
			2797 => x"fe902c01",
			2798 => x"00011e10",
			2799 => x"04001804",
			2800 => x"01c72c01",
			2801 => x"0d001508",
			2802 => x"04001d04",
			2803 => x"ff252c01",
			2804 => x"01012c01",
			2805 => x"012d2c01",
			2806 => x"0600c904",
			2807 => x"fe692c01",
			2808 => x"00762c01",
			2809 => x"0100060c",
			2810 => x"04002608",
			2811 => x"04000d04",
			2812 => x"ffc72c01",
			2813 => x"01122c01",
			2814 => x"fef82c01",
			2815 => x"fe782c01",
			2816 => x"0700301c",
			2817 => x"09001b18",
			2818 => x"00010314",
			2819 => x"0700290c",
			2820 => x"05001a08",
			2821 => x"02006b04",
			2822 => x"ff582c75",
			2823 => x"01282c75",
			2824 => x"fe912c75",
			2825 => x"07002c04",
			2826 => x"00b82c75",
			2827 => x"01742c75",
			2828 => x"fe902c75",
			2829 => x"fe882c75",
			2830 => x"0200f708",
			2831 => x"09002204",
			2832 => x"01892c75",
			2833 => x"fefc2c75",
			2834 => x"08001f10",
			2835 => x"01000c08",
			2836 => x"01000a04",
			2837 => x"00902c75",
			2838 => x"fe702c75",
			2839 => x"0e009e04",
			2840 => x"ffd12c75",
			2841 => x"011f2c75",
			2842 => x"00010e04",
			2843 => x"00d22c75",
			2844 => x"fe802c75",
			2845 => x"03002a2c",
			2846 => x"0e009320",
			2847 => x"0000eb14",
			2848 => x"0e006a0c",
			2849 => x"09001808",
			2850 => x"0a001b04",
			2851 => x"ffcc2d09",
			2852 => x"00692d09",
			2853 => x"ff682d09",
			2854 => x"09001c04",
			2855 => x"00a22d09",
			2856 => x"00052d09",
			2857 => x"0a002f04",
			2858 => x"ff492d09",
			2859 => x"0a003104",
			2860 => x"00462d09",
			2861 => x"ffe32d09",
			2862 => x"08001f08",
			2863 => x"00013404",
			2864 => x"00b82d09",
			2865 => x"ffd12d09",
			2866 => x"ffca2d09",
			2867 => x"09001c10",
			2868 => x"00013108",
			2869 => x"0000e704",
			2870 => x"00032d09",
			2871 => x"ff022d09",
			2872 => x"00013904",
			2873 => x"005a2d09",
			2874 => x"ffec2d09",
			2875 => x"0e009308",
			2876 => x"05002e04",
			2877 => x"002c2d09",
			2878 => x"ff6b2d09",
			2879 => x"00012a04",
			2880 => x"00bb2d09",
			2881 => x"ffd32d09",
			2882 => x"0600b028",
			2883 => x"0200eb1c",
			2884 => x"0e007b18",
			2885 => x"09001808",
			2886 => x"0e005704",
			2887 => x"ff2e2d75",
			2888 => x"010c2d75",
			2889 => x"0e006a04",
			2890 => x"fe892d75",
			2891 => x"03002304",
			2892 => x"00f72d75",
			2893 => x"01000a04",
			2894 => x"ffeb2d75",
			2895 => x"fec12d75",
			2896 => x"01642d75",
			2897 => x"08001808",
			2898 => x"04002204",
			2899 => x"ff192d75",
			2900 => x"009b2d75",
			2901 => x"fe662d75",
			2902 => x"0001320c",
			2903 => x"07003304",
			2904 => x"010f2d75",
			2905 => x"0600b604",
			2906 => x"01762d75",
			2907 => x"ffa92d75",
			2908 => x"fed72d75",
			2909 => x"0500262c",
			2910 => x"0201121c",
			2911 => x"0700290c",
			2912 => x"05001a08",
			2913 => x"07002504",
			2914 => x"ffef2e11",
			2915 => x"00232e11",
			2916 => x"ffd62e11",
			2917 => x"07003308",
			2918 => x"06007704",
			2919 => x"fffb2e11",
			2920 => x"00852e11",
			2921 => x"07003404",
			2922 => x"ffe82e11",
			2923 => x"00172e11",
			2924 => x"00013108",
			2925 => x"03002604",
			2926 => x"00112e11",
			2927 => x"ffb02e11",
			2928 => x"00013c04",
			2929 => x"00232e11",
			2930 => x"fff22e11",
			2931 => x"05002e18",
			2932 => x"0f00bf10",
			2933 => x"06008e08",
			2934 => x"0b001704",
			2935 => x"fff32e11",
			2936 => x"00052e11",
			2937 => x"01000b04",
			2938 => x"00172e11",
			2939 => x"fffd2e11",
			2940 => x"09001d04",
			2941 => x"ff942e11",
			2942 => x"00032e11",
			2943 => x"0600ab04",
			2944 => x"ffd32e11",
			2945 => x"0c001904",
			2946 => x"00442e11",
			2947 => x"fff62e11",
			2948 => x"0600770c",
			2949 => x"09001808",
			2950 => x"06004904",
			2951 => x"fe852e7d",
			2952 => x"01942e7d",
			2953 => x"fe5c2e7d",
			2954 => x"0200f714",
			2955 => x"05002e10",
			2956 => x"08001d0c",
			2957 => x"08001b08",
			2958 => x"0000cc04",
			2959 => x"02092e7d",
			2960 => x"01912e7d",
			2961 => x"027e2e7d",
			2962 => x"00982e7d",
			2963 => x"fe702e7d",
			2964 => x"0e009104",
			2965 => x"fe602e7d",
			2966 => x"00013210",
			2967 => x"05002e08",
			2968 => x"0e009e04",
			2969 => x"feb92e7d",
			2970 => x"015b2e7d",
			2971 => x"0c002004",
			2972 => x"03de2e7d",
			2973 => x"fe902e7d",
			2974 => x"fe672e7d",
			2975 => x"09001f30",
			2976 => x"0700290c",
			2977 => x"09001808",
			2978 => x"07002504",
			2979 => x"fe642f01",
			2980 => x"027e2f01",
			2981 => x"fe532f01",
			2982 => x"00011e18",
			2983 => x"05002910",
			2984 => x"0200f70c",
			2985 => x"05002508",
			2986 => x"0a002504",
			2987 => x"04202f01",
			2988 => x"032a2f01",
			2989 => x"045f2f01",
			2990 => x"025c2f01",
			2991 => x"07003104",
			2992 => x"fe492f01",
			2993 => x"03842f01",
			2994 => x"0e00a408",
			2995 => x"07003204",
			2996 => x"fe5b2f01",
			2997 => x"003b2f01",
			2998 => x"03902f01",
			2999 => x"01000608",
			3000 => x"07002d04",
			3001 => x"fe622f01",
			3002 => x"02802f01",
			3003 => x"09002108",
			3004 => x"07003404",
			3005 => x"fe5d2f01",
			3006 => x"02302f01",
			3007 => x"fe5a2f01",
			3008 => x"08001c20",
			3009 => x"07002b0c",
			3010 => x"0000a608",
			3011 => x"0e005604",
			3012 => x"ffe52f95",
			3013 => x"00272f95",
			3014 => x"ffce2f95",
			3015 => x"00013210",
			3016 => x"0a003408",
			3017 => x"05002704",
			3018 => x"00742f95",
			3019 => x"00012f95",
			3020 => x"0a004304",
			3021 => x"fff92f95",
			3022 => x"00072f95",
			3023 => x"ffe72f95",
			3024 => x"0e009e20",
			3025 => x"0b001308",
			3026 => x"05002404",
			3027 => x"fff72f95",
			3028 => x"00112f95",
			3029 => x"0200eb0c",
			3030 => x"07003004",
			3031 => x"ffcf2f95",
			3032 => x"05002a04",
			3033 => x"003e2f95",
			3034 => x"fff72f95",
			3035 => x"03003404",
			3036 => x"ff812f95",
			3037 => x"05003b04",
			3038 => x"00172f95",
			3039 => x"fff52f95",
			3040 => x"0a003104",
			3041 => x"00482f95",
			3042 => x"0d001804",
			3043 => x"ffac2f95",
			3044 => x"00292f95",
			3045 => x"0600bd30",
			3046 => x"0200f720",
			3047 => x"0e007b18",
			3048 => x"01000814",
			3049 => x"0000b70c",
			3050 => x"00008904",
			3051 => x"fff33009",
			3052 => x"0b001504",
			3053 => x"00333009",
			3054 => x"ffff3009",
			3055 => x"01000504",
			3056 => x"ffe53009",
			3057 => x"00083009",
			3058 => x"ffc23009",
			3059 => x"07003304",
			3060 => x"003f3009",
			3061 => x"00003009",
			3062 => x"0c001704",
			3063 => x"ff993009",
			3064 => x"0e009104",
			3065 => x"ffe63009",
			3066 => x"0b001904",
			3067 => x"00313009",
			3068 => x"fffb3009",
			3069 => x"0b001304",
			3070 => x"ffed3009",
			3071 => x"01001004",
			3072 => x"00603009",
			3073 => x"ffe33009",
			3074 => x"08001c28",
			3075 => x"0d00141c",
			3076 => x"07002e10",
			3077 => x"0000b708",
			3078 => x"06006b04",
			3079 => x"ffbf30ad",
			3080 => x"008230ad",
			3081 => x"0b001504",
			3082 => x"ff8a30ad",
			3083 => x"000530ad",
			3084 => x"00013308",
			3085 => x"0d001204",
			3086 => x"002930ad",
			3087 => x"00c730ad",
			3088 => x"ffdb30ad",
			3089 => x"00010308",
			3090 => x"0f008d04",
			3091 => x"ffe230ad",
			3092 => x"002330ad",
			3093 => x"ff9a30ad",
			3094 => x"0a002f14",
			3095 => x"0e009410",
			3096 => x"0000f30c",
			3097 => x"0000bc04",
			3098 => x"ffa130ad",
			3099 => x"07002f04",
			3100 => x"ffed30ad",
			3101 => x"006e30ad",
			3102 => x"ff6230ad",
			3103 => x"009530ad",
			3104 => x"0d001810",
			3105 => x"03003408",
			3106 => x"00010704",
			3107 => x"000f30ad",
			3108 => x"ff2730ad",
			3109 => x"05004a04",
			3110 => x"002230ad",
			3111 => x"ffee30ad",
			3112 => x"08001f04",
			3113 => x"004f30ad",
			3114 => x"ffa830ad",
			3115 => x"05002628",
			3116 => x"0201121c",
			3117 => x"0e008314",
			3118 => x"01000b10",
			3119 => x"06006b04",
			3120 => x"ffae3131",
			3121 => x"0000b704",
			3122 => x"008b3131",
			3123 => x"0000d904",
			3124 => x"00053131",
			3125 => x"ffdf3131",
			3126 => x"ff7d3131",
			3127 => x"0c001504",
			3128 => x"010c3131",
			3129 => x"001f3131",
			3130 => x"0b001304",
			3131 => x"ff613131",
			3132 => x"09001b04",
			3133 => x"00733131",
			3134 => x"ffa03131",
			3135 => x"07003304",
			3136 => x"ff303131",
			3137 => x"08001d08",
			3138 => x"03003d04",
			3139 => x"00ac3131",
			3140 => x"ffef3131",
			3141 => x"00010e0c",
			3142 => x"01001108",
			3143 => x"03004904",
			3144 => x"00513131",
			3145 => x"fff73131",
			3146 => x"ffe83131",
			3147 => x"ff3e3131",
			3148 => x"0600bd38",
			3149 => x"00010320",
			3150 => x"0e007714",
			3151 => x"01000810",
			3152 => x"0f007404",
			3153 => x"ff4d31b5",
			3154 => x"0000b704",
			3155 => x"011431b5",
			3156 => x"07002b04",
			3157 => x"ff5931b5",
			3158 => x"fffd31b5",
			3159 => x"fee331b5",
			3160 => x"0b001404",
			3161 => x"fff631b5",
			3162 => x"0e007d04",
			3163 => x"000331b5",
			3164 => x"013231b5",
			3165 => x"03003810",
			3166 => x"0e009e0c",
			3167 => x"01000608",
			3168 => x"04002204",
			3169 => x"ff7631b5",
			3170 => x"004431b5",
			3171 => x"feaa31b5",
			3172 => x"000431b5",
			3173 => x"03003a04",
			3174 => x"009d31b5",
			3175 => x"ffaf31b5",
			3176 => x"0b001304",
			3177 => x"ffe331b5",
			3178 => x"01001004",
			3179 => x"011431b5",
			3180 => x"ff4731b5",
			3181 => x"04001928",
			3182 => x"0700331c",
			3183 => x"0700290c",
			3184 => x"02009008",
			3185 => x"00008904",
			3186 => x"ffe43259",
			3187 => x"00353259",
			3188 => x"ffc73259",
			3189 => x"00011d08",
			3190 => x"09001f04",
			3191 => x"00a53259",
			3192 => x"fffb3259",
			3193 => x"00013104",
			3194 => x"ffc13259",
			3195 => x"00323259",
			3196 => x"07003508",
			3197 => x"08001f04",
			3198 => x"ff993259",
			3199 => x"00073259",
			3200 => x"004b3259",
			3201 => x"04002320",
			3202 => x"00010114",
			3203 => x"0e007d10",
			3204 => x"0b00180c",
			3205 => x"03002108",
			3206 => x"03001e04",
			3207 => x"ffff3259",
			3208 => x"00013259",
			3209 => x"ffbf3259",
			3210 => x"00023259",
			3211 => x"00543259",
			3212 => x"07003904",
			3213 => x"ff713259",
			3214 => x"07003b04",
			3215 => x"00033259",
			3216 => x"fffc3259",
			3217 => x"0e009104",
			3218 => x"ffbf3259",
			3219 => x"00012704",
			3220 => x"00513259",
			3221 => x"fff13259",
			3222 => x"0e009330",
			3223 => x"00010a2c",
			3224 => x"0e006f18",
			3225 => x"09001808",
			3226 => x"00008904",
			3227 => x"ff6a32ed",
			3228 => x"00a632ed",
			3229 => x"0d001108",
			3230 => x"08001804",
			3231 => x"001a32ed",
			3232 => x"fff232ed",
			3233 => x"08001604",
			3234 => x"fffc32ed",
			3235 => x"feb432ed",
			3236 => x"08001d08",
			3237 => x"03003304",
			3238 => x"013e32ed",
			3239 => x"ffb832ed",
			3240 => x"0000f008",
			3241 => x"0200d904",
			3242 => x"ffd532ed",
			3243 => x"00e132ed",
			3244 => x"fec432ed",
			3245 => x"fea332ed",
			3246 => x"08001f10",
			3247 => x"03002a08",
			3248 => x"0b001304",
			3249 => x"007932ed",
			3250 => x"015e32ed",
			3251 => x"0e00a004",
			3252 => x"009d32ed",
			3253 => x"ff7632ed",
			3254 => x"0f00c708",
			3255 => x"08002a04",
			3256 => x"00d532ed",
			3257 => x"ffeb32ed",
			3258 => x"fed932ed",
			3259 => x"0e009334",
			3260 => x"0000f81c",
			3261 => x"0e007918",
			3262 => x"01000810",
			3263 => x"0f007404",
			3264 => x"ff6e3389",
			3265 => x"0000b704",
			3266 => x"00f43389",
			3267 => x"0b001804",
			3268 => x"ff9c3389",
			3269 => x"00213389",
			3270 => x"08001804",
			3271 => x"fffb3389",
			3272 => x"fefc3389",
			3273 => x"00f33389",
			3274 => x"01000608",
			3275 => x"0b001504",
			3276 => x"ffb13389",
			3277 => x"003e3389",
			3278 => x"0800190c",
			3279 => x"08001804",
			3280 => x"ffbe3389",
			3281 => x"0f00c204",
			3282 => x"002e3389",
			3283 => x"fff53389",
			3284 => x"febf3389",
			3285 => x"03002a08",
			3286 => x"00013404",
			3287 => x"00fc3389",
			3288 => x"ff943389",
			3289 => x"03002f08",
			3290 => x"08001c04",
			3291 => x"002a3389",
			3292 => x"fedb3389",
			3293 => x"0e00a008",
			3294 => x"02011f04",
			3295 => x"013a3389",
			3296 => x"ffda3389",
			3297 => x"ff573389",
			3298 => x"0600770c",
			3299 => x"09001708",
			3300 => x"0d001004",
			3301 => x"fe983415",
			3302 => x"012a3415",
			3303 => x"fe5f3415",
			3304 => x"00011628",
			3305 => x"08001c14",
			3306 => x"07002904",
			3307 => x"fe9c3415",
			3308 => x"0a00340c",
			3309 => x"0e008508",
			3310 => x"0000cc04",
			3311 => x"01d53415",
			3312 => x"00cd3415",
			3313 => x"028a3415",
			3314 => x"ffc83415",
			3315 => x"0e008008",
			3316 => x"01000a04",
			3317 => x"ffbd3415",
			3318 => x"fe3a3415",
			3319 => x"0200ec04",
			3320 => x"01f83415",
			3321 => x"03002f04",
			3322 => x"ff143415",
			3323 => x"02223415",
			3324 => x"0600c90c",
			3325 => x"01000a08",
			3326 => x"0e009104",
			3327 => x"fe713415",
			3328 => x"013a3415",
			3329 => x"fe563415",
			3330 => x"03002d04",
			3331 => x"01b43415",
			3332 => x"fe7b3415",
			3333 => x"0600770c",
			3334 => x"09001808",
			3335 => x"03001704",
			3336 => x"fee13481",
			3337 => x"013f3481",
			3338 => x"fe5e3481",
			3339 => x"00013228",
			3340 => x"0e008510",
			3341 => x"01000b0c",
			3342 => x"0200e408",
			3343 => x"05002a04",
			3344 => x"018a3481",
			3345 => x"fefb3481",
			3346 => x"fe7e3481",
			3347 => x"fe513481",
			3348 => x"0d001914",
			3349 => x"0d00150c",
			3350 => x"08001c08",
			3351 => x"08001904",
			3352 => x"00933481",
			3353 => x"017e3481",
			3354 => x"fff43481",
			3355 => x"03002e04",
			3356 => x"01d33481",
			3357 => x"01103481",
			3358 => x"fea93481",
			3359 => x"fe783481",
			3360 => x"09002034",
			3361 => x"0e00630c",
			3362 => x"0b001208",
			3363 => x"07001b04",
			3364 => x"fe8a34fd",
			3365 => x"00d534fd",
			3366 => x"fe5e34fd",
			3367 => x"00011e20",
			3368 => x"0e008010",
			3369 => x"01000b0c",
			3370 => x"0200d808",
			3371 => x"05002104",
			3372 => x"023d34fd",
			3373 => x"018734fd",
			3374 => x"fe6f34fd",
			3375 => x"fe0a34fd",
			3376 => x"03002a0c",
			3377 => x"08001d08",
			3378 => x"0000e304",
			3379 => x"020434fd",
			3380 => x"030b34fd",
			3381 => x"01b434fd",
			3382 => x"016534fd",
			3383 => x"0600c904",
			3384 => x"fe4f34fd",
			3385 => x"01c934fd",
			3386 => x"0c001a08",
			3387 => x"05002a04",
			3388 => x"00ef34fd",
			3389 => x"fe6f34fd",
			3390 => x"fe6234fd",
			3391 => x"0e009334",
			3392 => x"00010a30",
			3393 => x"0e006f18",
			3394 => x"09001808",
			3395 => x"00008904",
			3396 => x"ff713599",
			3397 => x"00a13599",
			3398 => x"0d001108",
			3399 => x"08001804",
			3400 => x"001b3599",
			3401 => x"fff33599",
			3402 => x"01000204",
			3403 => x"00003599",
			3404 => x"febe3599",
			3405 => x"08001d0c",
			3406 => x"03003308",
			3407 => x"07002d04",
			3408 => x"00653599",
			3409 => x"014d3599",
			3410 => x"ffbc3599",
			3411 => x"0000f008",
			3412 => x"0200d904",
			3413 => x"ffdf3599",
			3414 => x"00d43599",
			3415 => x"fed33599",
			3416 => x"feab3599",
			3417 => x"08001f10",
			3418 => x"04001708",
			3419 => x"05002304",
			3420 => x"01083599",
			3421 => x"ffad3599",
			3422 => x"01000c04",
			3423 => x"00173599",
			3424 => x"01443599",
			3425 => x"0f00c708",
			3426 => x"08002a04",
			3427 => x"00c93599",
			3428 => x"ffed3599",
			3429 => x"fee63599",
			3430 => x"07002e1c",
			3431 => x"05001f10",
			3432 => x"0a001c04",
			3433 => x"ffd2364d",
			3434 => x"0000b708",
			3435 => x"00008904",
			3436 => x"fffc364d",
			3437 => x"0068364d",
			3438 => x"ffd7364d",
			3439 => x"03001d04",
			3440 => x"0001364d",
			3441 => x"04001504",
			3442 => x"fffe364d",
			3443 => x"ff6c364d",
			3444 => x"0a00311c",
			3445 => x"05002910",
			3446 => x"0d00180c",
			3447 => x"0d001408",
			3448 => x"0600b004",
			3449 => x"ffcf364d",
			3450 => x"0050364d",
			3451 => x"00e4364d",
			3452 => x"ffcc364d",
			3453 => x"0f00c608",
			3454 => x"0600a104",
			3455 => x"ffef364d",
			3456 => x"002b364d",
			3457 => x"ffae364d",
			3458 => x"01000a08",
			3459 => x"05004104",
			3460 => x"0071364d",
			3461 => x"ffed364d",
			3462 => x"0e00a510",
			3463 => x"04002308",
			3464 => x"0f00b804",
			3465 => x"0005364d",
			3466 => x"ff44364d",
			3467 => x"0f00d804",
			3468 => x"ffc7364d",
			3469 => x"0038364d",
			3470 => x"0e00ac08",
			3471 => x"03003104",
			3472 => x"004b364d",
			3473 => x"fff9364d",
			3474 => x"ffdf364d",
			3475 => x"0e008628",
			3476 => x"01000b24",
			3477 => x"04001f1c",
			3478 => x"07002910",
			3479 => x"05001a0c",
			3480 => x"07002504",
			3481 => x"ffc536f1",
			3482 => x"05001304",
			3483 => x"fffb36f1",
			3484 => x"008d36f1",
			3485 => x"ff5c36f1",
			3486 => x"00010c08",
			3487 => x"06007704",
			3488 => x"fff436f1",
			3489 => x"00ce36f1",
			3490 => x"ffbb36f1",
			3491 => x"05002b04",
			3492 => x"000136f1",
			3493 => x"ff7336f1",
			3494 => x"ff1936f1",
			3495 => x"0a003118",
			3496 => x"05002910",
			3497 => x"0d00140c",
			3498 => x"0c001408",
			3499 => x"02012e04",
			3500 => x"00b336f1",
			3501 => x"ffc836f1",
			3502 => x"ff8736f1",
			3503 => x"012036f1",
			3504 => x"0600ae04",
			3505 => x"002c36f1",
			3506 => x"ff8036f1",
			3507 => x"05002e08",
			3508 => x"07003404",
			3509 => x"002436f1",
			3510 => x"ff5536f1",
			3511 => x"09002008",
			3512 => x"00013c04",
			3513 => x"00d536f1",
			3514 => x"fff136f1",
			3515 => x"ff9436f1",
			3516 => x"0e008b30",
			3517 => x"05001a08",
			3518 => x"00008904",
			3519 => x"ffe33795",
			3520 => x"00413795",
			3521 => x"07003120",
			3522 => x"0e008618",
			3523 => x"05001f10",
			3524 => x"05001c08",
			3525 => x"04001304",
			3526 => x"00003795",
			3527 => x"ffe13795",
			3528 => x"04001304",
			3529 => x"fffc3795",
			3530 => x"001c3795",
			3531 => x"04001604",
			3532 => x"000a3795",
			3533 => x"ff733795",
			3534 => x"04002004",
			3535 => x"fff13795",
			3536 => x"000f3795",
			3537 => x"04001e04",
			3538 => x"00283795",
			3539 => x"ffd33795",
			3540 => x"00011e0c",
			3541 => x"05002704",
			3542 => x"00c63795",
			3543 => x"05002c04",
			3544 => x"fff13795",
			3545 => x"00533795",
			3546 => x"0600ca10",
			3547 => x"03003108",
			3548 => x"03002404",
			3549 => x"00003795",
			3550 => x"ff5f3795",
			3551 => x"0a003704",
			3552 => x"002c3795",
			3553 => x"fff83795",
			3554 => x"03002d04",
			3555 => x"006e3795",
			3556 => x"ffc33795",
			3557 => x"0600770c",
			3558 => x"09001708",
			3559 => x"0b001104",
			3560 => x"ff2b3809",
			3561 => x"00f23809",
			3562 => x"fe723809",
			3563 => x"0001322c",
			3564 => x"0500230c",
			3565 => x"09001a08",
			3566 => x"0a002104",
			3567 => x"00a73809",
			3568 => x"018f3809",
			3569 => x"006c3809",
			3570 => x"0700300c",
			3571 => x"00010108",
			3572 => x"07002c04",
			3573 => x"feda3809",
			3574 => x"009b3809",
			3575 => x"fe803809",
			3576 => x"01000804",
			3577 => x"01773809",
			3578 => x"0200ec08",
			3579 => x"0e007904",
			3580 => x"ff893809",
			3581 => x"017d3809",
			3582 => x"0600b004",
			3583 => x"fea23809",
			3584 => x"00323809",
			3585 => x"fe963809",
			3586 => x"08001c24",
			3587 => x"06006b04",
			3588 => x"ffc938a5",
			3589 => x"0001321c",
			3590 => x"04001908",
			3591 => x"08001604",
			3592 => x"fff938a5",
			3593 => x"008c38a5",
			3594 => x"03002a08",
			3595 => x"07002b04",
			3596 => x"ffe738a5",
			3597 => x"004738a5",
			3598 => x"09001e04",
			3599 => x"ffbe38a5",
			3600 => x"08001904",
			3601 => x"fff938a5",
			3602 => x"001138a5",
			3603 => x"ffce38a5",
			3604 => x"0f00d420",
			3605 => x"0200eb14",
			3606 => x"0700300c",
			3607 => x"04001408",
			3608 => x"04001304",
			3609 => x"fffa38a5",
			3610 => x"000638a5",
			3611 => x"ffab38a5",
			3612 => x"09002104",
			3613 => x"005f38a5",
			3614 => x"fff338a5",
			3615 => x"03003404",
			3616 => x"ff5a38a5",
			3617 => x"04002a04",
			3618 => x"002138a5",
			3619 => x"fff038a5",
			3620 => x"04001804",
			3621 => x"ffb638a5",
			3622 => x"01001004",
			3623 => x"008138a5",
			3624 => x"ffe638a5",
			3625 => x"0f007a0c",
			3626 => x"0b001208",
			3627 => x"0b001004",
			3628 => x"feb43931",
			3629 => x"00ce3931",
			3630 => x"fe653931",
			3631 => x"00011e28",
			3632 => x"05004024",
			3633 => x"0400170c",
			3634 => x"0c001404",
			3635 => x"02453931",
			3636 => x"0000e904",
			3637 => x"01c03931",
			3638 => x"01123931",
			3639 => x"0700300c",
			3640 => x"0d001408",
			3641 => x"00010104",
			3642 => x"01553931",
			3643 => x"fe803931",
			3644 => x"fe4b3931",
			3645 => x"0d001908",
			3646 => x"01000a04",
			3647 => x"02233931",
			3648 => x"01033931",
			3649 => x"fe953931",
			3650 => x"fe753931",
			3651 => x"0600c90c",
			3652 => x"0d001108",
			3653 => x"05002e04",
			3654 => x"fe9b3931",
			3655 => x"016a3931",
			3656 => x"fe5e3931",
			3657 => x"03002a04",
			3658 => x"01963931",
			3659 => x"fe623931",
			3660 => x"0e008534",
			3661 => x"0400191c",
			3662 => x"01000910",
			3663 => x"06006b04",
			3664 => x"ff6d39d5",
			3665 => x"0000b704",
			3666 => x"012c39d5",
			3667 => x"09001904",
			3668 => x"ff9139d5",
			3669 => x"002939d5",
			3670 => x"07002c04",
			3671 => x"ff1a39d5",
			3672 => x"0a002004",
			3673 => x"ffd939d5",
			3674 => x"001d39d5",
			3675 => x"07003410",
			3676 => x"0300210c",
			3677 => x"03001f08",
			3678 => x"05002204",
			3679 => x"ffcb39d5",
			3680 => x"fffe39d5",
			3681 => x"002239d5",
			3682 => x"feba39d5",
			3683 => x"05002904",
			3684 => x"006439d5",
			3685 => x"ff9139d5",
			3686 => x"0001321c",
			3687 => x"05002304",
			3688 => x"011439d5",
			3689 => x"05002504",
			3690 => x"ff4439d5",
			3691 => x"0200f704",
			3692 => x"014c39d5",
			3693 => x"03002f08",
			3694 => x"0e00a104",
			3695 => x"ff2339d5",
			3696 => x"008139d5",
			3697 => x"0600b004",
			3698 => x"ff8539d5",
			3699 => x"012f39d5",
			3700 => x"fefe39d5",
			3701 => x"0f007404",
			3702 => x"fe6f3a41",
			3703 => x"05003028",
			3704 => x"00013224",
			3705 => x"01000810",
			3706 => x"02011208",
			3707 => x"0b001304",
			3708 => x"00eb3a41",
			3709 => x"01a43a41",
			3710 => x"05002504",
			3711 => x"009a3a41",
			3712 => x"fee23a41",
			3713 => x"0e007d08",
			3714 => x"01000b04",
			3715 => x"ff8f3a41",
			3716 => x"fe423a41",
			3717 => x"0000f804",
			3718 => x"01ae3a41",
			3719 => x"0600b004",
			3720 => x"fe763a41",
			3721 => x"00bc3a41",
			3722 => x"fe863a41",
			3723 => x"0e009604",
			3724 => x"fe703a41",
			3725 => x"0f00c704",
			3726 => x"01853a41",
			3727 => x"fe9c3a41",
			3728 => x"0c001208",
			3729 => x"08001b04",
			3730 => x"ff4e3ad5",
			3731 => x"018b3ad5",
			3732 => x"05002010",
			3733 => x"06007008",
			3734 => x"0b001304",
			3735 => x"00833ad5",
			3736 => x"fef73ad5",
			3737 => x"0b001304",
			3738 => x"00693ad5",
			3739 => x"014f3ad5",
			3740 => x"07002e10",
			3741 => x"04001604",
			3742 => x"00153ad5",
			3743 => x"08001504",
			3744 => x"00033ad5",
			3745 => x"0a002304",
			3746 => x"ffe63ad5",
			3747 => x"fe9e3ad5",
			3748 => x"00011e14",
			3749 => x"0a00340c",
			3750 => x"05002404",
			3751 => x"ff313ad5",
			3752 => x"0200f704",
			3753 => x"014c3ad5",
			3754 => x"00273ad5",
			3755 => x"01000804",
			3756 => x"00283ad5",
			3757 => x"feb43ad5",
			3758 => x"01000a08",
			3759 => x"0d001304",
			3760 => x"00f63ad5",
			3761 => x"ff7b3ad5",
			3762 => x"03002604",
			3763 => x"00803ad5",
			3764 => x"fe7e3ad5",
			3765 => x"0c001208",
			3766 => x"08001b04",
			3767 => x"ff583b71",
			3768 => x"01743b71",
			3769 => x"05002010",
			3770 => x"06007008",
			3771 => x"0b001304",
			3772 => x"00823b71",
			3773 => x"ff053b71",
			3774 => x"0b001304",
			3775 => x"005e3b71",
			3776 => x"01463b71",
			3777 => x"07002e10",
			3778 => x"04001604",
			3779 => x"00183b71",
			3780 => x"08001504",
			3781 => x"00033b71",
			3782 => x"0a002304",
			3783 => x"ffe73b71",
			3784 => x"fea63b71",
			3785 => x"00011e18",
			3786 => x"0a003410",
			3787 => x"0d001508",
			3788 => x"08001b04",
			3789 => x"011f3b71",
			3790 => x"ff903b71",
			3791 => x"0e008004",
			3792 => x"ff543b71",
			3793 => x"01263b71",
			3794 => x"01000804",
			3795 => x"00273b71",
			3796 => x"fec13b71",
			3797 => x"01000a08",
			3798 => x"00013b04",
			3799 => x"00ed3b71",
			3800 => x"ff823b71",
			3801 => x"03002604",
			3802 => x"00813b71",
			3803 => x"fe853b71",
			3804 => x"0f007404",
			3805 => x"fe6d3bd7",
			3806 => x"0001322c",
			3807 => x"05004028",
			3808 => x"01000a14",
			3809 => x"0200f708",
			3810 => x"05002704",
			3811 => x"01b63bd7",
			3812 => x"01233bd7",
			3813 => x"0a002d04",
			3814 => x"fe6b3bd7",
			3815 => x"0e008304",
			3816 => x"feb63bd7",
			3817 => x"01ca3bd7",
			3818 => x"0e008508",
			3819 => x"07003304",
			3820 => x"fe4d3bd7",
			3821 => x"00d83bd7",
			3822 => x"05002304",
			3823 => x"01ee3bd7",
			3824 => x"00010f04",
			3825 => x"012a3bd7",
			3826 => x"ffc03bd7",
			3827 => x"fe7b3bd7",
			3828 => x"fe713bd7",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1331, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2571, initial_addr_3'length));
	end generate gen_rom_1;

	gen_rom_2: if SELECT_ROM = 2 generate
		bank <= (
			0 => x"09001d2c",
			1 => x"00012110",
			2 => x"0a00370c",
			3 => x"0a003104",
			4 => x"ce1d007d",
			5 => x"01000804",
			6 => x"d351007d",
			7 => x"ce2b007d",
			8 => x"da40007d",
			9 => x"0500280c",
			10 => x"05002504",
			11 => x"ce23007d",
			12 => x"08001b04",
			13 => x"dc41007d",
			14 => x"ce2f007d",
			15 => x"01000a08",
			16 => x"05002c04",
			17 => x"e5bb007d",
			18 => x"ed92007d",
			19 => x"0f00cb04",
			20 => x"de43007d",
			21 => x"ce36007d",
			22 => x"0c001a10",
			23 => x"0a003d04",
			24 => x"ce1d007d",
			25 => x"01000908",
			26 => x"06007004",
			27 => x"ce23007d",
			28 => x"d038007d",
			29 => x"d562007d",
			30 => x"ce1c007d",
			31 => x"09001c28",
			32 => x"0500270c",
			33 => x"08001504",
			34 => x"001f0101",
			35 => x"03002a04",
			36 => x"ff8e0101",
			37 => x"00030101",
			38 => x"0c001408",
			39 => x"0600a504",
			40 => x"ff9c0101",
			41 => x"00440101",
			42 => x"01000b10",
			43 => x"00010a04",
			44 => x"ffdc0101",
			45 => x"0600a504",
			46 => x"00a10101",
			47 => x"0f00c904",
			48 => x"ffc20101",
			49 => x"00730101",
			50 => x"ffc90101",
			51 => x"08001808",
			52 => x"0f006f04",
			53 => x"ffe40101",
			54 => x"00320101",
			55 => x"0e004d08",
			56 => x"00009f04",
			57 => x"ffef0101",
			58 => x"00210101",
			59 => x"0a004504",
			60 => x"ff920101",
			61 => x"0a004704",
			62 => x"00160101",
			63 => x"ffeb0101",
			64 => x"09001d28",
			65 => x"00010708",
			66 => x"03003104",
			67 => x"fe560175",
			68 => x"ff5b0175",
			69 => x"05002708",
			70 => x"04001a04",
			71 => x"fe5b0175",
			72 => x"00dc0175",
			73 => x"01000b10",
			74 => x"08001c0c",
			75 => x"0f00b304",
			76 => x"0a610175",
			77 => x"02013004",
			78 => x"04f70175",
			79 => x"075b0175",
			80 => x"01da0175",
			81 => x"07003104",
			82 => x"fe570175",
			83 => x"00b80175",
			84 => x"0c001a10",
			85 => x"0a003d04",
			86 => x"fe560175",
			87 => x"05004e08",
			88 => x"06006404",
			89 => x"00640175",
			90 => x"05f90175",
			91 => x"fe5a0175",
			92 => x"fe550175",
			93 => x"09001d20",
			94 => x"0000e704",
			95 => x"fe6201d9",
			96 => x"0e009018",
			97 => x"05002504",
			98 => x"fe6c01d9",
			99 => x"0a00340c",
			100 => x"08001c08",
			101 => x"02012f04",
			102 => x"00e901d9",
			103 => x"027c01d9",
			104 => x"fdf401d9",
			105 => x"0d001204",
			106 => x"021c01d9",
			107 => x"02f301d9",
			108 => x"fe5101d9",
			109 => x"0c001a10",
			110 => x"0a003d04",
			111 => x"fe6301d9",
			112 => x"01000908",
			113 => x"04004304",
			114 => x"fe5c01d9",
			115 => x"018201d9",
			116 => x"024201d9",
			117 => x"fe6101d9",
			118 => x"09001d30",
			119 => x"0001070c",
			120 => x"0000e704",
			121 => x"fe57025d",
			122 => x"0000f304",
			123 => x"00ad025d",
			124 => x"fe6e025d",
			125 => x"04001d10",
			126 => x"03002708",
			127 => x"02013704",
			128 => x"fe42025d",
			129 => x"ffde025d",
			130 => x"0e009904",
			131 => x"03ef025d",
			132 => x"fe70025d",
			133 => x"0e009210",
			134 => x"02011204",
			135 => x"07a1025d",
			136 => x"08001c08",
			137 => x"04002004",
			138 => x"03ad025d",
			139 => x"04dc025d",
			140 => x"0233025d",
			141 => x"fe46025d",
			142 => x"0b001810",
			143 => x"0a003d04",
			144 => x"fe59025d",
			145 => x"04003604",
			146 => x"0309025d",
			147 => x"04004304",
			148 => x"fe5c025d",
			149 => x"00a2025d",
			150 => x"fe57025d",
			151 => x"0c001a28",
			152 => x"0600670c",
			153 => x"08001c04",
			154 => x"fe6402b1",
			155 => x"0d001304",
			156 => x"01b102b1",
			157 => x"fe7d02b1",
			158 => x"0e009018",
			159 => x"05002504",
			160 => x"fe7102b1",
			161 => x"0d001610",
			162 => x"0a003408",
			163 => x"09001c04",
			164 => x"00ef02b1",
			165 => x"fef302b1",
			166 => x"05004e04",
			167 => x"01cf02b1",
			168 => x"fe9e02b1",
			169 => x"fe6d02b1",
			170 => x"fe5302b1",
			171 => x"fe6702b1",
			172 => x"07002b1c",
			173 => x"02011614",
			174 => x"0a003d08",
			175 => x"08001504",
			176 => x"00080345",
			177 => x"ffa10345",
			178 => x"00009f04",
			179 => x"fff20345",
			180 => x"05004e04",
			181 => x"004f0345",
			182 => x"fff60345",
			183 => x"01000804",
			184 => x"00840345",
			185 => x"fff60345",
			186 => x"02012f28",
			187 => x"0600a114",
			188 => x"0f00a70c",
			189 => x"01000c04",
			190 => x"ffba0345",
			191 => x"01000d04",
			192 => x"00140345",
			193 => x"fff90345",
			194 => x"01000b04",
			195 => x"003f0345",
			196 => x"fff30345",
			197 => x"07002e04",
			198 => x"ff6f0345",
			199 => x"0700320c",
			200 => x"08001f08",
			201 => x"04001d04",
			202 => x"fffa0345",
			203 => x"00390345",
			204 => x"fff70345",
			205 => x"ffec0345",
			206 => x"07002f04",
			207 => x"006c0345",
			208 => x"ffce0345",
			209 => x"0e008a3c",
			210 => x"00012f28",
			211 => x"0900190c",
			212 => x"08001804",
			213 => x"ff0603e1",
			214 => x"08001b04",
			215 => x"000103e1",
			216 => x"ffe503e1",
			217 => x"0c001508",
			218 => x"0a002d04",
			219 => x"ffec03e1",
			220 => x"00cb03e1",
			221 => x"00012710",
			222 => x"0a004308",
			223 => x"0e004d04",
			224 => x"003703e1",
			225 => x"ff1603e1",
			226 => x"05004e04",
			227 => x"009c03e1",
			228 => x"ffc703e1",
			229 => x"007b03e1",
			230 => x"0d00130c",
			231 => x"08001908",
			232 => x"0f00c804",
			233 => x"00fb03e1",
			234 => x"005003e1",
			235 => x"000c03e1",
			236 => x"0f00c504",
			237 => x"005a03e1",
			238 => x"ff4403e1",
			239 => x"0b001308",
			240 => x"0a002f04",
			241 => x"ffed03e1",
			242 => x"003b03e1",
			243 => x"01000904",
			244 => x"ff1603e1",
			245 => x"01000b04",
			246 => x"002603e1",
			247 => x"ffc503e1",
			248 => x"08001c2c",
			249 => x"02012f24",
			250 => x"02012b20",
			251 => x"00012f18",
			252 => x"0b00150c",
			253 => x"0d000e04",
			254 => x"00370465",
			255 => x"0a003404",
			256 => x"ff590465",
			257 => x"002f0465",
			258 => x"00010a08",
			259 => x"03003b04",
			260 => x"ffa40465",
			261 => x"00250465",
			262 => x"00730465",
			263 => x"04001f04",
			264 => x"00030465",
			265 => x"00990465",
			266 => x"ff890465",
			267 => x"05002704",
			268 => x"ffcb0465",
			269 => x"00a50465",
			270 => x"03003308",
			271 => x"05003e04",
			272 => x"ff750465",
			273 => x"00050465",
			274 => x"0c001a0c",
			275 => x"0a003704",
			276 => x"fff40465",
			277 => x"01000904",
			278 => x"fff90465",
			279 => x"00400465",
			280 => x"ffe10465",
			281 => x"09001d34",
			282 => x"0001070c",
			283 => x"0000e704",
			284 => x"fe5a04f1",
			285 => x"0c001504",
			286 => x"00c304f1",
			287 => x"fe6c04f1",
			288 => x"04001d10",
			289 => x"03002708",
			290 => x"02013704",
			291 => x"fe4504f1",
			292 => x"ffd804f1",
			293 => x"0f00d504",
			294 => x"032a04f1",
			295 => x"fe7304f1",
			296 => x"0e009214",
			297 => x"08001c10",
			298 => x"04002008",
			299 => x"0f00c504",
			300 => x"01e904f1",
			301 => x"03b304f1",
			302 => x"0f00b904",
			303 => x"04da04f1",
			304 => x"03bb04f1",
			305 => x"016904f1",
			306 => x"fe4b04f1",
			307 => x"0b001810",
			308 => x"0a003d04",
			309 => x"fe5c04f1",
			310 => x"01000908",
			311 => x"04004304",
			312 => x"fe5d04f1",
			313 => x"00d404f1",
			314 => x"02b104f1",
			315 => x"fe5904f1",
			316 => x"0d001330",
			317 => x"0e008a28",
			318 => x"00012f20",
			319 => x"0a003410",
			320 => x"0b001204",
			321 => x"001e0585",
			322 => x"0b001608",
			323 => x"04001804",
			324 => x"ffff0585",
			325 => x"ff8a0585",
			326 => x"000b0585",
			327 => x"0900200c",
			328 => x"06005504",
			329 => x"fff90585",
			330 => x"05004e04",
			331 => x"004e0585",
			332 => x"fffc0585",
			333 => x"ffeb0585",
			334 => x"01000804",
			335 => x"00720585",
			336 => x"fffd0585",
			337 => x"0b001304",
			338 => x"00100585",
			339 => x"ffa30585",
			340 => x"08001808",
			341 => x"0f00a504",
			342 => x"fff80585",
			343 => x"00300585",
			344 => x"0a00450c",
			345 => x"0b001408",
			346 => x"0c001404",
			347 => x"ffed0585",
			348 => x"000d0585",
			349 => x"ff910585",
			350 => x"03004004",
			351 => x"00140585",
			352 => x"fff00585",
			353 => x"0e008a40",
			354 => x"0c001410",
			355 => x"0600a50c",
			356 => x"04002008",
			357 => x"08001504",
			358 => x"00130629",
			359 => x"ff5c0629",
			360 => x"00260629",
			361 => x"002a0629",
			362 => x"00010714",
			363 => x"05004c0c",
			364 => x"0e004d08",
			365 => x"00009f04",
			366 => x"ffe30629",
			367 => x"00280629",
			368 => x"ff6f0629",
			369 => x"05004e04",
			370 => x"00620629",
			371 => x"ffd30629",
			372 => x"0100090c",
			373 => x"04002908",
			374 => x"0f00c604",
			375 => x"00c00629",
			376 => x"00110629",
			377 => x"fff40629",
			378 => x"05003108",
			379 => x"00013b04",
			380 => x"ff790629",
			381 => x"00100629",
			382 => x"09001e04",
			383 => x"00640629",
			384 => x"ffe50629",
			385 => x"0b001308",
			386 => x"0f00dd04",
			387 => x"00280629",
			388 => x"fff90629",
			389 => x"01000904",
			390 => x"ff7e0629",
			391 => x"01000b04",
			392 => x"000b0629",
			393 => x"ffe80629",
			394 => x"09001c30",
			395 => x"05002708",
			396 => x"03002a04",
			397 => x"fe6906bd",
			398 => x"00e706bd",
			399 => x"08001c20",
			400 => x"01000508",
			401 => x"0f00bc04",
			402 => x"fe9206bd",
			403 => x"00b506bd",
			404 => x"05002c0c",
			405 => x"0f00ca08",
			406 => x"07002b04",
			407 => x"00e306bd",
			408 => x"ff6306bd",
			409 => x"018806bd",
			410 => x"0a002d04",
			411 => x"008d06bd",
			412 => x"06007304",
			413 => x"ff4a06bd",
			414 => x"01d206bd",
			415 => x"0f00bf04",
			416 => x"ff9006bd",
			417 => x"fe5106bd",
			418 => x"0a003708",
			419 => x"08001804",
			420 => x"fff806bd",
			421 => x"fe5806bd",
			422 => x"09002110",
			423 => x"0e006508",
			424 => x"06005804",
			425 => x"016306bd",
			426 => x"fe6406bd",
			427 => x"08001b04",
			428 => x"ff9f06bd",
			429 => x"01cc06bd",
			430 => x"fe7d06bd",
			431 => x"02010218",
			432 => x"0a003404",
			433 => x"fe5a0761",
			434 => x"04002704",
			435 => x"01df0761",
			436 => x"01000408",
			437 => x"08001904",
			438 => x"fe790761",
			439 => x"024a0761",
			440 => x"08001804",
			441 => x"008e0761",
			442 => x"fe5a0761",
			443 => x"08001c2c",
			444 => x"03002714",
			445 => x"0d00120c",
			446 => x"04001d08",
			447 => x"09001804",
			448 => x"fe1c0761",
			449 => x"00770761",
			450 => x"025c0761",
			451 => x"07002d04",
			452 => x"fdfa0761",
			453 => x"ff9d0761",
			454 => x"0e008a10",
			455 => x"0c001404",
			456 => x"01470761",
			457 => x"06009f04",
			458 => x"02b70761",
			459 => x"0f00c104",
			460 => x"01230761",
			461 => x"021a0761",
			462 => x"02012d04",
			463 => x"febe0761",
			464 => x"01350761",
			465 => x"0a003708",
			466 => x"07002e04",
			467 => x"fdf00761",
			468 => x"fe670761",
			469 => x"0e008804",
			470 => x"01c90761",
			471 => x"fe5e0761",
			472 => x"01000d28",
			473 => x"01000308",
			474 => x"0d001104",
			475 => x"fe3907b5",
			476 => x"ffce07b5",
			477 => x"03002204",
			478 => x"fe8d07b5",
			479 => x"0e009018",
			480 => x"00013a10",
			481 => x"0a003408",
			482 => x"01000904",
			483 => x"005907b5",
			484 => x"fec607b5",
			485 => x"05004e04",
			486 => x"010407b5",
			487 => x"fea507b5",
			488 => x"0d001304",
			489 => x"019107b5",
			490 => x"002907b5",
			491 => x"fe9007b5",
			492 => x"fe7107b5",
			493 => x"0a002d1c",
			494 => x"07002e10",
			495 => x"0e007e08",
			496 => x"0f00ba04",
			497 => x"ff630871",
			498 => x"00900871",
			499 => x"00013f04",
			500 => x"fef40871",
			501 => x"000d0871",
			502 => x"0b001508",
			503 => x"0e009104",
			504 => x"00b60871",
			505 => x"ffcd0871",
			506 => x"ffb60871",
			507 => x"01000b2c",
			508 => x"0600a21c",
			509 => x"07002b14",
			510 => x"0e005d0c",
			511 => x"08001c04",
			512 => x"ff860871",
			513 => x"06005904",
			514 => x"00550871",
			515 => x"ffe50871",
			516 => x"0d001204",
			517 => x"ffe30871",
			518 => x"00cc0871",
			519 => x"0a003204",
			520 => x"00090871",
			521 => x"ff500871",
			522 => x"0e008b08",
			523 => x"05003504",
			524 => x"01220871",
			525 => x"00140871",
			526 => x"0b001404",
			527 => x"00370871",
			528 => x"ff860871",
			529 => x"0000c808",
			530 => x"0200ad04",
			531 => x"fff00871",
			532 => x"004a0871",
			533 => x"07003104",
			534 => x"ff510871",
			535 => x"07003308",
			536 => x"0f00b804",
			537 => x"003a0871",
			538 => x"fff30871",
			539 => x"ffc40871",
			540 => x"0e008a3c",
			541 => x"00012f2c",
			542 => x"05002c14",
			543 => x"0c00170c",
			544 => x"0b001208",
			545 => x"06005404",
			546 => x"ffd00905",
			547 => x"01080905",
			548 => x"fe730905",
			549 => x"09001c04",
			550 => x"012d0905",
			551 => x"ff760905",
			552 => x"04003814",
			553 => x"05004c10",
			554 => x"0e006f08",
			555 => x"07002604",
			556 => x"009a0905",
			557 => x"fe910905",
			558 => x"03002c04",
			559 => x"ff800905",
			560 => x"011b0905",
			561 => x"017f0905",
			562 => x"fec10905",
			563 => x"0d001204",
			564 => x"018b0905",
			565 => x"0a002d04",
			566 => x"fee40905",
			567 => x"01000a04",
			568 => x"01540905",
			569 => x"ff330905",
			570 => x"09001b0c",
			571 => x"00013f08",
			572 => x"0f00c704",
			573 => x"00900905",
			574 => x"fef30905",
			575 => x"00a90905",
			576 => x"fea00905",
			577 => x"0d001338",
			578 => x"04001d10",
			579 => x"0300270c",
			580 => x"03002308",
			581 => x"03002104",
			582 => x"fff309a1",
			583 => x"002109a1",
			584 => x"ff4809a1",
			585 => x"001609a1",
			586 => x"0f00c420",
			587 => x"07002b14",
			588 => x"01000a10",
			589 => x"0c001608",
			590 => x"07002504",
			591 => x"fff609a1",
			592 => x"00ab09a1",
			593 => x"03003504",
			594 => x"ffab09a1",
			595 => x"005d09a1",
			596 => x"ffc309a1",
			597 => x"04002204",
			598 => x"ff7d09a1",
			599 => x"00011404",
			600 => x"ffd709a1",
			601 => x"004809a1",
			602 => x"01000704",
			603 => x"002409a1",
			604 => x"00b609a1",
			605 => x"08001804",
			606 => x"006109a1",
			607 => x"0b001408",
			608 => x"03002c04",
			609 => x"ffdd09a1",
			610 => x"003d09a1",
			611 => x"0a004504",
			612 => x"ff2f09a1",
			613 => x"03004004",
			614 => x"002709a1",
			615 => x"ffe709a1",
			616 => x"0a002d24",
			617 => x"0f00c918",
			618 => x"05002b0c",
			619 => x"03002308",
			620 => x"03002104",
			621 => x"ffab0a5d",
			622 => x"00070a5d",
			623 => x"feb00a5d",
			624 => x"04001f04",
			625 => x"00e60a5d",
			626 => x"03002604",
			627 => x"00520a5d",
			628 => x"ff290a5d",
			629 => x"0e008a04",
			630 => x"00980a5d",
			631 => x"0b001304",
			632 => x"002e0a5d",
			633 => x"ff2d0a5d",
			634 => x"02012328",
			635 => x"05004c20",
			636 => x"0e006f0c",
			637 => x"0e004d08",
			638 => x"08001c04",
			639 => x"ffb60a5d",
			640 => x"00ab0a5d",
			641 => x"fec70a5d",
			642 => x"02012110",
			643 => x"07002c08",
			644 => x"0e007b04",
			645 => x"00460a5d",
			646 => x"00d70a5d",
			647 => x"0d001304",
			648 => x"00030a5d",
			649 => x"ff3f0a5d",
			650 => x"ff3b0a5d",
			651 => x"05004e04",
			652 => x"00ea0a5d",
			653 => x"ff760a5d",
			654 => x"08001c08",
			655 => x"0e008904",
			656 => x"015a0a5d",
			657 => x"ffb50a5d",
			658 => x"0a003b04",
			659 => x"ff2e0a5d",
			660 => x"03003404",
			661 => x"002c0a5d",
			662 => x"fff50a5d",
			663 => x"01000a3c",
			664 => x"01000308",
			665 => x"0d001104",
			666 => x"fe7f0b01",
			667 => x"00400b01",
			668 => x"06009b18",
			669 => x"0d001208",
			670 => x"01000804",
			671 => x"feb00b01",
			672 => x"ffdd0b01",
			673 => x"0400360c",
			674 => x"0a003104",
			675 => x"fecd0b01",
			676 => x"03003504",
			677 => x"00380b01",
			678 => x"01510b01",
			679 => x"fecd0b01",
			680 => x"0b00140c",
			681 => x"05002504",
			682 => x"ff4a0b01",
			683 => x"03002904",
			684 => x"00d30b01",
			685 => x"018a0b01",
			686 => x"0e008004",
			687 => x"00e60b01",
			688 => x"0e008304",
			689 => x"fef40b01",
			690 => x"0e008a04",
			691 => x"01170b01",
			692 => x"ff250b01",
			693 => x"0d001208",
			694 => x"08001904",
			695 => x"00fc0b01",
			696 => x"ff6a0b01",
			697 => x"0b001308",
			698 => x"0600b304",
			699 => x"ff350b01",
			700 => x"007e0b01",
			701 => x"0c001404",
			702 => x"ffd00b01",
			703 => x"fe810b01",
			704 => x"0e008a48",
			705 => x"00011e24",
			706 => x"05004c1c",
			707 => x"0700260c",
			708 => x"00009f04",
			709 => x"ffb90bad",
			710 => x"08001b04",
			711 => x"ffe90bad",
			712 => x"007f0bad",
			713 => x"00010a04",
			714 => x"ff260bad",
			715 => x"0d001404",
			716 => x"ffa30bad",
			717 => x"0f00b004",
			718 => x"00750bad",
			719 => x"ffe40bad",
			720 => x"05004e04",
			721 => x"008c0bad",
			722 => x"ffb50bad",
			723 => x"01000910",
			724 => x"03002608",
			725 => x"02012904",
			726 => x"00480bad",
			727 => x"ffbf0bad",
			728 => x"0a002d04",
			729 => x"00340bad",
			730 => x"01110bad",
			731 => x"03002c08",
			732 => x"00013904",
			733 => x"ff3c0bad",
			734 => x"004b0bad",
			735 => x"05003604",
			736 => x"00850bad",
			737 => x"04002904",
			738 => x"ffc00bad",
			739 => x"000b0bad",
			740 => x"01000904",
			741 => x"ff570bad",
			742 => x"09001a08",
			743 => x"0f00d404",
			744 => x"00480bad",
			745 => x"fff10bad",
			746 => x"ffc10bad",
			747 => x"00012f44",
			748 => x"0a003424",
			749 => x"0b001208",
			750 => x"0c001304",
			751 => x"fffc0c69",
			752 => x"00430c69",
			753 => x"0400190c",
			754 => x"06009c08",
			755 => x"0e007804",
			756 => x"fff70c69",
			757 => x"00400c69",
			758 => x"ffda0c69",
			759 => x"05003008",
			760 => x"0600a804",
			761 => x"ff3a0c69",
			762 => x"000c0c69",
			763 => x"06009104",
			764 => x"ffca0c69",
			765 => x"00380c69",
			766 => x"09001e08",
			767 => x"04003104",
			768 => x"00850c69",
			769 => x"ffe20c69",
			770 => x"0f007c14",
			771 => x"0400380c",
			772 => x"01000904",
			773 => x"ffe50c69",
			774 => x"03003804",
			775 => x"fff60c69",
			776 => x"00820c69",
			777 => x"06007204",
			778 => x"ffb40c69",
			779 => x"00300c69",
			780 => x"ff850c69",
			781 => x"0800190c",
			782 => x"0d001308",
			783 => x"04001d04",
			784 => x"00280c69",
			785 => x"00d00c69",
			786 => x"ffea0c69",
			787 => x"08001c08",
			788 => x"0a002d04",
			789 => x"ffcb0c69",
			790 => x"00550c69",
			791 => x"0a003b04",
			792 => x"ff870c69",
			793 => x"00090c69",
			794 => x"0c001414",
			795 => x"0600a50c",
			796 => x"08001504",
			797 => x"002e0d15",
			798 => x"0d001304",
			799 => x"feb30d15",
			800 => x"003b0d15",
			801 => x"01000804",
			802 => x"01120d15",
			803 => x"ff770d15",
			804 => x"0e008a38",
			805 => x"01000920",
			806 => x"0e007410",
			807 => x"04004308",
			808 => x"0c001504",
			809 => x"00570d15",
			810 => x"feef0d15",
			811 => x"01000604",
			812 => x"00c40d15",
			813 => x"ffe10d15",
			814 => x"03002608",
			815 => x"0d001204",
			816 => x"00880d15",
			817 => x"ff800d15",
			818 => x"00012104",
			819 => x"004c0d15",
			820 => x"01590d15",
			821 => x"05003108",
			822 => x"0f00c604",
			823 => x"fea80d15",
			824 => x"00780d15",
			825 => x"0d00160c",
			826 => x"04003808",
			827 => x"01000d04",
			828 => x"00ee0d15",
			829 => x"ffca0d15",
			830 => x"ff850d15",
			831 => x"ff5e0d15",
			832 => x"0c001608",
			833 => x"0600b604",
			834 => x"00a70d15",
			835 => x"ff700d15",
			836 => x"fef90d15",
			837 => x"01000d28",
			838 => x"05002504",
			839 => x"fe990d69",
			840 => x"08001504",
			841 => x"01390d69",
			842 => x"05004c14",
			843 => x"04003410",
			844 => x"0a003708",
			845 => x"08001c04",
			846 => x"00080d69",
			847 => x"fe6e0d69",
			848 => x"00010c04",
			849 => x"00840d69",
			850 => x"018a0d69",
			851 => x"fe750d69",
			852 => x"05004f08",
			853 => x"0f006d04",
			854 => x"ff770d69",
			855 => x"01b50d69",
			856 => x"fec10d69",
			857 => x"fe820d69",
			858 => x"0d00163c",
			859 => x"0a003724",
			860 => x"08001c20",
			861 => x"02012f14",
			862 => x"0100090c",
			863 => x"02012c08",
			864 => x"0c001404",
			865 => x"ff740de5",
			866 => x"00f70de5",
			867 => x"fec80de5",
			868 => x"05003104",
			869 => x"fe580de5",
			870 => x"015a0de5",
			871 => x"0600b608",
			872 => x"00014204",
			873 => x"00e30de5",
			874 => x"01910de5",
			875 => x"febb0de5",
			876 => x"fe790de5",
			877 => x"01000910",
			878 => x"0e006504",
			879 => x"feb60de5",
			880 => x"01000504",
			881 => x"011a0de5",
			882 => x"00011004",
			883 => x"fec90de5",
			884 => x"00930de5",
			885 => x"04003804",
			886 => x"01b60de5",
			887 => x"fee10de5",
			888 => x"fe950de5",
			889 => x"0d001340",
			890 => x"00012f2c",
			891 => x"0a003418",
			892 => x"0b001204",
			893 => x"00360e99",
			894 => x"0e008310",
			895 => x"04001808",
			896 => x"07002904",
			897 => x"fff00e99",
			898 => x"00110e99",
			899 => x"07002804",
			900 => x"00040e99",
			901 => x"ff5d0e99",
			902 => x"000b0e99",
			903 => x"09002010",
			904 => x"05004e0c",
			905 => x"06005504",
			906 => x"fff80e99",
			907 => x"0d001204",
			908 => x"00040e99",
			909 => x"005b0e99",
			910 => x"fff60e99",
			911 => x"ffea0e99",
			912 => x"04001904",
			913 => x"ffb10e99",
			914 => x"08001b0c",
			915 => x"00013904",
			916 => x"00ac0e99",
			917 => x"00014004",
			918 => x"00070e99",
			919 => x"00380e99",
			920 => x"fffa0e99",
			921 => x"08001808",
			922 => x"04003604",
			923 => x"00620e99",
			924 => x"fff30e99",
			925 => x"0b001408",
			926 => x"03002c04",
			927 => x"ffe70e99",
			928 => x"00210e99",
			929 => x"0a004504",
			930 => x"ff7c0e99",
			931 => x"03004104",
			932 => x"001b0e99",
			933 => x"ffee0e99",
			934 => x"0b001830",
			935 => x"0e00902c",
			936 => x"0a003718",
			937 => x"08001c14",
			938 => x"00013c10",
			939 => x"08001508",
			940 => x"0000c704",
			941 => x"ff7b0efd",
			942 => x"02080efd",
			943 => x"0f00c604",
			944 => x"00330efd",
			945 => x"fe840efd",
			946 => x"018f0efd",
			947 => x"fe5b0efd",
			948 => x"0400360c",
			949 => x"01000908",
			950 => x"00010704",
			951 => x"fec10efd",
			952 => x"01850efd",
			953 => x"01e40efd",
			954 => x"04004304",
			955 => x"fe8b0efd",
			956 => x"01bf0efd",
			957 => x"fe7b0efd",
			958 => x"fe740efd",
			959 => x"08001508",
			960 => x"09001804",
			961 => x"ffe40f81",
			962 => x"00830f81",
			963 => x"05002708",
			964 => x"03002c04",
			965 => x"ff530f81",
			966 => x"00080f81",
			967 => x"00013a28",
			968 => x"07002a14",
			969 => x"01000508",
			970 => x"08001804",
			971 => x"ffbf0f81",
			972 => x"00010f81",
			973 => x"00009f04",
			974 => x"ffc20f81",
			975 => x"0a003e04",
			976 => x"008b0f81",
			977 => x"ffe50f81",
			978 => x"03002c08",
			979 => x"0e007c04",
			980 => x"00200f81",
			981 => x"ff1a0f81",
			982 => x"0b001404",
			983 => x"00760f81",
			984 => x"08001904",
			985 => x"ff6a0f81",
			986 => x"00120f81",
			987 => x"0d001304",
			988 => x"00b30f81",
			989 => x"04001e04",
			990 => x"001b0f81",
			991 => x"ff8f0f81",
			992 => x"04001d1c",
			993 => x"03002710",
			994 => x"0201370c",
			995 => x"03002308",
			996 => x"03002104",
			997 => x"ffd3104d",
			998 => x"0038104d",
			999 => x"fed8104d",
			1000 => x"0023104d",
			1001 => x"0e008908",
			1002 => x"07002904",
			1003 => x"ffd7104d",
			1004 => x"00db104d",
			1005 => x"ff84104d",
			1006 => x"01000a28",
			1007 => x"00011e1c",
			1008 => x"0d001204",
			1009 => x"ff41104d",
			1010 => x"0d00130c",
			1011 => x"09002008",
			1012 => x"00009f04",
			1013 => x"fff0104d",
			1014 => x"00e5104d",
			1015 => x"ffd3104d",
			1016 => x"08001804",
			1017 => x"0072104d",
			1018 => x"05002e04",
			1019 => x"0007104d",
			1020 => x"ff40104d",
			1021 => x"05002a04",
			1022 => x"0011104d",
			1023 => x"08001b04",
			1024 => x"0114104d",
			1025 => x"0048104d",
			1026 => x"03003318",
			1027 => x"0c001404",
			1028 => x"0021104d",
			1029 => x"0f00c20c",
			1030 => x"05003904",
			1031 => x"ff25104d",
			1032 => x"05003b04",
			1033 => x"0007104d",
			1034 => x"fff8104d",
			1035 => x"0600ab04",
			1036 => x"0028104d",
			1037 => x"ffd5104d",
			1038 => x"0e006704",
			1039 => x"ff77104d",
			1040 => x"0d001604",
			1041 => x"00b8104d",
			1042 => x"ffbb104d",
			1043 => x"03003b34",
			1044 => x"09001e30",
			1045 => x"0a003424",
			1046 => x"01000b20",
			1047 => x"0c001410",
			1048 => x"0600a508",
			1049 => x"08001504",
			1050 => x"003410d1",
			1051 => x"fe8510d1",
			1052 => x"0600af04",
			1053 => x"010c10d1",
			1054 => x"ff3e10d1",
			1055 => x"0e008a08",
			1056 => x"0e007404",
			1057 => x"fedb10d1",
			1058 => x"00a410d1",
			1059 => x"0600ae04",
			1060 => x"fecd10d1",
			1061 => x"fff410d1",
			1062 => x"feae10d1",
			1063 => x"04002e08",
			1064 => x"01000704",
			1065 => x"002b10d1",
			1066 => x"015610d1",
			1067 => x"ff3010d1",
			1068 => x"fe9710d1",
			1069 => x"05004e0c",
			1070 => x"0f006f04",
			1071 => x"ff8410d1",
			1072 => x"0600a304",
			1073 => x"017c10d1",
			1074 => x"fff210d1",
			1075 => x"ff2e10d1",
			1076 => x"07002b2c",
			1077 => x"03002710",
			1078 => x"04001d04",
			1079 => x"fef51195",
			1080 => x"01000704",
			1081 => x"00ba1195",
			1082 => x"04001e04",
			1083 => x"000c1195",
			1084 => x"ffb71195",
			1085 => x"01000b18",
			1086 => x"05003508",
			1087 => x"0f008404",
			1088 => x"fff31195",
			1089 => x"01141195",
			1090 => x"0a003d08",
			1091 => x"08001804",
			1092 => x"000f1195",
			1093 => x"ff371195",
			1094 => x"05004e04",
			1095 => x"00bd1195",
			1096 => x"ffc61195",
			1097 => x"ff521195",
			1098 => x"00013d2c",
			1099 => x"09001908",
			1100 => x"01000a04",
			1101 => x"fed11195",
			1102 => x"00221195",
			1103 => x"08001808",
			1104 => x"00012504",
			1105 => x"ffab1195",
			1106 => x"00961195",
			1107 => x"0a002d0c",
			1108 => x"0e007908",
			1109 => x"06007f04",
			1110 => x"fff51195",
			1111 => x"005e1195",
			1112 => x"febd1195",
			1113 => x"09001d08",
			1114 => x"00011e04",
			1115 => x"ffcd1195",
			1116 => x"00d81195",
			1117 => x"0a004504",
			1118 => x"ff191195",
			1119 => x"00621195",
			1120 => x"0e009008",
			1121 => x"0c001704",
			1122 => x"010d1195",
			1123 => x"ffb81195",
			1124 => x"ff641195",
			1125 => x"06007104",
			1126 => x"ff131221",
			1127 => x"0e008b38",
			1128 => x"01000924",
			1129 => x"09001910",
			1130 => x"08001808",
			1131 => x"0b001304",
			1132 => x"00481221",
			1133 => x"fef81221",
			1134 => x"05002504",
			1135 => x"fff01221",
			1136 => x"00c81221",
			1137 => x"04002908",
			1138 => x"03002404",
			1139 => x"ffba1221",
			1140 => x"01071221",
			1141 => x"03003b04",
			1142 => x"ff761221",
			1143 => x"0a004504",
			1144 => x"00731221",
			1145 => x"ffec1221",
			1146 => x"0300330c",
			1147 => x"02013008",
			1148 => x"05003904",
			1149 => x"fee01221",
			1150 => x"00061221",
			1151 => x"00291221",
			1152 => x"0d001704",
			1153 => x"00cf1221",
			1154 => x"ffa71221",
			1155 => x"09001908",
			1156 => x"0a002d04",
			1157 => x"00501221",
			1158 => x"ffd11221",
			1159 => x"ff0b1221",
			1160 => x"0e008a50",
			1161 => x"0e008338",
			1162 => x"05002b14",
			1163 => x"04001a0c",
			1164 => x"04001804",
			1165 => x"ff6d12dd",
			1166 => x"0a002704",
			1167 => x"fff412dd",
			1168 => x"00aa12dd",
			1169 => x"04002004",
			1170 => x"fefe12dd",
			1171 => x"ffee12dd",
			1172 => x"0400230c",
			1173 => x"08001c08",
			1174 => x"00011e04",
			1175 => x"002c12dd",
			1176 => x"011e12dd",
			1177 => x"ffb012dd",
			1178 => x"0a003d0c",
			1179 => x"09001b04",
			1180 => x"004312dd",
			1181 => x"08001804",
			1182 => x"000d12dd",
			1183 => x"ff1912dd",
			1184 => x"0d001204",
			1185 => x"ffa012dd",
			1186 => x"05004e04",
			1187 => x"008f12dd",
			1188 => x"ffac12dd",
			1189 => x"01000904",
			1190 => x"012512dd",
			1191 => x"03002c08",
			1192 => x"05002904",
			1193 => x"fff312dd",
			1194 => x"ff7112dd",
			1195 => x"05003504",
			1196 => x"008f12dd",
			1197 => x"0a003704",
			1198 => x"000412dd",
			1199 => x"ffd012dd",
			1200 => x"01000704",
			1201 => x"ff1012dd",
			1202 => x"05002a04",
			1203 => x"ffa912dd",
			1204 => x"09001c04",
			1205 => x"008012dd",
			1206 => x"ffce12dd",
			1207 => x"07002b30",
			1208 => x"0a002d18",
			1209 => x"0c00150c",
			1210 => x"04001d04",
			1211 => x"ff6513c1",
			1212 => x"01000b04",
			1213 => x"002413c1",
			1214 => x"fff713c1",
			1215 => x"07002904",
			1216 => x"ffc713c1",
			1217 => x"03002304",
			1218 => x"fff613c1",
			1219 => x"007d13c1",
			1220 => x"0e005d0c",
			1221 => x"08001c04",
			1222 => x"ff9713c1",
			1223 => x"0e004d04",
			1224 => x"004913c1",
			1225 => x"ffe213c1",
			1226 => x"05004e08",
			1227 => x"02010204",
			1228 => x"003b13c1",
			1229 => x"00ca13c1",
			1230 => x"fff413c1",
			1231 => x"00013d38",
			1232 => x"02012b2c",
			1233 => x"00012e20",
			1234 => x"0f00b610",
			1235 => x"0f00a708",
			1236 => x"01000c04",
			1237 => x"ff7613c1",
			1238 => x"002e13c1",
			1239 => x"09001d04",
			1240 => x"008713c1",
			1241 => x"ffdf13c1",
			1242 => x"03002f08",
			1243 => x"05003004",
			1244 => x"ff2013c1",
			1245 => x"fffc13c1",
			1246 => x"03003104",
			1247 => x"001013c1",
			1248 => x"ffee13c1",
			1249 => x"01000904",
			1250 => x"00ad13c1",
			1251 => x"03003404",
			1252 => x"ff6d13c1",
			1253 => x"000e13c1",
			1254 => x"05003104",
			1255 => x"ff2e13c1",
			1256 => x"05003b04",
			1257 => x"001513c1",
			1258 => x"fff413c1",
			1259 => x"0e009008",
			1260 => x"08001c04",
			1261 => x"00b313c1",
			1262 => x"ffe213c1",
			1263 => x"ff8a13c1",
			1264 => x"05002708",
			1265 => x"03002c04",
			1266 => x"ff0c1455",
			1267 => x"001a1455",
			1268 => x"08001608",
			1269 => x"09001904",
			1270 => x"ff421455",
			1271 => x"00851455",
			1272 => x"01000a20",
			1273 => x"07002c10",
			1274 => x"03002604",
			1275 => x"ffeb1455",
			1276 => x"0f00b808",
			1277 => x"0d001204",
			1278 => x"ff781455",
			1279 => x"008a1455",
			1280 => x"013b1455",
			1281 => x"00013a0c",
			1282 => x"08001904",
			1283 => x"001e1455",
			1284 => x"03003104",
			1285 => x"fefe1455",
			1286 => x"ffe41455",
			1287 => x"008c1455",
			1288 => x"03003310",
			1289 => x"0c001404",
			1290 => x"ffed1455",
			1291 => x"05003904",
			1292 => x"ff361455",
			1293 => x"05003a04",
			1294 => x"000b1455",
			1295 => x"fff31455",
			1296 => x"0e006704",
			1297 => x"ff641455",
			1298 => x"0d001604",
			1299 => x"00c71455",
			1300 => x"ffb71455",
			1301 => x"0e008a54",
			1302 => x"0d001330",
			1303 => x"0e008228",
			1304 => x"09001914",
			1305 => x"0b001208",
			1306 => x"0b001104",
			1307 => x"ffde1521",
			1308 => x"003a1521",
			1309 => x"08001504",
			1310 => x"000f1521",
			1311 => x"08001804",
			1312 => x"ff7f1521",
			1313 => x"000d1521",
			1314 => x"0a002a08",
			1315 => x"09001a04",
			1316 => x"00141521",
			1317 => x"ffb31521",
			1318 => x"09002008",
			1319 => x"00009f04",
			1320 => x"fff61521",
			1321 => x"00751521",
			1322 => x"ffe21521",
			1323 => x"01000904",
			1324 => x"009b1521",
			1325 => x"00041521",
			1326 => x"08001808",
			1327 => x"06006704",
			1328 => x"fff81521",
			1329 => x"00391521",
			1330 => x"03002c04",
			1331 => x"ff8d1521",
			1332 => x"00010a0c",
			1333 => x"0a004504",
			1334 => x"ff901521",
			1335 => x"05004e04",
			1336 => x"00191521",
			1337 => x"fff31521",
			1338 => x"0f00b908",
			1339 => x"03003404",
			1340 => x"00601521",
			1341 => x"fff51521",
			1342 => x"ffea1521",
			1343 => x"0b001308",
			1344 => x"0f00da04",
			1345 => x"00241521",
			1346 => x"fffa1521",
			1347 => x"01000904",
			1348 => x"ff8a1521",
			1349 => x"01000b04",
			1350 => x"00091521",
			1351 => x"ffec1521",
			1352 => x"0100051c",
			1353 => x"08001b14",
			1354 => x"09001908",
			1355 => x"0c001404",
			1356 => x"fe7e1605",
			1357 => x"ffee1605",
			1358 => x"09001b04",
			1359 => x"00d61605",
			1360 => x"04001c04",
			1361 => x"00461605",
			1362 => x"fe961605",
			1363 => x"09002004",
			1364 => x"01151605",
			1365 => x"ffbb1605",
			1366 => x"08001928",
			1367 => x"01000b24",
			1368 => x"04001d10",
			1369 => x"04001a0c",
			1370 => x"04001808",
			1371 => x"0d001304",
			1372 => x"ff2a1605",
			1373 => x"00191605",
			1374 => x"01811605",
			1375 => x"ff4a1605",
			1376 => x"04003610",
			1377 => x"02012d08",
			1378 => x"00011204",
			1379 => x"00891605",
			1380 => x"01a21605",
			1381 => x"0e008504",
			1382 => x"011c1605",
			1383 => x"ff951605",
			1384 => x"ff101605",
			1385 => x"feb41605",
			1386 => x"03002c10",
			1387 => x"00014208",
			1388 => x"0a003204",
			1389 => x"fe691605",
			1390 => x"00721605",
			1391 => x"00014704",
			1392 => x"012e1605",
			1393 => x"ff0a1605",
			1394 => x"09001c08",
			1395 => x"08001c04",
			1396 => x"014e1605",
			1397 => x"ff051605",
			1398 => x"03003308",
			1399 => x"0b001604",
			1400 => x"ffba1605",
			1401 => x"fea51605",
			1402 => x"0e006708",
			1403 => x"0e004d04",
			1404 => x"00ed1605",
			1405 => x"fe981605",
			1406 => x"0d001604",
			1407 => x"012c1605",
			1408 => x"fef91605",
			1409 => x"06007104",
			1410 => x"ff0a1691",
			1411 => x"0e008b38",
			1412 => x"00013d30",
			1413 => x"0e007e14",
			1414 => x"02012110",
			1415 => x"06007408",
			1416 => x"0c001b04",
			1417 => x"00f81691",
			1418 => x"fffb1691",
			1419 => x"04001904",
			1420 => x"00741691",
			1421 => x"ff6b1691",
			1422 => x"01231691",
			1423 => x"04002010",
			1424 => x"02011f08",
			1425 => x"0a002c04",
			1426 => x"ffad1691",
			1427 => x"00ab1691",
			1428 => x"0e008304",
			1429 => x"feaf1691",
			1430 => x"00021691",
			1431 => x"00013808",
			1432 => x"01000d04",
			1433 => x"00f31691",
			1434 => x"ffa31691",
			1435 => x"ffb11691",
			1436 => x"08001c04",
			1437 => x"011a1691",
			1438 => x"ff9a1691",
			1439 => x"09001908",
			1440 => x"0a002d04",
			1441 => x"00521691",
			1442 => x"ffcd1691",
			1443 => x"ff011691",
			1444 => x"01000d58",
			1445 => x"01000308",
			1446 => x"0d001104",
			1447 => x"fe491747",
			1448 => x"ffd21747",
			1449 => x"00012f30",
			1450 => x"0a00341c",
			1451 => x"0e008010",
			1452 => x"04001808",
			1453 => x"03002704",
			1454 => x"febd1747",
			1455 => x"01311747",
			1456 => x"0d001404",
			1457 => x"fe631747",
			1458 => x"ff181747",
			1459 => x"0c001404",
			1460 => x"fe2f1747",
			1461 => x"01000a04",
			1462 => x"016e1747",
			1463 => x"feac1747",
			1464 => x"05004e10",
			1465 => x"01000708",
			1466 => x"01000404",
			1467 => x"01531747",
			1468 => x"ff331747",
			1469 => x"04003804",
			1470 => x"015a1747",
			1471 => x"fef31747",
			1472 => x"feac1747",
			1473 => x"07002c0c",
			1474 => x"0f00c704",
			1475 => x"01b21747",
			1476 => x"0f00cc04",
			1477 => x"ff881747",
			1478 => x"012c1747",
			1479 => x"00013a08",
			1480 => x"00013504",
			1481 => x"00921747",
			1482 => x"fe721747",
			1483 => x"0e009008",
			1484 => x"0d001304",
			1485 => x"016f1747",
			1486 => x"00181747",
			1487 => x"fea71747",
			1488 => x"fe761747",
			1489 => x"09001d20",
			1490 => x"00010708",
			1491 => x"03003104",
			1492 => x"fe5d17a9",
			1493 => x"ff9c17a9",
			1494 => x"01000b14",
			1495 => x"05002504",
			1496 => x"fe6417a9",
			1497 => x"0e008a0c",
			1498 => x"03002604",
			1499 => x"019817a9",
			1500 => x"0c001404",
			1501 => x"022317a9",
			1502 => x"037a17a9",
			1503 => x"001b17a9",
			1504 => x"fe4f17a9",
			1505 => x"0c001a10",
			1506 => x"0a003d04",
			1507 => x"fe5d17a9",
			1508 => x"01000908",
			1509 => x"04004304",
			1510 => x"fe5f17a9",
			1511 => x"00e817a9",
			1512 => x"02fc17a9",
			1513 => x"fe5b17a9",
			1514 => x"00011e20",
			1515 => x"0a003d14",
			1516 => x"08001504",
			1517 => x"0009183d",
			1518 => x"0c00150c",
			1519 => x"07002604",
			1520 => x"0013183d",
			1521 => x"0c001404",
			1522 => x"ffe6183d",
			1523 => x"0004183d",
			1524 => x"ff95183d",
			1525 => x"01000904",
			1526 => x"ffc8183d",
			1527 => x"09002104",
			1528 => x"0045183d",
			1529 => x"ffeb183d",
			1530 => x"0e008a18",
			1531 => x"0100090c",
			1532 => x"0c001404",
			1533 => x"ffee183d",
			1534 => x"05002704",
			1535 => x"ffe7183d",
			1536 => x"00b1183d",
			1537 => x"0f00b904",
			1538 => x"0028183d",
			1539 => x"00013f04",
			1540 => x"ff95183d",
			1541 => x"000e183d",
			1542 => x"0b001308",
			1543 => x"0f00e104",
			1544 => x"001f183d",
			1545 => x"fffc183d",
			1546 => x"01000904",
			1547 => x"ff9e183d",
			1548 => x"01000b04",
			1549 => x"0009183d",
			1550 => x"fff3183d",
			1551 => x"05002708",
			1552 => x"03002c04",
			1553 => x"fe8e1891",
			1554 => x"009f1891",
			1555 => x"00013d1c",
			1556 => x"0f00c718",
			1557 => x"0d001614",
			1558 => x"00013710",
			1559 => x"0a002d08",
			1560 => x"08001804",
			1561 => x"005d1891",
			1562 => x"fed51891",
			1563 => x"01000504",
			1564 => x"ff681891",
			1565 => x"00981891",
			1566 => x"01181891",
			1567 => x"feb81891",
			1568 => x"fe621891",
			1569 => x"07002f04",
			1570 => x"01771891",
			1571 => x"fecc1891",
			1572 => x"09001d24",
			1573 => x"00010708",
			1574 => x"03003104",
			1575 => x"fe5e18fd",
			1576 => x"ffb318fd",
			1577 => x"01000b18",
			1578 => x"05002504",
			1579 => x"fe6718fd",
			1580 => x"0e008a10",
			1581 => x"0a002d08",
			1582 => x"0d001204",
			1583 => x"028f18fd",
			1584 => x"002018fd",
			1585 => x"0d001204",
			1586 => x"026f18fd",
			1587 => x"037118fd",
			1588 => x"000b18fd",
			1589 => x"fe5218fd",
			1590 => x"0c001a10",
			1591 => x"0a003d04",
			1592 => x"fe5f18fd",
			1593 => x"05004e08",
			1594 => x"08001b04",
			1595 => x"ffff18fd",
			1596 => x"03c018fd",
			1597 => x"fe6218fd",
			1598 => x"fe5d18fd",
			1599 => x"09001d28",
			1600 => x"00010a08",
			1601 => x"03003104",
			1602 => x"fe611971",
			1603 => x"00151971",
			1604 => x"0e008a18",
			1605 => x"03002204",
			1606 => x"fe691971",
			1607 => x"01000b10",
			1608 => x"0a002d08",
			1609 => x"0d001204",
			1610 => x"02151971",
			1611 => x"00731971",
			1612 => x"0f00c704",
			1613 => x"028b1971",
			1614 => x"02041971",
			1615 => x"ff8c1971",
			1616 => x"07002e04",
			1617 => x"00791971",
			1618 => x"fe271971",
			1619 => x"0c001a10",
			1620 => x"0a003d04",
			1621 => x"fe621971",
			1622 => x"0e006508",
			1623 => x"0000b004",
			1624 => x"01461971",
			1625 => x"fe5a1971",
			1626 => x"03af1971",
			1627 => x"fe601971",
			1628 => x"0c001a28",
			1629 => x"0600670c",
			1630 => x"08001c04",
			1631 => x"fe6719c5",
			1632 => x"05004704",
			1633 => x"fe8119c5",
			1634 => x"01a319c5",
			1635 => x"0e009018",
			1636 => x"05002504",
			1637 => x"fe7419c5",
			1638 => x"01000d10",
			1639 => x"05004c08",
			1640 => x"09001e04",
			1641 => x"00f319c5",
			1642 => x"fe5019c5",
			1643 => x"05005404",
			1644 => x"03c819c5",
			1645 => x"fec719c5",
			1646 => x"fe6719c5",
			1647 => x"fe5719c5",
			1648 => x"fe6819c5",
			1649 => x"04001d1c",
			1650 => x"0300270c",
			1651 => x"0a002808",
			1652 => x"0a002704",
			1653 => x"fff41a59",
			1654 => x"000e1a59",
			1655 => x"ff8a1a59",
			1656 => x"09001a08",
			1657 => x"0600bd04",
			1658 => x"00331a59",
			1659 => x"fffc1a59",
			1660 => x"0600a004",
			1661 => x"00031a59",
			1662 => x"ffe91a59",
			1663 => x"08001c20",
			1664 => x"0d00151c",
			1665 => x"0a002a08",
			1666 => x"04002004",
			1667 => x"ffcf1a59",
			1668 => x"000e1a59",
			1669 => x"01000b10",
			1670 => x"0e006f08",
			1671 => x"05004c04",
			1672 => x"ffc41a59",
			1673 => x"00371a59",
			1674 => x"0e008a04",
			1675 => x"00b41a59",
			1676 => x"fff51a59",
			1677 => x"ffd91a59",
			1678 => x"ffd01a59",
			1679 => x"0a003704",
			1680 => x"ffa41a59",
			1681 => x"0c001a08",
			1682 => x"0e006704",
			1683 => x"fffe1a59",
			1684 => x"00281a59",
			1685 => x"ffec1a59",
			1686 => x"05002c28",
			1687 => x"00014220",
			1688 => x"0d001110",
			1689 => x"0100070c",
			1690 => x"09001908",
			1691 => x"0d000e04",
			1692 => x"002f1af5",
			1693 => x"ff6e1af5",
			1694 => x"00341af5",
			1695 => x"006c1af5",
			1696 => x"08001604",
			1697 => x"002f1af5",
			1698 => x"07002a08",
			1699 => x"03002704",
			1700 => x"ffe01af5",
			1701 => x"003b1af5",
			1702 => x"ff2c1af5",
			1703 => x"0f00d404",
			1704 => x"007a1af5",
			1705 => x"ffba1af5",
			1706 => x"08001c18",
			1707 => x"0f006f04",
			1708 => x"ffa71af5",
			1709 => x"0d001510",
			1710 => x"01000508",
			1711 => x"07002b04",
			1712 => x"00431af5",
			1713 => x"ffc41af5",
			1714 => x"04003704",
			1715 => x"00b71af5",
			1716 => x"ffeb1af5",
			1717 => x"ffbf1af5",
			1718 => x"0a003704",
			1719 => x"ff7b1af5",
			1720 => x"08001f08",
			1721 => x"04003904",
			1722 => x"005f1af5",
			1723 => x"ffef1af5",
			1724 => x"ffde1af5",
			1725 => x"08001c2c",
			1726 => x"02012f24",
			1727 => x"02012b20",
			1728 => x"00012f18",
			1729 => x"0b00150c",
			1730 => x"0d000e04",
			1731 => x"00381b79",
			1732 => x"0a003404",
			1733 => x"ff611b79",
			1734 => x"002f1b79",
			1735 => x"00010a08",
			1736 => x"03003b04",
			1737 => x"ffa81b79",
			1738 => x"00251b79",
			1739 => x"006f1b79",
			1740 => x"04001f04",
			1741 => x"00051b79",
			1742 => x"00931b79",
			1743 => x"ff8f1b79",
			1744 => x"05002704",
			1745 => x"ffcd1b79",
			1746 => x"009e1b79",
			1747 => x"03003308",
			1748 => x"05003e04",
			1749 => x"ff791b79",
			1750 => x"00051b79",
			1751 => x"0c001a0c",
			1752 => x"0a003704",
			1753 => x"fff51b79",
			1754 => x"01000904",
			1755 => x"fffa1b79",
			1756 => x"003d1b79",
			1757 => x"ffe21b79",
			1758 => x"01000b3c",
			1759 => x"07002b1c",
			1760 => x"00012214",
			1761 => x"0a003408",
			1762 => x"08001504",
			1763 => x"00571c05",
			1764 => x"fe6e1c05",
			1765 => x"01000908",
			1766 => x"06007204",
			1767 => x"feb21c05",
			1768 => x"00bf1c05",
			1769 => x"01781c05",
			1770 => x"0f00c204",
			1771 => x"01b01c05",
			1772 => x"006f1c05",
			1773 => x"00013d18",
			1774 => x"02012c14",
			1775 => x"00012d0c",
			1776 => x"0c001404",
			1777 => x"fe2f1c05",
			1778 => x"09001c04",
			1779 => x"00b51c05",
			1780 => x"fe9d1c05",
			1781 => x"01000904",
			1782 => x"00f61c05",
			1783 => x"fe901c05",
			1784 => x"fedc1c05",
			1785 => x"0e008b04",
			1786 => x"01821c05",
			1787 => x"00151c05",
			1788 => x"07003104",
			1789 => x"fe6a1c05",
			1790 => x"07003204",
			1791 => x"01111c05",
			1792 => x"febe1c05",
			1793 => x"0a003d3c",
			1794 => x"00011f14",
			1795 => x"0c00150c",
			1796 => x"08001904",
			1797 => x"ff3e1ca1",
			1798 => x"0a002d04",
			1799 => x"ffd81ca1",
			1800 => x"00a31ca1",
			1801 => x"08001804",
			1802 => x"ff831ca1",
			1803 => x"fea61ca1",
			1804 => x"0e007e08",
			1805 => x"00012a04",
			1806 => x"ff531ca1",
			1807 => x"01171ca1",
			1808 => x"00013d14",
			1809 => x"0a002d08",
			1810 => x"07002e04",
			1811 => x"fe8b1ca1",
			1812 => x"00b31ca1",
			1813 => x"0f00c708",
			1814 => x"0f00c004",
			1815 => x"ffb31ca1",
			1816 => x"01351ca1",
			1817 => x"febe1ca1",
			1818 => x"0e009008",
			1819 => x"08001c04",
			1820 => x"01291ca1",
			1821 => x"ff511ca1",
			1822 => x"ff0c1ca1",
			1823 => x"09002110",
			1824 => x"08001b08",
			1825 => x"08001804",
			1826 => x"00a21ca1",
			1827 => x"ff401ca1",
			1828 => x"05004e04",
			1829 => x"01471ca1",
			1830 => x"ffc81ca1",
			1831 => x"ff361ca1",
			1832 => x"0e008a40",
			1833 => x"0001071c",
			1834 => x"0700260c",
			1835 => x"00009f04",
			1836 => x"ffe71d45",
			1837 => x"08001b04",
			1838 => x"fff71d45",
			1839 => x"00341d45",
			1840 => x"05004c04",
			1841 => x"ff8a1d45",
			1842 => x"01000904",
			1843 => x"ffd81d45",
			1844 => x"05004f04",
			1845 => x"003a1d45",
			1846 => x"fff21d45",
			1847 => x"0c001408",
			1848 => x"0600a504",
			1849 => x"ff971d45",
			1850 => x"00231d45",
			1851 => x"01000b10",
			1852 => x"08001c0c",
			1853 => x"03002608",
			1854 => x"0d001204",
			1855 => x"002f1d45",
			1856 => x"ffc71d45",
			1857 => x"00ae1d45",
			1858 => x"ffd21d45",
			1859 => x"07003104",
			1860 => x"ffbd1d45",
			1861 => x"05003404",
			1862 => x"00191d45",
			1863 => x"fff91d45",
			1864 => x"0b001308",
			1865 => x"01000c04",
			1866 => x"000d1d45",
			1867 => x"fffc1d45",
			1868 => x"01000904",
			1869 => x"ff961d45",
			1870 => x"01000b04",
			1871 => x"000a1d45",
			1872 => x"ffef1d45",
			1873 => x"01000a34",
			1874 => x"01000308",
			1875 => x"0d001104",
			1876 => x"fe8a1dd9",
			1877 => x"003e1dd9",
			1878 => x"06009b14",
			1879 => x"0a003104",
			1880 => x"fea31dd9",
			1881 => x"0100090c",
			1882 => x"0e007108",
			1883 => x"0c001604",
			1884 => x"00d51dd9",
			1885 => x"fea81dd9",
			1886 => x"012f1dd9",
			1887 => x"01041dd9",
			1888 => x"07002a04",
			1889 => x"01791dd9",
			1890 => x"0b001408",
			1891 => x"03002904",
			1892 => x"ffef1dd9",
			1893 => x"017d1dd9",
			1894 => x"04001d04",
			1895 => x"fede1dd9",
			1896 => x"00013404",
			1897 => x"ff931dd9",
			1898 => x"00e81dd9",
			1899 => x"0d001208",
			1900 => x"08001904",
			1901 => x"00ef1dd9",
			1902 => x"ff701dd9",
			1903 => x"0b001308",
			1904 => x"0600b304",
			1905 => x"ff3f1dd9",
			1906 => x"00711dd9",
			1907 => x"0c001404",
			1908 => x"ffd11dd9",
			1909 => x"fe8a1dd9",
			1910 => x"0e008a44",
			1911 => x"00011e28",
			1912 => x"0a003d10",
			1913 => x"0c00150c",
			1914 => x"08001804",
			1915 => x"ffbc1e7d",
			1916 => x"07002504",
			1917 => x"fff61e7d",
			1918 => x"004d1e7d",
			1919 => x"ff5f1e7d",
			1920 => x"0100090c",
			1921 => x"04004304",
			1922 => x"ff771e7d",
			1923 => x"08001b04",
			1924 => x"fff11e7d",
			1925 => x"004f1e7d",
			1926 => x"04003808",
			1927 => x"01000e04",
			1928 => x"00971e7d",
			1929 => x"fff71e7d",
			1930 => x"ffca1e7d",
			1931 => x"05002b10",
			1932 => x"0d001004",
			1933 => x"00851e7d",
			1934 => x"0600ab08",
			1935 => x"07002b04",
			1936 => x"00091e7d",
			1937 => x"ff231e7d",
			1938 => x"00691e7d",
			1939 => x"08001c04",
			1940 => x"01051e7d",
			1941 => x"03003104",
			1942 => x"ff741e7d",
			1943 => x"00401e7d",
			1944 => x"01000904",
			1945 => x"ff4f1e7d",
			1946 => x"09001a08",
			1947 => x"0f00d404",
			1948 => x"004b1e7d",
			1949 => x"fff11e7d",
			1950 => x"ffc01e7d",
			1951 => x"0c00141c",
			1952 => x"0600a510",
			1953 => x"08001504",
			1954 => x"00271f29",
			1955 => x"0d001308",
			1956 => x"07002804",
			1957 => x"ffc91f29",
			1958 => x"fe801f29",
			1959 => x"00431f29",
			1960 => x"09001908",
			1961 => x"08001b04",
			1962 => x"01271f29",
			1963 => x"ffb31f29",
			1964 => x"ff631f29",
			1965 => x"0e008a30",
			1966 => x"01000918",
			1967 => x"0e00740c",
			1968 => x"04004304",
			1969 => x"feda1f29",
			1970 => x"08001b04",
			1971 => x"ffe01f29",
			1972 => x"00ee1f29",
			1973 => x"0f00c608",
			1974 => x"05002704",
			1975 => x"ff5a1f29",
			1976 => x"01651f29",
			1977 => x"00171f29",
			1978 => x"05003108",
			1979 => x"0f00c604",
			1980 => x"fe961f29",
			1981 => x"00561f29",
			1982 => x"0d00160c",
			1983 => x"04003808",
			1984 => x"00009f04",
			1985 => x"ffbc1f29",
			1986 => x"01111f29",
			1987 => x"ff741f29",
			1988 => x"ff411f29",
			1989 => x"01000904",
			1990 => x"fedb1f29",
			1991 => x"09001b04",
			1992 => x"00b01f29",
			1993 => x"ff691f29",
			1994 => x"0f006f04",
			1995 => x"fe751f9d",
			1996 => x"0e008a28",
			1997 => x"0c00140c",
			1998 => x"0d001208",
			1999 => x"0f00be04",
			2000 => x"fe021f9d",
			2001 => x"ffe31f9d",
			2002 => x"014d1f9d",
			2003 => x"0800180c",
			2004 => x"0b001404",
			2005 => x"00f71f9d",
			2006 => x"03003d04",
			2007 => x"02001f9d",
			2008 => x"ff471f9d",
			2009 => x"07002904",
			2010 => x"fe871f9d",
			2011 => x"01000404",
			2012 => x"01ae1f9d",
			2013 => x"03002c04",
			2014 => x"ff3b1f9d",
			2015 => x"00931f9d",
			2016 => x"0b00140c",
			2017 => x"09001904",
			2018 => x"feeb1f9d",
			2019 => x"0f00d804",
			2020 => x"00b61f9d",
			2021 => x"ff841f9d",
			2022 => x"fe661f9d",
			2023 => x"0a003d38",
			2024 => x"00011f10",
			2025 => x"0c00150c",
			2026 => x"08001904",
			2027 => x"ff362031",
			2028 => x"0a002d04",
			2029 => x"ffd72031",
			2030 => x"00aa2031",
			2031 => x"febb2031",
			2032 => x"0e007e08",
			2033 => x"00012a04",
			2034 => x"ff482031",
			2035 => x"01232031",
			2036 => x"00013d14",
			2037 => x"07002b04",
			2038 => x"007f2031",
			2039 => x"0600ae08",
			2040 => x"03002f04",
			2041 => x"fedc2031",
			2042 => x"00912031",
			2043 => x"04002004",
			2044 => x"ff802031",
			2045 => x"00e52031",
			2046 => x"0e009008",
			2047 => x"08001c04",
			2048 => x"01352031",
			2049 => x"ff472031",
			2050 => x"ff052031",
			2051 => x"09002110",
			2052 => x"0d001204",
			2053 => x"ff672031",
			2054 => x"05004e08",
			2055 => x"0f006f04",
			2056 => x"00742031",
			2057 => x"015c2031",
			2058 => x"ff982031",
			2059 => x"ff2d2031",
			2060 => x"0d001338",
			2061 => x"04001d10",
			2062 => x"0300270c",
			2063 => x"03002308",
			2064 => x"03002104",
			2065 => x"fff320cd",
			2066 => x"001f20cd",
			2067 => x"ff5120cd",
			2068 => x"001820cd",
			2069 => x"0f00c420",
			2070 => x"07002b14",
			2071 => x"01000a10",
			2072 => x"0c001608",
			2073 => x"07002504",
			2074 => x"fff620cd",
			2075 => x"00a620cd",
			2076 => x"03003504",
			2077 => x"ffad20cd",
			2078 => x"005920cd",
			2079 => x"ffc520cd",
			2080 => x"04002204",
			2081 => x"ff8420cd",
			2082 => x"00011404",
			2083 => x"ffd820cd",
			2084 => x"004420cd",
			2085 => x"01000704",
			2086 => x"002020cd",
			2087 => x"00af20cd",
			2088 => x"08001804",
			2089 => x"005c20cd",
			2090 => x"0b001408",
			2091 => x"03002c04",
			2092 => x"ffde20cd",
			2093 => x"003b20cd",
			2094 => x"0a004504",
			2095 => x"ff3920cd",
			2096 => x"03004004",
			2097 => x"002620cd",
			2098 => x"ffe720cd",
			2099 => x"0d001624",
			2100 => x"05002504",
			2101 => x"fe742119",
			2102 => x"0e00901c",
			2103 => x"00009f04",
			2104 => x"fe822119",
			2105 => x"0c001408",
			2106 => x"0600a504",
			2107 => x"fee12119",
			2108 => x"01692119",
			2109 => x"08001808",
			2110 => x"09001904",
			2111 => x"00632119",
			2112 => x"01e22119",
			2113 => x"0d001304",
			2114 => x"00f32119",
			2115 => x"ffe32119",
			2116 => x"fe6e2119",
			2117 => x"fe6c2119",
			2118 => x"0a002c18",
			2119 => x"08001504",
			2120 => x"007621bd",
			2121 => x"05002a0c",
			2122 => x"0d001404",
			2123 => x"fef021bd",
			2124 => x"0f00ba04",
			2125 => x"fff121bd",
			2126 => x"004f21bd",
			2127 => x"04001e04",
			2128 => x"008821bd",
			2129 => x"ff9021bd",
			2130 => x"0d001524",
			2131 => x"01000b20",
			2132 => x"0100050c",
			2133 => x"0d001208",
			2134 => x"0a003704",
			2135 => x"ff4821bd",
			2136 => x"000b21bd",
			2137 => x"007421bd",
			2138 => x"04003610",
			2139 => x"0e008b08",
			2140 => x"00010704",
			2141 => x"002e21bd",
			2142 => x"010121bd",
			2143 => x"0c001504",
			2144 => x"004621bd",
			2145 => x"ff9921bd",
			2146 => x"ff8621bd",
			2147 => x"ff6321bd",
			2148 => x"0a004510",
			2149 => x"0e008708",
			2150 => x"0c001704",
			2151 => x"000121bd",
			2152 => x"ff4a21bd",
			2153 => x"0e008a04",
			2154 => x"001f21bd",
			2155 => x"ffdd21bd",
			2156 => x"03004104",
			2157 => x"004921bd",
			2158 => x"ffe221bd",
			2159 => x"07002b28",
			2160 => x"02011620",
			2161 => x"0a003d14",
			2162 => x"08001504",
			2163 => x"00082269",
			2164 => x"07002608",
			2165 => x"07002504",
			2166 => x"fff02269",
			2167 => x"000d2269",
			2168 => x"03003504",
			2169 => x"ff982269",
			2170 => x"00042269",
			2171 => x"00009f04",
			2172 => x"fff22269",
			2173 => x"05004e04",
			2174 => x"004c2269",
			2175 => x"fff72269",
			2176 => x"01000804",
			2177 => x"00802269",
			2178 => x"fff62269",
			2179 => x"02012f28",
			2180 => x"0600a114",
			2181 => x"0f00a70c",
			2182 => x"01000c04",
			2183 => x"ffbb2269",
			2184 => x"01000d04",
			2185 => x"00142269",
			2186 => x"fff92269",
			2187 => x"01000b04",
			2188 => x"003c2269",
			2189 => x"fff42269",
			2190 => x"07002e04",
			2191 => x"ff782269",
			2192 => x"0700320c",
			2193 => x"08001f08",
			2194 => x"04001d04",
			2195 => x"fffa2269",
			2196 => x"00372269",
			2197 => x"fff72269",
			2198 => x"ffec2269",
			2199 => x"07002f04",
			2200 => x"00682269",
			2201 => x"ffcf2269",
			2202 => x"05002c24",
			2203 => x"0201301c",
			2204 => x"0d000e04",
			2205 => x"00122325",
			2206 => x"0300270c",
			2207 => x"03002308",
			2208 => x"03002104",
			2209 => x"fff52325",
			2210 => x"00042325",
			2211 => x"ff6f2325",
			2212 => x"04001a04",
			2213 => x"00232325",
			2214 => x"0e008104",
			2215 => x"ffc62325",
			2216 => x"001c2325",
			2217 => x"0f00d404",
			2218 => x"00452325",
			2219 => x"ffcd2325",
			2220 => x"05003514",
			2221 => x"0e008a0c",
			2222 => x"09001d08",
			2223 => x"0000e704",
			2224 => x"fffc2325",
			2225 => x"008a2325",
			2226 => x"fff52325",
			2227 => x"00013f04",
			2228 => x"ffdd2325",
			2229 => x"00042325",
			2230 => x"03003b1c",
			2231 => x"0201020c",
			2232 => x"0e004d08",
			2233 => x"06005204",
			2234 => x"fff72325",
			2235 => x"00142325",
			2236 => x"ff962325",
			2237 => x"08001c04",
			2238 => x"00372325",
			2239 => x"0a003b04",
			2240 => x"ffcf2325",
			2241 => x"03003404",
			2242 => x"000a2325",
			2243 => x"fffd2325",
			2244 => x"05004e08",
			2245 => x"0f006f04",
			2246 => x"fff22325",
			2247 => x"00562325",
			2248 => x"ffe22325",
			2249 => x"0c001a34",
			2250 => x"06006710",
			2251 => x"08001c04",
			2252 => x"fe602391",
			2253 => x"0d001308",
			2254 => x"00005e04",
			2255 => x"fed02391",
			2256 => x"03b12391",
			2257 => x"fe742391",
			2258 => x"0e009020",
			2259 => x"0300240c",
			2260 => x"0d001108",
			2261 => x"07002a04",
			2262 => x"fe5e2391",
			2263 => x"01f42391",
			2264 => x"fe3d2391",
			2265 => x"01000d10",
			2266 => x"0a003408",
			2267 => x"00013a04",
			2268 => x"00312391",
			2269 => x"01cc2391",
			2270 => x"05004e04",
			2271 => x"021a2391",
			2272 => x"fe8b2391",
			2273 => x"fe5e2391",
			2274 => x"fe4b2391",
			2275 => x"fe652391",
			2276 => x"05002708",
			2277 => x"03002c04",
			2278 => x"ff152425",
			2279 => x"00182425",
			2280 => x"0e008a30",
			2281 => x"0e00821c",
			2282 => x"0e007e10",
			2283 => x"00012a0c",
			2284 => x"0a003104",
			2285 => x"ff1c2425",
			2286 => x"05003704",
			2287 => x"00b92425",
			2288 => x"fffa2425",
			2289 => x"00ef2425",
			2290 => x"0b001404",
			2291 => x"003d2425",
			2292 => x"04002204",
			2293 => x"fedb2425",
			2294 => x"ffdc2425",
			2295 => x"01000904",
			2296 => x"00f52425",
			2297 => x"03002904",
			2298 => x"ff882425",
			2299 => x"05003404",
			2300 => x"00a72425",
			2301 => x"00012804",
			2302 => x"00062425",
			2303 => x"ff9e2425",
			2304 => x"04001e08",
			2305 => x"04001b04",
			2306 => x"ff872425",
			2307 => x"007d2425",
			2308 => x"00014c04",
			2309 => x"ff422425",
			2310 => x"00014e04",
			2311 => x"000d2425",
			2312 => x"fff92425",
			2313 => x"0201223c",
			2314 => x"03003b30",
			2315 => x"0b001208",
			2316 => x"0b001104",
			2317 => x"fffa24e1",
			2318 => x"005824e1",
			2319 => x"0d001418",
			2320 => x"0e008310",
			2321 => x"07002608",
			2322 => x"04002304",
			2323 => x"002624e1",
			2324 => x"ffe824e1",
			2325 => x"04001804",
			2326 => x"fffc24e1",
			2327 => x"ff2e24e1",
			2328 => x"0a003104",
			2329 => x"ffd724e1",
			2330 => x"002e24e1",
			2331 => x"00010a04",
			2332 => x"ff8824e1",
			2333 => x"09001e08",
			2334 => x"0600a204",
			2335 => x"008e24e1",
			2336 => x"ffee24e1",
			2337 => x"ffdf24e1",
			2338 => x"05004e08",
			2339 => x"0f006f04",
			2340 => x"ffda24e1",
			2341 => x"009024e1",
			2342 => x"ffc524e1",
			2343 => x"0e008a14",
			2344 => x"01000908",
			2345 => x"04001f04",
			2346 => x"004824e1",
			2347 => x"00d924e1",
			2348 => x"0a002d04",
			2349 => x"ffa824e1",
			2350 => x"05003304",
			2351 => x"003924e1",
			2352 => x"ffdf24e1",
			2353 => x"0b001304",
			2354 => x"004424e1",
			2355 => x"01000904",
			2356 => x"ff6c24e1",
			2357 => x"01000c04",
			2358 => x"000e24e1",
			2359 => x"ffe324e1",
			2360 => x"0b001838",
			2361 => x"08001c2c",
			2362 => x"05002c14",
			2363 => x"00012a04",
			2364 => x"fe402555",
			2365 => x"08001908",
			2366 => x"09001904",
			2367 => x"00152555",
			2368 => x"01c92555",
			2369 => x"09001a04",
			2370 => x"00f62555",
			2371 => x"fe812555",
			2372 => x"0d001514",
			2373 => x"06006704",
			2374 => x"fe912555",
			2375 => x"0d001208",
			2376 => x"00012d04",
			2377 => x"ff082555",
			2378 => x"01682555",
			2379 => x"05004e04",
			2380 => x"01f62555",
			2381 => x"ff2f2555",
			2382 => x"fe8e2555",
			2383 => x"0a003704",
			2384 => x"fe562555",
			2385 => x"04003404",
			2386 => x"01852555",
			2387 => x"fe872555",
			2388 => x"fe712555",
			2389 => x"04001d1c",
			2390 => x"03002710",
			2391 => x"0a002808",
			2392 => x"03002404",
			2393 => x"ffe72611",
			2394 => x"00212611",
			2395 => x"03002304",
			2396 => x"001e2611",
			2397 => x"ff402611",
			2398 => x"09001c08",
			2399 => x"08001b04",
			2400 => x"007a2611",
			2401 => x"ffeb2611",
			2402 => x"ffe12611",
			2403 => x"04001e0c",
			2404 => x"06009e04",
			2405 => x"ffe32611",
			2406 => x"07002f04",
			2407 => x"00a12611",
			2408 => x"fffb2611",
			2409 => x"07002b1c",
			2410 => x"0e005d0c",
			2411 => x"08001c04",
			2412 => x"ffba2611",
			2413 => x"07002604",
			2414 => x"00282611",
			2415 => x"ffea2611",
			2416 => x"01000a0c",
			2417 => x"06009908",
			2418 => x"06007404",
			2419 => x"005c2611",
			2420 => x"ffc82611",
			2421 => x"008c2611",
			2422 => x"fff32611",
			2423 => x"0b001404",
			2424 => x"001b2611",
			2425 => x"0e00840c",
			2426 => x"0a004504",
			2427 => x"ff772611",
			2428 => x"0200be04",
			2429 => x"00282611",
			2430 => x"ffe72611",
			2431 => x"0e008b08",
			2432 => x"01000d04",
			2433 => x"00682611",
			2434 => x"ffe92611",
			2435 => x"ff942611",
			2436 => x"0500270c",
			2437 => x"03002c04",
			2438 => x"febf26c5",
			2439 => x"03002d04",
			2440 => x"004d26c5",
			2441 => x"fff626c5",
			2442 => x"0600a32c",
			2443 => x"00011e20",
			2444 => x"0a003d10",
			2445 => x"0100060c",
			2446 => x"0b001608",
			2447 => x"0a003104",
			2448 => x"ff8426c5",
			2449 => x"00ad26c5",
			2450 => x"ff4626c5",
			2451 => x"fed526c5",
			2452 => x"05004e0c",
			2453 => x"05004c08",
			2454 => x"05004904",
			2455 => x"00f626c5",
			2456 => x"ff0326c5",
			2457 => x"014226c5",
			2458 => x"ff4e26c5",
			2459 => x"0c001504",
			2460 => x"006e26c5",
			2461 => x"09001d04",
			2462 => x"016826c5",
			2463 => x"ff9626c5",
			2464 => x"00013c18",
			2465 => x"03002c0c",
			2466 => x"04002208",
			2467 => x"0f00c304",
			2468 => x"ff6a26c5",
			2469 => x"fea326c5",
			2470 => x"008b26c5",
			2471 => x"0600ad08",
			2472 => x"09001d04",
			2473 => x"013e26c5",
			2474 => x"ffa426c5",
			2475 => x"ff4326c5",
			2476 => x"07002f08",
			2477 => x"07002b04",
			2478 => x"000626c5",
			2479 => x"015026c5",
			2480 => x"ff2826c5",
			2481 => x"0c001940",
			2482 => x"0000cf0c",
			2483 => x"08001c04",
			2484 => x"fe652749",
			2485 => x"0c001804",
			2486 => x"fe8c2749",
			2487 => x"01d82749",
			2488 => x"07002b14",
			2489 => x"0b001510",
			2490 => x"0600a008",
			2491 => x"05002c04",
			2492 => x"fe492749",
			2493 => x"00bf2749",
			2494 => x"03002404",
			2495 => x"ff6e2749",
			2496 => x"01e82749",
			2497 => x"029b2749",
			2498 => x"02012f14",
			2499 => x"0400220c",
			2500 => x"0e007e04",
			2501 => x"00af2749",
			2502 => x"0e008304",
			2503 => x"fda62749",
			2504 => x"ff4b2749",
			2505 => x"09001d04",
			2506 => x"01012749",
			2507 => x"fe7a2749",
			2508 => x"07002f08",
			2509 => x"09001a04",
			2510 => x"01dc2749",
			2511 => x"00e92749",
			2512 => x"fe6e2749",
			2513 => x"fe642749",
			2514 => x"03003b44",
			2515 => x"01000514",
			2516 => x"0c001404",
			2517 => x"feb827ed",
			2518 => x"09001b08",
			2519 => x"03002304",
			2520 => x"ff6627ed",
			2521 => x"011e27ed",
			2522 => x"0d001304",
			2523 => x"feeb27ed",
			2524 => x"001d27ed",
			2525 => x"0d001524",
			2526 => x"01000b20",
			2527 => x"0a002c10",
			2528 => x"0c001408",
			2529 => x"0c001304",
			2530 => x"fff927ed",
			2531 => x"fea527ed",
			2532 => x"08001904",
			2533 => x"00c427ed",
			2534 => x"ff8027ed",
			2535 => x"0f00c708",
			2536 => x"04003404",
			2537 => x"011027ed",
			2538 => x"fef527ed",
			2539 => x"00013d04",
			2540 => x"fe9927ed",
			2541 => x"00ca27ed",
			2542 => x"feaf27ed",
			2543 => x"0e008704",
			2544 => x"feb027ed",
			2545 => x"0600a304",
			2546 => x"00f827ed",
			2547 => x"ff4d27ed",
			2548 => x"05004e0c",
			2549 => x"0f006f04",
			2550 => x"ff8a27ed",
			2551 => x"0600a304",
			2552 => x"016b27ed",
			2553 => x"fff227ed",
			2554 => x"ff3a27ed",
			2555 => x"07002b30",
			2556 => x"0a002d18",
			2557 => x"0c00150c",
			2558 => x"04001d04",
			2559 => x"ff5f28c9",
			2560 => x"01000b04",
			2561 => x"002428c9",
			2562 => x"fff628c9",
			2563 => x"07002904",
			2564 => x"ffc528c9",
			2565 => x"03002304",
			2566 => x"fff628c9",
			2567 => x"008528c9",
			2568 => x"0e005d0c",
			2569 => x"08001c04",
			2570 => x"ff9428c9",
			2571 => x"0e004d04",
			2572 => x"004c28c9",
			2573 => x"ffe228c9",
			2574 => x"02010208",
			2575 => x"0e006604",
			2576 => x"009428c9",
			2577 => x"ffa828c9",
			2578 => x"00d528c9",
			2579 => x"00013d34",
			2580 => x"0400221c",
			2581 => x"05003418",
			2582 => x"0600ae10",
			2583 => x"0e007b08",
			2584 => x"0b001504",
			2585 => x"002128c9",
			2586 => x"ffe628c9",
			2587 => x"02011604",
			2588 => x"ffff28c9",
			2589 => x"ff2028c9",
			2590 => x"0b001404",
			2591 => x"ffd728c9",
			2592 => x"004d28c9",
			2593 => x"003f28c9",
			2594 => x"09001c04",
			2595 => x"007b28c9",
			2596 => x"01000c08",
			2597 => x"0e008004",
			2598 => x"ff4f28c9",
			2599 => x"000b28c9",
			2600 => x"01000d08",
			2601 => x"08001d04",
			2602 => x"fff028c9",
			2603 => x"006328c9",
			2604 => x"ffd928c9",
			2605 => x"0e009008",
			2606 => x"0b001504",
			2607 => x"00c128c9",
			2608 => x"fff428c9",
			2609 => x"ff8628c9",
			2610 => x"0e008a40",
			2611 => x"0600ab3c",
			2612 => x"05002b18",
			2613 => x"03002710",
			2614 => x"0d00110c",
			2615 => x"0d000f04",
			2616 => x"ff81296d",
			2617 => x"03002104",
			2618 => x"fffa296d",
			2619 => x"0052296d",
			2620 => x"fefd296d",
			2621 => x"08001b04",
			2622 => x"0093296d",
			2623 => x"ff7c296d",
			2624 => x"0d001514",
			2625 => x"08001c0c",
			2626 => x"00012d08",
			2627 => x"0d001204",
			2628 => x"ff79296d",
			2629 => x"009e296d",
			2630 => x"010a296d",
			2631 => x"0e004d04",
			2632 => x"006a296d",
			2633 => x"ff47296d",
			2634 => x"01000c04",
			2635 => x"ff65296d",
			2636 => x"01000d08",
			2637 => x"03003304",
			2638 => x"ffe3296d",
			2639 => x"0076296d",
			2640 => x"ffc6296d",
			2641 => x"00bd296d",
			2642 => x"0b001308",
			2643 => x"0f00df04",
			2644 => x"005c296d",
			2645 => x"fff0296d",
			2646 => x"01000904",
			2647 => x"ff15296d",
			2648 => x"01000b04",
			2649 => x"0027296d",
			2650 => x"ffc9296d",
			2651 => x"0f006f04",
			2652 => x"fe7929f1",
			2653 => x"0e008a30",
			2654 => x"0c00140c",
			2655 => x"0d001208",
			2656 => x"0f00be04",
			2657 => x"fe1f29f1",
			2658 => x"ffdf29f1",
			2659 => x"013129f1",
			2660 => x"08001810",
			2661 => x"05002504",
			2662 => x"ff3229f1",
			2663 => x"0b001404",
			2664 => x"00ed29f1",
			2665 => x"03003d04",
			2666 => x"01fb29f1",
			2667 => x"ff5229f1",
			2668 => x"00014110",
			2669 => x"0a003708",
			2670 => x"09001b04",
			2671 => x"005d29f1",
			2672 => x"fead29f1",
			2673 => x"0e006504",
			2674 => x"fe8529f1",
			2675 => x"013929f1",
			2676 => x"018329f1",
			2677 => x"0b00140c",
			2678 => x"09001904",
			2679 => x"fef729f1",
			2680 => x"0f00d804",
			2681 => x"00af29f1",
			2682 => x"ff8c29f1",
			2683 => x"fe7029f1",
			2684 => x"0c001944",
			2685 => x"0000cf10",
			2686 => x"08001c04",
			2687 => x"fe682a7d",
			2688 => x"08001d08",
			2689 => x"0d001304",
			2690 => x"024f2a7d",
			2691 => x"ff142a7d",
			2692 => x"fe912a7d",
			2693 => x"07002b14",
			2694 => x"04001804",
			2695 => x"fe6f2a7d",
			2696 => x"0b00150c",
			2697 => x"0e007004",
			2698 => x"fde22a7d",
			2699 => x"0a002c04",
			2700 => x"ffd22a7d",
			2701 => x"01882a7d",
			2702 => x"02532a7d",
			2703 => x"00013d14",
			2704 => x"0a00370c",
			2705 => x"0e007e04",
			2706 => x"008c2a7d",
			2707 => x"02012b04",
			2708 => x"ff6c2a7d",
			2709 => x"fe322a7d",
			2710 => x"09001d04",
			2711 => x"01fc2a7d",
			2712 => x"fe892a7d",
			2713 => x"07002f08",
			2714 => x"09001a04",
			2715 => x"01cb2a7d",
			2716 => x"01272a7d",
			2717 => x"fe742a7d",
			2718 => x"fe662a7d",
			2719 => x"08001508",
			2720 => x"09001804",
			2721 => x"ffe52b09",
			2722 => x"007e2b09",
			2723 => x"05002708",
			2724 => x"03002c04",
			2725 => x"ff572b09",
			2726 => x"00082b09",
			2727 => x"00013a2c",
			2728 => x"07002b10",
			2729 => x"01000b0c",
			2730 => x"02011608",
			2731 => x"0a003d04",
			2732 => x"ff902b09",
			2733 => x"00632b09",
			2734 => x"007e2b09",
			2735 => x"ff982b09",
			2736 => x"0600a10c",
			2737 => x"06009d08",
			2738 => x"01000c04",
			2739 => x"ff932b09",
			2740 => x"001d2b09",
			2741 => x"00752b09",
			2742 => x"03003108",
			2743 => x"0600a804",
			2744 => x"ff122b09",
			2745 => x"00092b09",
			2746 => x"0e008904",
			2747 => x"00452b09",
			2748 => x"fff52b09",
			2749 => x"0d001304",
			2750 => x"00ab2b09",
			2751 => x"04001e04",
			2752 => x"001a2b09",
			2753 => x"ff912b09",
			2754 => x"0d001644",
			2755 => x"0300240c",
			2756 => x"0d001108",
			2757 => x"0b001404",
			2758 => x"fe8a2b95",
			2759 => x"014d2b95",
			2760 => x"fe532b95",
			2761 => x"0e008a28",
			2762 => x"0c001408",
			2763 => x"0600a504",
			2764 => x"fecb2b95",
			2765 => x"012e2b95",
			2766 => x"02010210",
			2767 => x"03003808",
			2768 => x"06008e04",
			2769 => x"fe412b95",
			2770 => x"006a2b95",
			2771 => x"05004e04",
			2772 => x"01912b95",
			2773 => x"fe8f2b95",
			2774 => x"08001c08",
			2775 => x"03002c04",
			2776 => x"00cf2b95",
			2777 => x"01e72b95",
			2778 => x"03002f04",
			2779 => x"fe3a2b95",
			2780 => x"00dc2b95",
			2781 => x"0b001408",
			2782 => x"00013604",
			2783 => x"fed12b95",
			2784 => x"015d2b95",
			2785 => x"00014604",
			2786 => x"fdf62b95",
			2787 => x"00012b95",
			2788 => x"fe702b95",
			2789 => x"0d001630",
			2790 => x"05002504",
			2791 => x"fe712bf9",
			2792 => x"0e009028",
			2793 => x"07002914",
			2794 => x"05002904",
			2795 => x"fe502bf9",
			2796 => x"05003508",
			2797 => x"0000d204",
			2798 => x"feb42bf9",
			2799 => x"01d62bf9",
			2800 => x"09001f04",
			2801 => x"fe462bf9",
			2802 => x"00f52bf9",
			2803 => x"00014210",
			2804 => x"07002b08",
			2805 => x"0d001504",
			2806 => x"01652bf9",
			2807 => x"fe9b2bf9",
			2808 => x"09001904",
			2809 => x"ff1b2bf9",
			2810 => x"00962bf9",
			2811 => x"01b82bf9",
			2812 => x"fe692bf9",
			2813 => x"fe6b2bf9",
			2814 => x"0d001648",
			2815 => x"05002708",
			2816 => x"03002c04",
			2817 => x"fe6d2c8f",
			2818 => x"00f12c8f",
			2819 => x"09001c1c",
			2820 => x"08001c14",
			2821 => x"00013b10",
			2822 => x"0a003408",
			2823 => x"07002c04",
			2824 => x"00512c8f",
			2825 => x"ff0b2c8f",
			2826 => x"04002a04",
			2827 => x"01c92c8f",
			2828 => x"00ce2c8f",
			2829 => x"01962c8f",
			2830 => x"0e008604",
			2831 => x"ff632c8f",
			2832 => x"fe602c8f",
			2833 => x"0a004318",
			2834 => x"0b001508",
			2835 => x"01000804",
			2836 => x"012c2c8f",
			2837 => x"fec32c8f",
			2838 => x"0e004d08",
			2839 => x"08001c04",
			2840 => x"fefa2c8f",
			2841 => x"01cf2c8f",
			2842 => x"07003104",
			2843 => x"fe682c8f",
			2844 => x"00402c8f",
			2845 => x"08001b04",
			2846 => x"feb82c8f",
			2847 => x"03004404",
			2848 => x"029f2c8f",
			2849 => x"ff532c8f",
			2850 => x"fe742c8f",
			2851 => x"09001c28",
			2852 => x"0500270c",
			2853 => x"08001504",
			2854 => x"00202d11",
			2855 => x"03002a04",
			2856 => x"ff8a2d11",
			2857 => x"00032d11",
			2858 => x"0c001408",
			2859 => x"0600a504",
			2860 => x"ff992d11",
			2861 => x"00472d11",
			2862 => x"01000b10",
			2863 => x"00010a04",
			2864 => x"ffdb2d11",
			2865 => x"0600a504",
			2866 => x"00a92d11",
			2867 => x"0f00c904",
			2868 => x"ffbe2d11",
			2869 => x"00762d11",
			2870 => x"ffc72d11",
			2871 => x"08001808",
			2872 => x"0f006f04",
			2873 => x"ffe32d11",
			2874 => x"00332d11",
			2875 => x"0e004d08",
			2876 => x"00009f04",
			2877 => x"ffee2d11",
			2878 => x"00222d11",
			2879 => x"0a004504",
			2880 => x"ff8d2d11",
			2881 => x"0a004704",
			2882 => x"00172d11",
			2883 => x"ffea2d11",
			2884 => x"00011e1c",
			2885 => x"0a003d10",
			2886 => x"08001504",
			2887 => x"00092da5",
			2888 => x"07002608",
			2889 => x"07002504",
			2890 => x"fff02da5",
			2891 => x"000e2da5",
			2892 => x"ff922da5",
			2893 => x"01000904",
			2894 => x"ffc62da5",
			2895 => x"09002104",
			2896 => x"00482da5",
			2897 => x"ffeb2da5",
			2898 => x"0a002c10",
			2899 => x"05002a0c",
			2900 => x"0d001408",
			2901 => x"0600ad04",
			2902 => x"ff812da5",
			2903 => x"fff42da5",
			2904 => x"00182da5",
			2905 => x"00302da5",
			2906 => x"0e008a14",
			2907 => x"01000908",
			2908 => x"01000504",
			2909 => x"fffb2da5",
			2910 => x"00ab2da5",
			2911 => x"0f00b904",
			2912 => x"00292da5",
			2913 => x"02013004",
			2914 => x"ffb52da5",
			2915 => x"000c2da5",
			2916 => x"0b001408",
			2917 => x"0f00e004",
			2918 => x"00252da5",
			2919 => x"fffb2da5",
			2920 => x"ffb52da5",
			2921 => x"05002708",
			2922 => x"03002c04",
			2923 => x"fe872e01",
			2924 => x"00a22e01",
			2925 => x"00013d20",
			2926 => x"0f00c71c",
			2927 => x"02012810",
			2928 => x"0f00c10c",
			2929 => x"09001904",
			2930 => x"ff662e01",
			2931 => x"00011e04",
			2932 => x"fff92e01",
			2933 => x"01562e01",
			2934 => x"feda2e01",
			2935 => x"01000904",
			2936 => x"01932e01",
			2937 => x"0f00c404",
			2938 => x"fea62e01",
			2939 => x"00402e01",
			2940 => x"fe542e01",
			2941 => x"07002f04",
			2942 => x"017f2e01",
			2943 => x"fec32e01",
			2944 => x"09001d24",
			2945 => x"00010a08",
			2946 => x"03003104",
			2947 => x"fe602e6d",
			2948 => x"00052e6d",
			2949 => x"0e008e18",
			2950 => x"05002504",
			2951 => x"fe6e2e6d",
			2952 => x"01000b10",
			2953 => x"0a002f08",
			2954 => x"02013004",
			2955 => x"00f82e6d",
			2956 => x"03452e6d",
			2957 => x"0f00c704",
			2958 => x"02dc2e6d",
			2959 => x"01f42e6d",
			2960 => x"ff7e2e6d",
			2961 => x"fe432e6d",
			2962 => x"0c001a10",
			2963 => x"0a003d04",
			2964 => x"fe602e6d",
			2965 => x"05004e08",
			2966 => x"0f006b04",
			2967 => x"00622e6d",
			2968 => x"03a42e6d",
			2969 => x"fe672e6d",
			2970 => x"fe5f2e6d",
			2971 => x"0c001a24",
			2972 => x"0a002808",
			2973 => x"0e008504",
			2974 => x"fe462eb9",
			2975 => x"00712eb9",
			2976 => x"01000304",
			2977 => x"fdfd2eb9",
			2978 => x"0e009014",
			2979 => x"01000d10",
			2980 => x"00013a08",
			2981 => x"04002004",
			2982 => x"ffbd2eb9",
			2983 => x"00ef2eb9",
			2984 => x"08001b04",
			2985 => x"01c82eb9",
			2986 => x"00692eb9",
			2987 => x"fe6e2eb9",
			2988 => x"fe622eb9",
			2989 => x"fe692eb9",
			2990 => x"0c001a28",
			2991 => x"0a00280c",
			2992 => x"0e008508",
			2993 => x"0f00be04",
			2994 => x"fe6d2f0d",
			2995 => x"fdb82f0d",
			2996 => x"00842f0d",
			2997 => x"01000304",
			2998 => x"fdc62f0d",
			2999 => x"0e009014",
			3000 => x"01000d10",
			3001 => x"06007108",
			3002 => x"04003604",
			3003 => x"00b92f0d",
			3004 => x"fe672f0d",
			3005 => x"08001c04",
			3006 => x"01202f0d",
			3007 => x"ffb32f0d",
			3008 => x"fe6a2f0d",
			3009 => x"fe5e2f0d",
			3010 => x"fe682f0d",
			3011 => x"04001d14",
			3012 => x"0300270c",
			3013 => x"0a002808",
			3014 => x"03002404",
			3015 => x"ffe42fa1",
			3016 => x"001f2fa1",
			3017 => x"ff6a2fa1",
			3018 => x"07002e04",
			3019 => x"005a2fa1",
			3020 => x"ffd72fa1",
			3021 => x"08001c28",
			3022 => x"00012f20",
			3023 => x"0a003410",
			3024 => x"0d001308",
			3025 => x"0d001104",
			3026 => x"00122fa1",
			3027 => x"ff732fa1",
			3028 => x"03002c04",
			3029 => x"ffdf2fa1",
			3030 => x"00322fa1",
			3031 => x"06006704",
			3032 => x"ffc62fa1",
			3033 => x"0d001508",
			3034 => x"0b001804",
			3035 => x"007a2fa1",
			3036 => x"ffef2fa1",
			3037 => x"ffd82fa1",
			3038 => x"07002c04",
			3039 => x"00982fa1",
			3040 => x"00252fa1",
			3041 => x"0000c70c",
			3042 => x"00009f04",
			3043 => x"fff02fa1",
			3044 => x"04003804",
			3045 => x"00442fa1",
			3046 => x"fff62fa1",
			3047 => x"ff872fa1",
			3048 => x"08001c40",
			3049 => x"02010214",
			3050 => x"03003b0c",
			3051 => x"0c001408",
			3052 => x"08001b04",
			3053 => x"fe7a3045",
			3054 => x"02b03045",
			3055 => x"fe4f3045",
			3056 => x"05004e04",
			3057 => x"02893045",
			3058 => x"fe713045",
			3059 => x"03002714",
			3060 => x"0d00120c",
			3061 => x"04001d08",
			3062 => x"09001804",
			3063 => x"fe2a3045",
			3064 => x"00663045",
			3065 => x"022a3045",
			3066 => x"07002d04",
			3067 => x"fe0d3045",
			3068 => x"ffa83045",
			3069 => x"0e008a10",
			3070 => x"0c001404",
			3071 => x"01203045",
			3072 => x"06009f04",
			3073 => x"028d3045",
			3074 => x"0f00c104",
			3075 => x"01013045",
			3076 => x"01ff3045",
			3077 => x"0d001204",
			3078 => x"ff473045",
			3079 => x"01953045",
			3080 => x"01000608",
			3081 => x"09002004",
			3082 => x"ffe83045",
			3083 => x"feac3045",
			3084 => x"03003304",
			3085 => x"fe573045",
			3086 => x"05003704",
			3087 => x"01713045",
			3088 => x"fe633045",
			3089 => x"05002c28",
			3090 => x"03002718",
			3091 => x"04001d0c",
			3092 => x"03002308",
			3093 => x"03002104",
			3094 => x"ffb630f9",
			3095 => x"004030f9",
			3096 => x"fea530f9",
			3097 => x"0d001204",
			3098 => x"00e430f9",
			3099 => x"07002e04",
			3100 => x"feec30f9",
			3101 => x"007530f9",
			3102 => x"04001b08",
			3103 => x"00012a04",
			3104 => x"ffb630f9",
			3105 => x"00f330f9",
			3106 => x"05002a04",
			3107 => x"ff2930f9",
			3108 => x"007530f9",
			3109 => x"04002310",
			3110 => x"08001c0c",
			3111 => x"0e008508",
			3112 => x"0e007404",
			3113 => x"006a30f9",
			3114 => x"014730f9",
			3115 => x"003d30f9",
			3116 => x"ff2630f9",
			3117 => x"0a003708",
			3118 => x"09001b04",
			3119 => x"000730f9",
			3120 => x"fee330f9",
			3121 => x"04002e08",
			3122 => x"09001e04",
			3123 => x"00f930f9",
			3124 => x"ffd230f9",
			3125 => x"03003b08",
			3126 => x"0e004f04",
			3127 => x"006b30f9",
			3128 => x"fef230f9",
			3129 => x"05004e08",
			3130 => x"0f006f04",
			3131 => x"ffb530f9",
			3132 => x"00e630f9",
			3133 => x"ff8030f9",
			3134 => x"0d001330",
			3135 => x"0e008a28",
			3136 => x"00012f20",
			3137 => x"0a003410",
			3138 => x"0b001204",
			3139 => x"001f318d",
			3140 => x"0b001608",
			3141 => x"04001804",
			3142 => x"fffe318d",
			3143 => x"ff86318d",
			3144 => x"000b318d",
			3145 => x"0900200c",
			3146 => x"06005504",
			3147 => x"fff9318d",
			3148 => x"05004e04",
			3149 => x"0051318d",
			3150 => x"fffc318d",
			3151 => x"ffea318d",
			3152 => x"01000804",
			3153 => x"0076318d",
			3154 => x"fffb318d",
			3155 => x"0b001304",
			3156 => x"0010318d",
			3157 => x"ff9e318d",
			3158 => x"08001808",
			3159 => x"0f00a504",
			3160 => x"fff8318d",
			3161 => x"0031318d",
			3162 => x"0a00450c",
			3163 => x"0b001408",
			3164 => x"0c001404",
			3165 => x"ffec318d",
			3166 => x"000e318d",
			3167 => x"ff8a318d",
			3168 => x"03004004",
			3169 => x"0014318d",
			3170 => x"fff0318d",
			3171 => x"09001d24",
			3172 => x"0000e704",
			3173 => x"fe6431f9",
			3174 => x"0e00901c",
			3175 => x"05002504",
			3176 => x"fe6f31f9",
			3177 => x"0a003410",
			3178 => x"00013d08",
			3179 => x"07002c04",
			3180 => x"012431f9",
			3181 => x"ff6c31f9",
			3182 => x"05002c04",
			3183 => x"028f31f9",
			3184 => x"01e931f9",
			3185 => x"05003804",
			3186 => x"02da31f9",
			3187 => x"020931f9",
			3188 => x"fe5331f9",
			3189 => x"0c001a10",
			3190 => x"0a003d04",
			3191 => x"fe6531f9",
			3192 => x"05004e08",
			3193 => x"08001b04",
			3194 => x"fffa31f9",
			3195 => x"028f31f9",
			3196 => x"fe6a31f9",
			3197 => x"fe6231f9",
			3198 => x"0e008a38",
			3199 => x"05002c10",
			3200 => x"00012a04",
			3201 => x"fe6b3285",
			3202 => x"01000908",
			3203 => x"02012c04",
			3204 => x"00d93285",
			3205 => x"ffa53285",
			3206 => x"fec83285",
			3207 => x"05002e08",
			3208 => x"0e007404",
			3209 => x"ff0d3285",
			3210 => x"01733285",
			3211 => x"05003008",
			3212 => x"07002b04",
			3213 => x"00b73285",
			3214 => x"fef13285",
			3215 => x"0201020c",
			3216 => x"06007408",
			3217 => x"06007104",
			3218 => x"ffdd3285",
			3219 => x"019a3285",
			3220 => x"fe773285",
			3221 => x"08001c04",
			3222 => x"01933285",
			3223 => x"03003104",
			3224 => x"fe9e3285",
			3225 => x"01183285",
			3226 => x"01000704",
			3227 => x"fe643285",
			3228 => x"0e009008",
			3229 => x"09001c04",
			3230 => x"014c3285",
			3231 => x"ff4b3285",
			3232 => x"feb03285",
			3233 => x"0e008a40",
			3234 => x"0001071c",
			3235 => x"0700260c",
			3236 => x"00009f04",
			3237 => x"ffe63319",
			3238 => x"08001b04",
			3239 => x"fff63319",
			3240 => x"00353319",
			3241 => x"05004c04",
			3242 => x"ff873319",
			3243 => x"01000904",
			3244 => x"ffd63319",
			3245 => x"05004f04",
			3246 => x"003b3319",
			3247 => x"fff23319",
			3248 => x"0c001408",
			3249 => x"0600a504",
			3250 => x"ff913319",
			3251 => x"00243319",
			3252 => x"01000b10",
			3253 => x"08001c0c",
			3254 => x"03002608",
			3255 => x"0d001204",
			3256 => x"00323319",
			3257 => x"ffc53319",
			3258 => x"00b73319",
			3259 => x"ffd03319",
			3260 => x"07003104",
			3261 => x"ffba3319",
			3262 => x"05003404",
			3263 => x"001a3319",
			3264 => x"fff93319",
			3265 => x"0b001308",
			3266 => x"01000c04",
			3267 => x"000e3319",
			3268 => x"fffc3319",
			3269 => x"ff973319",
			3270 => x"02012234",
			3271 => x"0c001408",
			3272 => x"04002004",
			3273 => x"ff2333bd",
			3274 => x"004233bd",
			3275 => x"08001810",
			3276 => x"0f006f04",
			3277 => x"ffcb33bd",
			3278 => x"03002604",
			3279 => x"ffd933bd",
			3280 => x"04003704",
			3281 => x"00be33bd",
			3282 => x"fff033bd",
			3283 => x"0a004310",
			3284 => x"00010a04",
			3285 => x"ff2a33bd",
			3286 => x"0600a208",
			3287 => x"09001e04",
			3288 => x"005833bd",
			3289 => x"ffe833bd",
			3290 => x"ffb333bd",
			3291 => x"0000d008",
			3292 => x"0f007404",
			3293 => x"fff633bd",
			3294 => x"006a33bd",
			3295 => x"ffd933bd",
			3296 => x"0e008a10",
			3297 => x"01000904",
			3298 => x"00b833bd",
			3299 => x"0a002d04",
			3300 => x"ffa533bd",
			3301 => x"05003304",
			3302 => x"003b33bd",
			3303 => x"ffde33bd",
			3304 => x"0b001304",
			3305 => x"004433bd",
			3306 => x"01000904",
			3307 => x"ff6833bd",
			3308 => x"01000c04",
			3309 => x"001033bd",
			3310 => x"ffe233bd",
			3311 => x"0a002d1c",
			3312 => x"0f00c810",
			3313 => x"05002b04",
			3314 => x"fec93469",
			3315 => x"04001f04",
			3316 => x"00ee3469",
			3317 => x"0c001604",
			3318 => x"00133469",
			3319 => x"ff0a3469",
			3320 => x"0e008a04",
			3321 => x"00a43469",
			3322 => x"0b001304",
			3323 => x"00313469",
			3324 => x"ff263469",
			3325 => x"02012328",
			3326 => x"05004c20",
			3327 => x"0e006f0c",
			3328 => x"0e004d08",
			3329 => x"08001c04",
			3330 => x"ffb13469",
			3331 => x"00ae3469",
			3332 => x"febd3469",
			3333 => x"07002b04",
			3334 => x"00a13469",
			3335 => x"0f00b608",
			3336 => x"04002304",
			3337 => x"009f3469",
			3338 => x"ff813469",
			3339 => x"00012e04",
			3340 => x"fef73469",
			3341 => x"003e3469",
			3342 => x"05004e04",
			3343 => x"00f93469",
			3344 => x"ff703469",
			3345 => x"08001c08",
			3346 => x"0e008904",
			3347 => x"01603469",
			3348 => x"ffab3469",
			3349 => x"0a003b04",
			3350 => x"ff223469",
			3351 => x"03003404",
			3352 => x"002e3469",
			3353 => x"fff43469",
			3354 => x"05002708",
			3355 => x"03002c04",
			3356 => x"ff4634ed",
			3357 => x"000834ed",
			3358 => x"08001c2c",
			3359 => x"00013a20",
			3360 => x"07002b10",
			3361 => x"0e005d04",
			3362 => x"ff9f34ed",
			3363 => x"0a002d04",
			3364 => x"ffeb34ed",
			3365 => x"04002e04",
			3366 => x"00c534ed",
			3367 => x"002d34ed",
			3368 => x"0600a108",
			3369 => x"00010a04",
			3370 => x"ff8934ed",
			3371 => x"007534ed",
			3372 => x"0600a804",
			3373 => x"ff4a34ed",
			3374 => x"ffff34ed",
			3375 => x"04002004",
			3376 => x"00c734ed",
			3377 => x"04002204",
			3378 => x"ffff34ed",
			3379 => x"003034ed",
			3380 => x"0200be0c",
			3381 => x"03003804",
			3382 => x"ffe534ed",
			3383 => x"04003804",
			3384 => x"006b34ed",
			3385 => x"ffeb34ed",
			3386 => x"ff5e34ed",
			3387 => x"0e008a40",
			3388 => x"00012f2c",
			3389 => x"05002c14",
			3390 => x"0c00170c",
			3391 => x"0b001208",
			3392 => x"06005404",
			3393 => x"ffd23589",
			3394 => x"00f73589",
			3395 => x"fe7b3589",
			3396 => x"09001c04",
			3397 => x"011a3589",
			3398 => x"ff7d3589",
			3399 => x"04003814",
			3400 => x"05004c10",
			3401 => x"0e006f08",
			3402 => x"07002604",
			3403 => x"00943589",
			3404 => x"fe983589",
			3405 => x"09001e04",
			3406 => x"00f93589",
			3407 => x"ff1b3589",
			3408 => x"01703589",
			3409 => x"feca3589",
			3410 => x"0d001308",
			3411 => x"01000804",
			3412 => x"018c3589",
			3413 => x"00273589",
			3414 => x"0a002d04",
			3415 => x"feb03589",
			3416 => x"05003304",
			3417 => x"00bf3589",
			3418 => x"ffd23589",
			3419 => x"09001b0c",
			3420 => x"00013f08",
			3421 => x"0a003104",
			3422 => x"fefd3589",
			3423 => x"00873589",
			3424 => x"00a73589",
			3425 => x"feab3589",
			3426 => x"05002c28",
			3427 => x"03002718",
			3428 => x"04001d0c",
			3429 => x"03002308",
			3430 => x"03002104",
			3431 => x"ffb9363d",
			3432 => x"0039363d",
			3433 => x"fead363d",
			3434 => x"0d001204",
			3435 => x"00d8363d",
			3436 => x"07002e04",
			3437 => x"fef5363d",
			3438 => x"006c363d",
			3439 => x"04001b08",
			3440 => x"00012a04",
			3441 => x"ffbb363d",
			3442 => x"00ea363d",
			3443 => x"05002a04",
			3444 => x"ff37363d",
			3445 => x"006a363d",
			3446 => x"0c001508",
			3447 => x"04002604",
			3448 => x"012f363d",
			3449 => x"0014363d",
			3450 => x"0800180c",
			3451 => x"0f006f04",
			3452 => x"ffa2363d",
			3453 => x"0a003e04",
			3454 => x"00d4363d",
			3455 => x"ffe0363d",
			3456 => x"0a004318",
			3457 => x"04002e10",
			3458 => x"0a003708",
			3459 => x"09001c04",
			3460 => x"004a363d",
			3461 => x"ff0c363d",
			3462 => x"09001f04",
			3463 => x"00df363d",
			3464 => x"ffd8363d",
			3465 => x"0e004d04",
			3466 => x"0082363d",
			3467 => x"fed3363d",
			3468 => x"05004e04",
			3469 => x"00e1363d",
			3470 => x"ffb6363d",
			3471 => x"05002708",
			3472 => x"03002c04",
			3473 => x"ff3e36c1",
			3474 => x"000836c1",
			3475 => x"08001c28",
			3476 => x"02012f20",
			3477 => x"07002b10",
			3478 => x"0e005d04",
			3479 => x"ff9a36c1",
			3480 => x"0a002d04",
			3481 => x"ffee36c1",
			3482 => x"04002e04",
			3483 => x"00d036c1",
			3484 => x"002c36c1",
			3485 => x"0600a108",
			3486 => x"00010a04",
			3487 => x"ff8336c1",
			3488 => x"008236c1",
			3489 => x"0e008504",
			3490 => x"ff6036c1",
			3491 => x"fff036c1",
			3492 => x"00014504",
			3493 => x"00d336c1",
			3494 => x"001036c1",
			3495 => x"0a003704",
			3496 => x"ff3f36c1",
			3497 => x"0c001904",
			3498 => x"005636c1",
			3499 => x"0a004504",
			3500 => x"ffac36c1",
			3501 => x"03004104",
			3502 => x"003f36c1",
			3503 => x"ffe936c1",
			3504 => x"0c001418",
			3505 => x"0600a50c",
			3506 => x"08001504",
			3507 => x"0031376d",
			3508 => x"0d001304",
			3509 => x"fe9a376d",
			3510 => x"0041376d",
			3511 => x"09001908",
			3512 => x"08001b04",
			3513 => x"011f376d",
			3514 => x"ffb8376d",
			3515 => x"ff6c376d",
			3516 => x"0e008a34",
			3517 => x"0100091c",
			3518 => x"0e00740c",
			3519 => x"04004304",
			3520 => x"fee5376d",
			3521 => x"08001b04",
			3522 => x"ffe2376d",
			3523 => x"00dd376d",
			3524 => x"0f00c60c",
			3525 => x"05002704",
			3526 => x"ff64376d",
			3527 => x"02011904",
			3528 => x"0087376d",
			3529 => x"0174376d",
			3530 => x"0017376d",
			3531 => x"05003108",
			3532 => x"0f00c404",
			3533 => x"fe9a376d",
			3534 => x"0046376d",
			3535 => x"0d00160c",
			3536 => x"04003808",
			3537 => x"00009f04",
			3538 => x"ffc0376d",
			3539 => x"0103376d",
			3540 => x"ff7a376d",
			3541 => x"ff4b376d",
			3542 => x"01000904",
			3543 => x"fee7376d",
			3544 => x"09001b04",
			3545 => x"00a7376d",
			3546 => x"ff73376d",
			3547 => x"0c00141c",
			3548 => x"0e008210",
			3549 => x"0400200c",
			3550 => x"08001504",
			3551 => x"000f3829",
			3552 => x"01000a04",
			3553 => x"ff303829",
			3554 => x"00073829",
			3555 => x"00293829",
			3556 => x"00014408",
			3557 => x"08001b04",
			3558 => x"006e3829",
			3559 => x"fff63829",
			3560 => x"ffca3829",
			3561 => x"01000b30",
			3562 => x"00010714",
			3563 => x"03003804",
			3564 => x"ff703829",
			3565 => x"07002b0c",
			3566 => x"09001f04",
			3567 => x"ffe43829",
			3568 => x"0b001804",
			3569 => x"00833829",
			3570 => x"ffeb3829",
			3571 => x"ffb43829",
			3572 => x"0600a50c",
			3573 => x"08001c08",
			3574 => x"07002c04",
			3575 => x"00d23829",
			3576 => x"001b3829",
			3577 => x"ffe43829",
			3578 => x"00013c08",
			3579 => x"00013504",
			3580 => x"005b3829",
			3581 => x"ff3b3829",
			3582 => x"0e008b04",
			3583 => x"00903829",
			3584 => x"ffed3829",
			3585 => x"0a00450c",
			3586 => x"07003104",
			3587 => x"ff683829",
			3588 => x"07003204",
			3589 => x"00223829",
			3590 => x"ffdd3829",
			3591 => x"07003104",
			3592 => x"002e3829",
			3593 => x"fff43829",
			3594 => x"05002c24",
			3595 => x"0201301c",
			3596 => x"0d000e04",
			3597 => x"001238e5",
			3598 => x"0300270c",
			3599 => x"03002308",
			3600 => x"03002104",
			3601 => x"fff538e5",
			3602 => x"000438e5",
			3603 => x"ff7538e5",
			3604 => x"04001a04",
			3605 => x"002238e5",
			3606 => x"0e008104",
			3607 => x"ffc738e5",
			3608 => x"001b38e5",
			3609 => x"0f00d404",
			3610 => x"004438e5",
			3611 => x"ffce38e5",
			3612 => x"05003514",
			3613 => x"0e008a0c",
			3614 => x"09001d08",
			3615 => x"0000e704",
			3616 => x"fffc38e5",
			3617 => x"008438e5",
			3618 => x"fff638e5",
			3619 => x"00013f04",
			3620 => x"ffde38e5",
			3621 => x"000438e5",
			3622 => x"03003b1c",
			3623 => x"0201020c",
			3624 => x"0e004d08",
			3625 => x"06005204",
			3626 => x"fff738e5",
			3627 => x"001438e5",
			3628 => x"ff9938e5",
			3629 => x"08001c04",
			3630 => x"003538e5",
			3631 => x"0a003b04",
			3632 => x"ffd038e5",
			3633 => x"03003404",
			3634 => x"000a38e5",
			3635 => x"fffd38e5",
			3636 => x"05004e08",
			3637 => x"0f006f04",
			3638 => x"fff238e5",
			3639 => x"005338e5",
			3640 => x"ffe238e5",
			3641 => x"0c001a34",
			3642 => x"06006710",
			3643 => x"08001c04",
			3644 => x"fe623951",
			3645 => x"0d001308",
			3646 => x"04001804",
			3647 => x"fed73951",
			3648 => x"030d3951",
			3649 => x"fe783951",
			3650 => x"0e009020",
			3651 => x"0300240c",
			3652 => x"0d001108",
			3653 => x"07002a04",
			3654 => x"fe663951",
			3655 => x"01cb3951",
			3656 => x"fe433951",
			3657 => x"01000d10",
			3658 => x"0a003408",
			3659 => x"00013a04",
			3660 => x"00293951",
			3661 => x"01b13951",
			3662 => x"05004e04",
			3663 => x"01f13951",
			3664 => x"fe923951",
			3665 => x"fe643951",
			3666 => x"fe4f3951",
			3667 => x"fe663951",
			3668 => x"01000b34",
			3669 => x"01000308",
			3670 => x"0d001104",
			3671 => x"fe5a39cd",
			3672 => x"006c39cd",
			3673 => x"05002504",
			3674 => x"fea839cd",
			3675 => x"0b00140c",
			3676 => x"06009704",
			3677 => x"febe39cd",
			3678 => x"08001b04",
			3679 => x"018e39cd",
			3680 => x"007f39cd",
			3681 => x"0e007e10",
			3682 => x"0200fb08",
			3683 => x"0e006604",
			3684 => x"007539cd",
			3685 => x"fe8539cd",
			3686 => x"06009804",
			3687 => x"011b39cd",
			3688 => x"01b639cd",
			3689 => x"0e008204",
			3690 => x"fe9439cd",
			3691 => x"0e008a04",
			3692 => x"00c239cd",
			3693 => x"ff1539cd",
			3694 => x"07003104",
			3695 => x"fe6439cd",
			3696 => x"07003204",
			3697 => x"012439cd",
			3698 => x"feb539cd",
			3699 => x"0300261c",
			3700 => x"0600ae14",
			3701 => x"05002d10",
			3702 => x"0300230c",
			3703 => x"0e007c08",
			3704 => x"03002104",
			3705 => x"ffec3a81",
			3706 => x"002d3a81",
			3707 => x"ffd73a81",
			3708 => x"ff393a81",
			3709 => x"00453a81",
			3710 => x"04001804",
			3711 => x"ffdd3a81",
			3712 => x"00603a81",
			3713 => x"09001c20",
			3714 => x"0c00140c",
			3715 => x"0e008204",
			3716 => x"ff9f3a81",
			3717 => x"08001b04",
			3718 => x"00543a81",
			3719 => x"ffdb3a81",
			3720 => x"01000b10",
			3721 => x"0e007404",
			3722 => x"ffbc3a81",
			3723 => x"0e008704",
			3724 => x"01003a81",
			3725 => x"0600af04",
			3726 => x"ffd23a81",
			3727 => x"00313a81",
			3728 => x"ffaf3a81",
			3729 => x"0a003704",
			3730 => x"ff723a81",
			3731 => x"0b001810",
			3732 => x"04003404",
			3733 => x"00603a81",
			3734 => x"03003b04",
			3735 => x"ff9c3a81",
			3736 => x"05004e04",
			3737 => x"00613a81",
			3738 => x"ffe53a81",
			3739 => x"0a004504",
			3740 => x"ffa53a81",
			3741 => x"05004e04",
			3742 => x"002f3a81",
			3743 => x"ffec3a81",
			3744 => x"0c001414",
			3745 => x"0600a50c",
			3746 => x"08001504",
			3747 => x"00303b25",
			3748 => x"0d001304",
			3749 => x"fea73b25",
			3750 => x"003e3b25",
			3751 => x"01000804",
			3752 => x"011d3b25",
			3753 => x"ff723b25",
			3754 => x"08001608",
			3755 => x"0e007604",
			3756 => x"ff893b25",
			3757 => x"01413b25",
			3758 => x"03002610",
			3759 => x"0e007c08",
			3760 => x"0a002a04",
			3761 => x"ffab3b25",
			3762 => x"00ed3b25",
			3763 => x"00014004",
			3764 => x"fea93b25",
			3765 => x"00563b25",
			3766 => x"09001c10",
			3767 => x"01000b0c",
			3768 => x"08001c08",
			3769 => x"00010a04",
			3770 => x"ff793b25",
			3771 => x"010b3b25",
			3772 => x"ff553b25",
			3773 => x"ff273b25",
			3774 => x"0a00370c",
			3775 => x"00013e04",
			3776 => x"fec63b25",
			3777 => x"00014204",
			3778 => x"001b3b25",
			3779 => x"ff9e3b25",
			3780 => x"0d001204",
			3781 => x"ff393b25",
			3782 => x"09002104",
			3783 => x"00a63b25",
			3784 => x"ff4b3b25",
			3785 => x"0e008a48",
			3786 => x"0d001328",
			3787 => x"0e008220",
			3788 => x"05002c10",
			3789 => x"0a002c0c",
			3790 => x"06009c08",
			3791 => x"09001904",
			3792 => x"ffeb3bd9",
			3793 => x"00113bd9",
			3794 => x"ff8e3bd9",
			3795 => x"00093bd9",
			3796 => x"00012d0c",
			3797 => x"08001b08",
			3798 => x"03003b04",
			3799 => x"ffb33bd9",
			3800 => x"fffd3bd9",
			3801 => x"00393bd9",
			3802 => x"00633bd9",
			3803 => x"01000904",
			3804 => x"00a03bd9",
			3805 => x"00033bd9",
			3806 => x"08001808",
			3807 => x"06006704",
			3808 => x"fff73bd9",
			3809 => x"003b3bd9",
			3810 => x"03002c04",
			3811 => x"ff893bd9",
			3812 => x"05003508",
			3813 => x"00010a04",
			3814 => x"fff13bd9",
			3815 => x"005b3bd9",
			3816 => x"0a004504",
			3817 => x"ffa43bd9",
			3818 => x"03004104",
			3819 => x"00193bd9",
			3820 => x"ffee3bd9",
			3821 => x"0b001308",
			3822 => x"0f00da04",
			3823 => x"00253bd9",
			3824 => x"fffa3bd9",
			3825 => x"01000904",
			3826 => x"ff853bd9",
			3827 => x"01000b04",
			3828 => x"000a3bd9",
			3829 => x"ffeb3bd9",
			3830 => x"0e009030",
			3831 => x"02013028",
			3832 => x"02012c24",
			3833 => x"00012f1c",
			3834 => x"0e008010",
			3835 => x"0a003d08",
			3836 => x"04001904",
			3837 => x"001c3c3d",
			3838 => x"ff813c3d",
			3839 => x"04003804",
			3840 => x"00413c3d",
			3841 => x"ffda3c3d",
			3842 => x"02011f08",
			3843 => x"01000d04",
			3844 => x"00633c3d",
			3845 => x"ffef3c3d",
			3846 => x"ffd63c3d",
			3847 => x"01000904",
			3848 => x"00933c3d",
			3849 => x"ff9a3c3d",
			3850 => x"ff983c3d",
			3851 => x"08001c04",
			3852 => x"00963c3d",
			3853 => x"ffee3c3d",
			3854 => x"ffa33c3d",
			3855 => x"0d001640",
			3856 => x"0300240c",
			3857 => x"0d001108",
			3858 => x"04001804",
			3859 => x"fe833cc1",
			3860 => x"01713cc1",
			3861 => x"fe503cc1",
			3862 => x"0e008a24",
			3863 => x"0f006f0c",
			3864 => x"0e004d08",
			3865 => x"00009904",
			3866 => x"feb53cc1",
			3867 => x"02123cc1",
			3868 => x"fe733cc1",
			3869 => x"0a00370c",
			3870 => x"08001c08",
			3871 => x"00013a04",
			3872 => x"00443cc1",
			3873 => x"01983cc1",
			3874 => x"fe273cc1",
			3875 => x"05004e08",
			3876 => x"0d001204",
			3877 => x"00223cc1",
			3878 => x"02373cc1",
			3879 => x"fea43cc1",
			3880 => x"0b001408",
			3881 => x"00013604",
			3882 => x"fec83cc1",
			3883 => x"01743cc1",
			3884 => x"00014604",
			3885 => x"fde33cc1",
			3886 => x"fffc3cc1",
			3887 => x"fe6e3cc1",
			3888 => x"05002c28",
			3889 => x"03002618",
			3890 => x"02013014",
			3891 => x"03002310",
			3892 => x"0d00110c",
			3893 => x"0d001004",
			3894 => x"ffc33d85",
			3895 => x"04001304",
			3896 => x"ffec3d85",
			3897 => x"009f3d85",
			3898 => x"ff403d85",
			3899 => x"fe8d3d85",
			3900 => x"003c3d85",
			3901 => x"00012a04",
			3902 => x"fed83d85",
			3903 => x"07002c04",
			3904 => x"011e3d85",
			3905 => x"01000904",
			3906 => x"ff043d85",
			3907 => x"00ba3d85",
			3908 => x"0e008a30",
			3909 => x"0e006510",
			3910 => x"0000af0c",
			3911 => x"03003804",
			3912 => x"ff263d85",
			3913 => x"0a003e04",
			3914 => x"01103d85",
			3915 => x"ff7d3d85",
			3916 => x"fef23d85",
			3917 => x"08001c10",
			3918 => x"0d00150c",
			3919 => x"05004e08",
			3920 => x"07002a04",
			3921 => x"00953d85",
			3922 => x"015b3d85",
			3923 => x"ffc23d85",
			3924 => x"ff5e3d85",
			3925 => x"0a003704",
			3926 => x"fed23d85",
			3927 => x"08001f08",
			3928 => x"04004304",
			3929 => x"01443d85",
			3930 => x"fff13d85",
			3931 => x"ff993d85",
			3932 => x"02013804",
			3933 => x"fefd3d85",
			3934 => x"02013a04",
			3935 => x"00133d85",
			3936 => x"ffd63d85",
			3937 => x"03003b3c",
			3938 => x"09001e38",
			3939 => x"0c001414",
			3940 => x"0600a50c",
			3941 => x"04002008",
			3942 => x"08001504",
			3943 => x"002c3e19",
			3944 => x"fe513e19",
			3945 => x"010c3e19",
			3946 => x"01000804",
			3947 => x"011f3e19",
			3948 => x"ff433e19",
			3949 => x"0e008a14",
			3950 => x"00010a04",
			3951 => x"fec73e19",
			3952 => x"03002608",
			3953 => x"0d001204",
			3954 => x"009b3e19",
			3955 => x"fee53e19",
			3956 => x"08001c04",
			3957 => x"01183e19",
			3958 => x"ffba3e19",
			3959 => x"01000904",
			3960 => x"fea43e19",
			3961 => x"0600b608",
			3962 => x"0a002d04",
			3963 => x"00fb3e19",
			3964 => x"fff63e19",
			3965 => x"ff7f3e19",
			3966 => x"fe913e19",
			3967 => x"05004e0c",
			3968 => x"0f006f04",
			3969 => x"ff7d3e19",
			3970 => x"09002504",
			3971 => x"01923e19",
			3972 => x"fff23e19",
			3973 => x"ff233e19",
			3974 => x"00012f40",
			3975 => x"05003018",
			3976 => x"0c00170c",
			3977 => x"0e008304",
			3978 => x"fee73ef5",
			3979 => x"03002c04",
			3980 => x"ff923ef5",
			3981 => x"00623ef5",
			3982 => x"07002a08",
			3983 => x"07002904",
			3984 => x"fff63ef5",
			3985 => x"006b3ef5",
			3986 => x"ffcd3ef5",
			3987 => x"0500350c",
			3988 => x"0a002f04",
			3989 => x"ffe73ef5",
			3990 => x"01000d04",
			3991 => x"00df3ef5",
			3992 => x"fff73ef5",
			3993 => x"0a004314",
			3994 => x"0e004d08",
			3995 => x"0f005804",
			3996 => x"ffe03ef5",
			3997 => x"00683ef5",
			3998 => x"08001804",
			3999 => x"00233ef5",
			4000 => x"00011404",
			4001 => x"fefe3ef5",
			4002 => x"fff13ef5",
			4003 => x"05004e04",
			4004 => x"009f3ef5",
			4005 => x"ffc53ef5",
			4006 => x"0e007f04",
			4007 => x"00fa3ef5",
			4008 => x"03002910",
			4009 => x"0600ad08",
			4010 => x"02013004",
			4011 => x"fefc3ef5",
			4012 => x"00513ef5",
			4013 => x"0600b604",
			4014 => x"00903ef5",
			4015 => x"ff6b3ef5",
			4016 => x"08001b08",
			4017 => x"08001804",
			4018 => x"001d3ef5",
			4019 => x"00f13ef5",
			4020 => x"0500390c",
			4021 => x"02013804",
			4022 => x"ff643ef5",
			4023 => x"00014c04",
			4024 => x"00163ef5",
			4025 => x"fff43ef5",
			4026 => x"0c001b04",
			4027 => x"00373ef5",
			4028 => x"fff63ef5",
			4029 => x"07002b30",
			4030 => x"03002710",
			4031 => x"04001d04",
			4032 => x"fefe3fc1",
			4033 => x"01000704",
			4034 => x"00b63fc1",
			4035 => x"04001e04",
			4036 => x"000c3fc1",
			4037 => x"ffba3fc1",
			4038 => x"01000b1c",
			4039 => x"07002910",
			4040 => x"07002608",
			4041 => x"00009f04",
			4042 => x"ffbe3fc1",
			4043 => x"00ce3fc1",
			4044 => x"04002e04",
			4045 => x"fff83fc1",
			4046 => x"ff4b3fc1",
			4047 => x"06006704",
			4048 => x"ffc73fc1",
			4049 => x"00010704",
			4050 => x"00603fc1",
			4051 => x"01203fc1",
			4052 => x"ff5a3fc1",
			4053 => x"02012f2c",
			4054 => x"09001908",
			4055 => x"0f00b604",
			4056 => x"00253fc1",
			4057 => x"fecb3fc1",
			4058 => x"08001808",
			4059 => x"00012504",
			4060 => x"ffaf3fc1",
			4061 => x"008e3fc1",
			4062 => x"0a002d0c",
			4063 => x"0e007908",
			4064 => x"07002c04",
			4065 => x"005e3fc1",
			4066 => x"fff53fc1",
			4067 => x"fecd3fc1",
			4068 => x"09001d08",
			4069 => x"00011e04",
			4070 => x"ffcc3fc1",
			4071 => x"00cc3fc1",
			4072 => x"0a004504",
			4073 => x"ff243fc1",
			4074 => x"005a3fc1",
			4075 => x"0e009008",
			4076 => x"08001c04",
			4077 => x"00f63fc1",
			4078 => x"ff9e3fc1",
			4079 => x"ff6a3fc1",
			4080 => x"05004c48",
			4081 => x"01000514",
			4082 => x"0c001404",
			4083 => x"fec8405d",
			4084 => x"09001b08",
			4085 => x"03002304",
			4086 => x"ff70405d",
			4087 => x"0116405d",
			4088 => x"0d001304",
			4089 => x"fef6405d",
			4090 => x"000f405d",
			4091 => x"0d001524",
			4092 => x"01000b20",
			4093 => x"0a002c10",
			4094 => x"0c001408",
			4095 => x"0c001304",
			4096 => x"fff9405d",
			4097 => x"feaf405d",
			4098 => x"00012a04",
			4099 => x"ff0b405d",
			4100 => x"0096405d",
			4101 => x"0c001508",
			4102 => x"05002704",
			4103 => x"ffc4405d",
			4104 => x"0159405d",
			4105 => x"0e008a04",
			4106 => x"0058405d",
			4107 => x"ff00405d",
			4108 => x"febb405d",
			4109 => x"0e008708",
			4110 => x"0b001504",
			4111 => x"ffc7405d",
			4112 => x"fead405d",
			4113 => x"0f00b704",
			4114 => x"00e6405d",
			4115 => x"ff55405d",
			4116 => x"05004e04",
			4117 => x"015d405d",
			4118 => x"ff33405d",
			4119 => x"01000b4c",
			4120 => x"0d001544",
			4121 => x"01000518",
			4122 => x"08001b10",
			4123 => x"0d00130c",
			4124 => x"0f00bc08",
			4125 => x"0a003704",
			4126 => x"ff6d4119",
			4127 => x"00044119",
			4128 => x"fff54119",
			4129 => x"00084119",
			4130 => x"07002904",
			4131 => x"fffc4119",
			4132 => x"004d4119",
			4133 => x"08001914",
			4134 => x"05002708",
			4135 => x"07002e04",
			4136 => x"ffa84119",
			4137 => x"00344119",
			4138 => x"04003608",
			4139 => x"0e005d04",
			4140 => x"fff34119",
			4141 => x"00d94119",
			4142 => x"ffd64119",
			4143 => x"0500310c",
			4144 => x"00013d08",
			4145 => x"0600ab04",
			4146 => x"ff594119",
			4147 => x"00164119",
			4148 => x"00334119",
			4149 => x"04003408",
			4150 => x"08001c04",
			4151 => x"006f4119",
			4152 => x"00024119",
			4153 => x"ffcd4119",
			4154 => x"0c001704",
			4155 => x"00084119",
			4156 => x"ff904119",
			4157 => x"0400370c",
			4158 => x"07003104",
			4159 => x"ff7c4119",
			4160 => x"07003204",
			4161 => x"001f4119",
			4162 => x"ffe14119",
			4163 => x"05004f04",
			4164 => x"00294119",
			4165 => x"fff44119",
			4166 => x"01000d30",
			4167 => x"05002504",
			4168 => x"fe93417d",
			4169 => x"08001504",
			4170 => x"0151417d",
			4171 => x"0a003714",
			4172 => x"08001c10",
			4173 => x"02012f08",
			4174 => x"0f00c704",
			4175 => x"0021417d",
			4176 => x"fe2a417d",
			4177 => x"0600ae04",
			4178 => x"0182417d",
			4179 => x"005a417d",
			4180 => x"fe67417d",
			4181 => x"0201020c",
			4182 => x"0f007c08",
			4183 => x"09001f04",
			4184 => x"fec0417d",
			4185 => x"0104417d",
			4186 => x"fe73417d",
			4187 => x"0600a204",
			4188 => x"01e0417d",
			4189 => x"0079417d",
			4190 => x"fe7c417d",
			4191 => x"0e008a4c",
			4192 => x"0600ab48",
			4193 => x"05002b18",
			4194 => x"03002710",
			4195 => x"0d00110c",
			4196 => x"0d000f04",
			4197 => x"ff854239",
			4198 => x"0e006f04",
			4199 => x"fffa4239",
			4200 => x"004f4239",
			4201 => x"ff064239",
			4202 => x"08001b04",
			4203 => x"008e4239",
			4204 => x"ff824239",
			4205 => x"01000a18",
			4206 => x"0f00bc10",
			4207 => x"0d001208",
			4208 => x"0d001104",
			4209 => x"00224239",
			4210 => x"ff2e4239",
			4211 => x"0d001504",
			4212 => x"009a4239",
			4213 => x"ffb54239",
			4214 => x"01000704",
			4215 => x"00f94239",
			4216 => x"00274239",
			4217 => x"0300330c",
			4218 => x"05002e04",
			4219 => x"000f4239",
			4220 => x"05003904",
			4221 => x"ff654239",
			4222 => x"ffff4239",
			4223 => x"0e006704",
			4224 => x"ff8b4239",
			4225 => x"0d001604",
			4226 => x"00ab4239",
			4227 => x"ffd34239",
			4228 => x"00b34239",
			4229 => x"0b001308",
			4230 => x"0f00df04",
			4231 => x"005b4239",
			4232 => x"fff04239",
			4233 => x"01000904",
			4234 => x"ff1e4239",
			4235 => x"01000b04",
			4236 => x"00224239",
			4237 => x"ffcb4239",
			4238 => x"0100051c",
			4239 => x"0c001404",
			4240 => x"fe774337",
			4241 => x"09001b08",
			4242 => x"05002b04",
			4243 => x"ff214337",
			4244 => x"016f4337",
			4245 => x"0d001308",
			4246 => x"08001804",
			4247 => x"ffd84337",
			4248 => x"fe774337",
			4249 => x"04002e04",
			4250 => x"008c4337",
			4251 => x"ff3c4337",
			4252 => x"08001928",
			4253 => x"01000b24",
			4254 => x"04001d10",
			4255 => x"04001a0c",
			4256 => x"04001808",
			4257 => x"0d001304",
			4258 => x"ff224337",
			4259 => x"001a4337",
			4260 => x"018f4337",
			4261 => x"ff374337",
			4262 => x"04003610",
			4263 => x"02012d08",
			4264 => x"00011204",
			4265 => x"008e4337",
			4266 => x"01aa4337",
			4267 => x"0600a904",
			4268 => x"01224337",
			4269 => x"ff894337",
			4270 => x"ff034337",
			4271 => x"fea84337",
			4272 => x"03002c10",
			4273 => x"00014208",
			4274 => x"0a003204",
			4275 => x"fe614337",
			4276 => x"00774337",
			4277 => x"00014704",
			4278 => x"013b4337",
			4279 => x"fefd4337",
			4280 => x"05003510",
			4281 => x"0a002f04",
			4282 => x"ff714337",
			4283 => x"09001d08",
			4284 => x"0600bd04",
			4285 => x"01974337",
			4286 => x"ffc94337",
			4287 => x"ff4d4337",
			4288 => x"0a003d0c",
			4289 => x"04002304",
			4290 => x"00284337",
			4291 => x"07002d04",
			4292 => x"feac4337",
			4293 => x"ff854337",
			4294 => x"05004908",
			4295 => x"05004504",
			4296 => x"ff934337",
			4297 => x"01634337",
			4298 => x"0a004504",
			4299 => x"fe924337",
			4300 => x"01074337",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1489, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2851, initial_addr_3'length));
	end generate gen_rom_2;

	gen_rom_3: if SELECT_ROM = 3 generate
		bank <= (
			0 => x"0d001a20",
			1 => x"09001404",
			2 => x"018c0055",
			3 => x"0a002308",
			4 => x"08001504",
			5 => x"ffd60055",
			6 => x"fe8c0055",
			7 => x"0a002404",
			8 => x"01480055",
			9 => x"0400330c",
			10 => x"04002e08",
			11 => x"0b001804",
			12 => x"fff00055",
			13 => x"009c0055",
			14 => x"01550055",
			15 => x"fe980055",
			16 => x"01000d08",
			17 => x"0000e704",
			18 => x"ffa90055",
			19 => x"01010055",
			20 => x"fe720055",
			21 => x"0f008b14",
			22 => x"04000808",
			23 => x"06003504",
			24 => x"fe8b00b9",
			25 => x"08b200b9",
			26 => x"0c001708",
			27 => x"0b001604",
			28 => x"fe6900b9",
			29 => x"018a00b9",
			30 => x"fe6700b9",
			31 => x"0900231c",
			32 => x"03003518",
			33 => x"0e006f04",
			34 => x"01ed00b9",
			35 => x"03002108",
			36 => x"00012204",
			37 => x"fe5500b9",
			38 => x"ff7000b9",
			39 => x"0200eb04",
			40 => x"fe7100b9",
			41 => x"0e009704",
			42 => x"00d700b9",
			43 => x"fe7f00b9",
			44 => x"ff2b00b9",
			45 => x"fe6b00b9",
			46 => x"0200fa18",
			47 => x"0f008b10",
			48 => x"09001504",
			49 => x"0004012d",
			50 => x"0c001708",
			51 => x"0b001704",
			52 => x"fe61012d",
			53 => x"0132012d",
			54 => x"fe5f012d",
			55 => x"07002b04",
			56 => x"01e5012d",
			57 => x"fe62012d",
			58 => x"09002320",
			59 => x"0e00971c",
			60 => x"0c001914",
			61 => x"0d001810",
			62 => x"07002c08",
			63 => x"05002c04",
			64 => x"01c1012d",
			65 => x"fe98012d",
			66 => x"01000704",
			67 => x"03e6012d",
			68 => x"01d6012d",
			69 => x"ff68012d",
			70 => x"0a003404",
			71 => x"0155012d",
			72 => x"0345012d",
			73 => x"fe6c012d",
			74 => x"fe61012d",
			75 => x"0400262c",
			76 => x"04002528",
			77 => x"08002218",
			78 => x"0a003614",
			79 => x"05003210",
			80 => x"0c001808",
			81 => x"04001604",
			82 => x"008201b9",
			83 => x"ffd101b9",
			84 => x"04001a04",
			85 => x"fef801b9",
			86 => x"00d601b9",
			87 => x"ff0301b9",
			88 => x"011a01b9",
			89 => x"04001b0c",
			90 => x"07003104",
			91 => x"ff9001b9",
			92 => x"07003304",
			93 => x"008b01b9",
			94 => x"ffed01b9",
			95 => x"feba01b9",
			96 => x"013d01b9",
			97 => x"04002e0c",
			98 => x"0b001804",
			99 => x"fec601b9",
			100 => x"0b001a04",
			101 => x"00d001b9",
			102 => x"feed01b9",
			103 => x"0400320c",
			104 => x"0f009c04",
			105 => x"ff7501b9",
			106 => x"03003504",
			107 => x"012201b9",
			108 => x"fff301b9",
			109 => x"ff0701b9",
			110 => x"0001111c",
			111 => x"0d001710",
			112 => x"09001f04",
			113 => x"ff81025d",
			114 => x"03002d04",
			115 => x"ffe9025d",
			116 => x"05004504",
			117 => x"003a025d",
			118 => x"ffef025d",
			119 => x"05002808",
			120 => x"09001e04",
			121 => x"0048025d",
			122 => x"fffa025d",
			123 => x"ffc9025d",
			124 => x"06009b08",
			125 => x"01000b04",
			126 => x"008b025d",
			127 => x"0004025d",
			128 => x"02011d0c",
			129 => x"02010f04",
			130 => x"001c025d",
			131 => x"0c001404",
			132 => x"0002025d",
			133 => x"ff6c025d",
			134 => x"0600a810",
			135 => x"00013a0c",
			136 => x"07002b04",
			137 => x"ffce025d",
			138 => x"05003804",
			139 => x"00a8025d",
			140 => x"fff9025d",
			141 => x"ffba025d",
			142 => x"01000704",
			143 => x"004d025d",
			144 => x"00014508",
			145 => x"05003404",
			146 => x"ff65025d",
			147 => x"fff6025d",
			148 => x"07003204",
			149 => x"0045025d",
			150 => x"ffc0025d",
			151 => x"04000808",
			152 => x"0e003304",
			153 => x"ff2202b9",
			154 => x"061f02b9",
			155 => x"0e004d04",
			156 => x"fe8902b9",
			157 => x"00008f04",
			158 => x"020202b9",
			159 => x"0f008b04",
			160 => x"fe8502b9",
			161 => x"0f00c010",
			162 => x"0d001308",
			163 => x"01000904",
			164 => x"005502b9",
			165 => x"019a02b9",
			166 => x"0c001604",
			167 => x"fe8602b9",
			168 => x"004a02b9",
			169 => x"00013104",
			170 => x"fe3e02b9",
			171 => x"0d001804",
			172 => x"004202b9",
			173 => x"ff3f02b9",
			174 => x"04002630",
			175 => x"0400252c",
			176 => x"04002324",
			177 => x"01000410",
			178 => x"07002b0c",
			179 => x"0d001108",
			180 => x"09001704",
			181 => x"00920355",
			182 => x"00040355",
			183 => x"ff320355",
			184 => x"00e80355",
			185 => x"0a003610",
			186 => x"0a003208",
			187 => x"00014504",
			188 => x"ffec0355",
			189 => x"00710355",
			190 => x"0d001704",
			191 => x"fefd0355",
			192 => x"fff10355",
			193 => x"00b60355",
			194 => x"09001f04",
			195 => x"001e0355",
			196 => x"feff0355",
			197 => x"01010355",
			198 => x"04002b0c",
			199 => x"05003904",
			200 => x"ff230355",
			201 => x"05003a04",
			202 => x"005f0355",
			203 => x"ff7e0355",
			204 => x"04003210",
			205 => x"0c001804",
			206 => x"ffb10355",
			207 => x"0200ef04",
			208 => x"ffdc0355",
			209 => x"07003a04",
			210 => x"00990355",
			211 => x"fff10355",
			212 => x"ff760355",
			213 => x"00010a1c",
			214 => x"0f008b10",
			215 => x"09001504",
			216 => x"cf4203f9",
			217 => x"0c001708",
			218 => x"0c001604",
			219 => x"cdde03f9",
			220 => x"ce4603f9",
			221 => x"cddc03f9",
			222 => x"07002b04",
			223 => x"d5cf03f9",
			224 => x"0200fa04",
			225 => x"cddf03f9",
			226 => x"cfe103f9",
			227 => x"09002230",
			228 => x"0e00962c",
			229 => x"09001d1c",
			230 => x"0a002f0c",
			231 => x"0e007704",
			232 => x"e86903f9",
			233 => x"03002104",
			234 => x"cded03f9",
			235 => x"dab003f9",
			236 => x"05003008",
			237 => x"0f00c204",
			238 => x"d82303f9",
			239 => x"cfe103f9",
			240 => x"00014204",
			241 => x"cde703f9",
			242 => x"cfff03f9",
			243 => x"07003208",
			244 => x"0f00ba04",
			245 => x"dc3403f9",
			246 => x"e8ff03f9",
			247 => x"0a003604",
			248 => x"d57703f9",
			249 => x"e12d03f9",
			250 => x"cde203f9",
			251 => x"0d001904",
			252 => x"d20803f9",
			253 => x"cddc03f9",
			254 => x"0f008b0c",
			255 => x"0c001708",
			256 => x"0b001704",
			257 => x"fe640485",
			258 => x"017b0485",
			259 => x"fe640485",
			260 => x"09002338",
			261 => x"0600ae20",
			262 => x"0f00c614",
			263 => x"0600a810",
			264 => x"01000908",
			265 => x"09001904",
			266 => x"01400485",
			267 => x"fea30485",
			268 => x"00012a04",
			269 => x"00b90485",
			270 => x"021b0485",
			271 => x"fdfe0485",
			272 => x"0c001504",
			273 => x"fe5d0485",
			274 => x"00013c04",
			275 => x"034c0485",
			276 => x"016f0485",
			277 => x"0b00150c",
			278 => x"0600b704",
			279 => x"fe0b0485",
			280 => x"0d001204",
			281 => x"01d60485",
			282 => x"fe500485",
			283 => x"07003404",
			284 => x"01560485",
			285 => x"05003304",
			286 => x"fe340485",
			287 => x"00a90485",
			288 => x"fe670485",
			289 => x"0600a948",
			290 => x"0e008130",
			291 => x"0e00802c",
			292 => x"0001191c",
			293 => x"0c00150c",
			294 => x"03001004",
			295 => x"00290551",
			296 => x"04002004",
			297 => x"ff480551",
			298 => x"00060551",
			299 => x"01000b08",
			300 => x"0200d104",
			301 => x"ffcb0551",
			302 => x"008c0551",
			303 => x"05002504",
			304 => x"00350551",
			305 => x"ff5f0551",
			306 => x"05002a08",
			307 => x"0600a004",
			308 => x"00bc0551",
			309 => x"fffd0551",
			310 => x"01000904",
			311 => x"ff940551",
			312 => x"00280551",
			313 => x"ff660551",
			314 => x"02011d0c",
			315 => x"00011808",
			316 => x"00010c04",
			317 => x"ffe70551",
			318 => x"00500551",
			319 => x"ff880551",
			320 => x"02012804",
			321 => x"00b10551",
			322 => x"0b001704",
			323 => x"ffad0551",
			324 => x"00580551",
			325 => x"00014514",
			326 => x"01000704",
			327 => x"fffe0551",
			328 => x"0b001b08",
			329 => x"04002604",
			330 => x"ff270551",
			331 => x"fff50551",
			332 => x"04002304",
			333 => x"00310551",
			334 => x"ffdd0551",
			335 => x"0e009408",
			336 => x"09001b04",
			337 => x"ffbb0551",
			338 => x"006d0551",
			339 => x"ff8e0551",
			340 => x"0d001854",
			341 => x"0c001628",
			342 => x"09001918",
			343 => x"00013c14",
			344 => x"0b001208",
			345 => x"04001504",
			346 => x"ffb2062d",
			347 => x"0012062d",
			348 => x"04002008",
			349 => x"09001804",
			350 => x"000c062d",
			351 => x"00ab062d",
			352 => x"ffda062d",
			353 => x"ff81062d",
			354 => x"0e009008",
			355 => x"0b001504",
			356 => x"ff5a062d",
			357 => x"0004062d",
			358 => x"0e009604",
			359 => x"007c062d",
			360 => x"ffe8062d",
			361 => x"01000814",
			362 => x"04001c08",
			363 => x"07002b04",
			364 => x"ffdd062d",
			365 => x"009b062d",
			366 => x"05002b04",
			367 => x"0007062d",
			368 => x"01000404",
			369 => x"ffff062d",
			370 => x"ff39062d",
			371 => x"0f00d014",
			372 => x"02012a10",
			373 => x"06009e08",
			374 => x"0a003604",
			375 => x"0082062d",
			376 => x"ffc1062d",
			377 => x"0b001704",
			378 => x"ff92062d",
			379 => x"002c062d",
			380 => x"00cb062d",
			381 => x"ffe2062d",
			382 => x"0900210c",
			383 => x"0c001908",
			384 => x"0c001804",
			385 => x"ff88062d",
			386 => x"fffc062d",
			387 => x"006f062d",
			388 => x"0400230c",
			389 => x"08002308",
			390 => x"08002004",
			391 => x"fffc062d",
			392 => x"0044062d",
			393 => x"ffd1062d",
			394 => x"ff42062d",
			395 => x"09001404",
			396 => x"01bc06a1",
			397 => x"0d001a2c",
			398 => x"0a002308",
			399 => x"08001504",
			400 => x"ffd306a1",
			401 => x"fe8706a1",
			402 => x"0a002404",
			403 => x"016406a1",
			404 => x"04001a10",
			405 => x"04001608",
			406 => x"01000c04",
			407 => x"00f006a1",
			408 => x"fe8f06a1",
			409 => x"09001904",
			410 => x"000b06a1",
			411 => x"fe4606a1",
			412 => x"03002708",
			413 => x"01000e04",
			414 => x"000406a1",
			415 => x"fe2b06a1",
			416 => x"02011d04",
			417 => x"ffb906a1",
			418 => x"009906a1",
			419 => x"01000d08",
			420 => x"0000e704",
			421 => x"ffa306a1",
			422 => x"011306a1",
			423 => x"fe6b06a1",
			424 => x"04002634",
			425 => x"04002530",
			426 => x"0800232c",
			427 => x"0600ae1c",
			428 => x"01000d10",
			429 => x"0c001708",
			430 => x"05002c04",
			431 => x"00c6074d",
			432 => x"fff7074d",
			433 => x"01000a04",
			434 => x"ff00074d",
			435 => x"0109074d",
			436 => x"0600a408",
			437 => x"07001f04",
			438 => x"004c074d",
			439 => x"fe81074d",
			440 => x"00ee074d",
			441 => x"00013604",
			442 => x"fe49074d",
			443 => x"09001d08",
			444 => x"0f00de04",
			445 => x"ff55074d",
			446 => x"00ba074d",
			447 => x"0072074d",
			448 => x"fe90074d",
			449 => x"019a074d",
			450 => x"04002b10",
			451 => x"00014108",
			452 => x"03003404",
			453 => x"fe85074d",
			454 => x"ff78074d",
			455 => x"0600b804",
			456 => x"0096074d",
			457 => x"fea0074d",
			458 => x"0f009c04",
			459 => x"feb9074d",
			460 => x"01000a04",
			461 => x"0127074d",
			462 => x"00012e04",
			463 => x"fe96074d",
			464 => x"00013204",
			465 => x"0171074d",
			466 => x"ff46074d",
			467 => x"04002350",
			468 => x"00010c20",
			469 => x"08001b10",
			470 => x"08001804",
			471 => x"ffa20831",
			472 => x"0f004b04",
			473 => x"ffeb0831",
			474 => x"07002b04",
			475 => x"00780831",
			476 => x"ffed0831",
			477 => x"0d001204",
			478 => x"00160831",
			479 => x"0e007c04",
			480 => x"ff690831",
			481 => x"0e009004",
			482 => x"00080831",
			483 => x"fff80831",
			484 => x"0f00c010",
			485 => x"07002a08",
			486 => x"0e007704",
			487 => x"005f0831",
			488 => x"ff870831",
			489 => x"05003304",
			490 => x"00960831",
			491 => x"fffc0831",
			492 => x"07002c0c",
			493 => x"03002608",
			494 => x"00013d04",
			495 => x"003c0831",
			496 => x"ffd10831",
			497 => x"ff500831",
			498 => x"07002e04",
			499 => x"00820831",
			500 => x"05002c08",
			501 => x"01000904",
			502 => x"00260831",
			503 => x"ff570831",
			504 => x"03002e04",
			505 => x"007a0831",
			506 => x"ffc50831",
			507 => x"04002508",
			508 => x"07003204",
			509 => x"00030831",
			510 => x"ff4b0831",
			511 => x"04002604",
			512 => x"006a0831",
			513 => x"04002b08",
			514 => x"03003404",
			515 => x"ff7e0831",
			516 => x"00050831",
			517 => x"0400320c",
			518 => x"0c001804",
			519 => x"ffda0831",
			520 => x"0200ef04",
			521 => x"ffec0831",
			522 => x"005e0831",
			523 => x"ffbe0831",
			524 => x"0600a844",
			525 => x"02011f34",
			526 => x"05002618",
			527 => x"03002108",
			528 => x"09001504",
			529 => x"003508fd",
			530 => x"ffa508fd",
			531 => x"01000e0c",
			532 => x"0000cc04",
			533 => x"fff008fd",
			534 => x"07002e04",
			535 => x"007708fd",
			536 => x"fffa08fd",
			537 => x"ffed08fd",
			538 => x"01000b14",
			539 => x"01000908",
			540 => x"0c001404",
			541 => x"001808fd",
			542 => x"ff9908fd",
			543 => x"0a003d08",
			544 => x"04002004",
			545 => x"fff608fd",
			546 => x"004f08fd",
			547 => x"ffec08fd",
			548 => x"0e008a04",
			549 => x"ff7608fd",
			550 => x"001108fd",
			551 => x"0e007d04",
			552 => x"ffa908fd",
			553 => x"00013b08",
			554 => x"0a003804",
			555 => x"009c08fd",
			556 => x"fff608fd",
			557 => x"ffd908fd",
			558 => x"01000704",
			559 => x"001908fd",
			560 => x"0c001808",
			561 => x"00014e04",
			562 => x"ff5b08fd",
			563 => x"000508fd",
			564 => x"09002004",
			565 => x"002e08fd",
			566 => x"0e00960c",
			567 => x"0b001b04",
			568 => x"ffa808fd",
			569 => x"0b001d04",
			570 => x"001708fd",
			571 => x"ffef08fd",
			572 => x"0e009804",
			573 => x"002308fd",
			574 => x"fff008fd",
			575 => x"0600a850",
			576 => x"0e008138",
			577 => x"09001914",
			578 => x"0001110c",
			579 => x"08001804",
			580 => x"ff0109e9",
			581 => x"0b001204",
			582 => x"ff9b09e9",
			583 => x"00bf09e9",
			584 => x"06009d04",
			585 => x"013409e9",
			586 => x"002609e9",
			587 => x"0c001610",
			588 => x"0b00150c",
			589 => x"0e007508",
			590 => x"04001c04",
			591 => x"004409e9",
			592 => x"ff8609e9",
			593 => x"feb309e9",
			594 => x"002609e9",
			595 => x"0e008010",
			596 => x"0a002f08",
			597 => x"04001a04",
			598 => x"ff5909e9",
			599 => x"00f009e9",
			600 => x"01000a04",
			601 => x"005709e9",
			602 => x"ff0f09e9",
			603 => x"ff4709e9",
			604 => x"02011d0c",
			605 => x"00011808",
			606 => x"02010104",
			607 => x"ffb909e9",
			608 => x"00b309e9",
			609 => x"ff0c09e9",
			610 => x"02012804",
			611 => x"014209e9",
			612 => x"01000a04",
			613 => x"fef209e9",
			614 => x"00ad09e9",
			615 => x"02012804",
			616 => x"fed909e9",
			617 => x"08002214",
			618 => x"09001b08",
			619 => x"01000804",
			620 => x"004b09e9",
			621 => x"fec409e9",
			622 => x"04002308",
			623 => x"0600b104",
			624 => x"00f009e9",
			625 => x"002009e9",
			626 => x"ffc109e9",
			627 => x"04002808",
			628 => x"03002904",
			629 => x"fffa09e9",
			630 => x"fee809e9",
			631 => x"04002904",
			632 => x"005d09e9",
			633 => x"ffea09e9",
			634 => x"0d001858",
			635 => x"0c00162c",
			636 => x"04002024",
			637 => x"0600a818",
			638 => x"00011910",
			639 => x"0c001508",
			640 => x"05001204",
			641 => x"00200aed",
			642 => x"ff760aed",
			643 => x"0e007104",
			644 => x"ffe80aed",
			645 => x"00450aed",
			646 => x"09001904",
			647 => x"00880aed",
			648 => x"00060aed",
			649 => x"04001908",
			650 => x"04001504",
			651 => x"ffc60aed",
			652 => x"00610aed",
			653 => x"ff740aed",
			654 => x"0b001504",
			655 => x"ff4b0aed",
			656 => x"ffff0aed",
			657 => x"0a003114",
			658 => x"03002104",
			659 => x"ffd10aed",
			660 => x"01000d0c",
			661 => x"07002604",
			662 => x"ffe40aed",
			663 => x"03002904",
			664 => x"00a70aed",
			665 => x"00190aed",
			666 => x"fff10aed",
			667 => x"08001d0c",
			668 => x"0d001504",
			669 => x"ff630aed",
			670 => x"0b001804",
			671 => x"00160aed",
			672 => x"fff10aed",
			673 => x"05003604",
			674 => x"ffcb0aed",
			675 => x"04003104",
			676 => x"00810aed",
			677 => x"ffeb0aed",
			678 => x"05003414",
			679 => x"00014c10",
			680 => x"0b001a08",
			681 => x"08002004",
			682 => x"ffec0aed",
			683 => x"ff590aed",
			684 => x"0b001b04",
			685 => x"00130aed",
			686 => x"fff10aed",
			687 => x"00210aed",
			688 => x"0500370c",
			689 => x"00012e04",
			690 => x"ffd50aed",
			691 => x"02013504",
			692 => x"007f0aed",
			693 => x"fff60aed",
			694 => x"00011808",
			695 => x"00011004",
			696 => x"fff20aed",
			697 => x"001a0aed",
			698 => x"ff8d0aed",
			699 => x"00010e24",
			700 => x"09001c18",
			701 => x"08001804",
			702 => x"ff1d0bd1",
			703 => x"08001b0c",
			704 => x"06004404",
			705 => x"ffd60bd1",
			706 => x"0e006a04",
			707 => x"00e20bd1",
			708 => x"00100bd1",
			709 => x"06009204",
			710 => x"ff610bd1",
			711 => x"006c0bd1",
			712 => x"0d001208",
			713 => x"04001e04",
			714 => x"00620bd1",
			715 => x"ffec0bd1",
			716 => x"fed60bd1",
			717 => x"0600a830",
			718 => x"01000a18",
			719 => x"09001908",
			720 => x"04001f04",
			721 => x"00c90bd1",
			722 => x"ffd20bd1",
			723 => x"03002404",
			724 => x"feff0bd1",
			725 => x"0600a308",
			726 => x"0f00b504",
			727 => x"00880bd1",
			728 => x"ff1d0bd1",
			729 => x"00880bd1",
			730 => x"00012d10",
			731 => x"0a002f04",
			732 => x"00a90bd1",
			733 => x"0b001804",
			734 => x"ff070bd1",
			735 => x"00012104",
			736 => x"00910bd1",
			737 => x"ffd40bd1",
			738 => x"05003804",
			739 => x"01030bd1",
			740 => x"002e0bd1",
			741 => x"02012804",
			742 => x"feed0bd1",
			743 => x"07002c04",
			744 => x"ff300bd1",
			745 => x"0400230c",
			746 => x"03002e08",
			747 => x"09001d04",
			748 => x"00210bd1",
			749 => x"01180bd1",
			750 => x"ff850bd1",
			751 => x"09002204",
			752 => x"ff4e0bd1",
			753 => x"03003304",
			754 => x"ffc30bd1",
			755 => x"00520bd1",
			756 => x"0600a95c",
			757 => x"0e008140",
			758 => x"05002614",
			759 => x"03002108",
			760 => x"09001504",
			761 => x"003f0cc5",
			762 => x"ff800cc5",
			763 => x"01000e08",
			764 => x"0000cc04",
			765 => x"ffe80cc5",
			766 => x"00a20cc5",
			767 => x"ffde0cc5",
			768 => x"04002110",
			769 => x"09001904",
			770 => x"fffe0cc5",
			771 => x"07002f08",
			772 => x"06008504",
			773 => x"00220cc5",
			774 => x"ff100cc5",
			775 => x"00340cc5",
			776 => x"0a00360c",
			777 => x"0d001608",
			778 => x"0d001204",
			779 => x"ffd20cc5",
			780 => x"00ad0cc5",
			781 => x"ffc30cc5",
			782 => x"0d001808",
			783 => x"08001d04",
			784 => x"ffa20cc5",
			785 => x"000b0cc5",
			786 => x"08001d04",
			787 => x"00250cc5",
			788 => x"ffe20cc5",
			789 => x"02011d0c",
			790 => x"00011808",
			791 => x"00010c04",
			792 => x"ffe80cc5",
			793 => x"004d0cc5",
			794 => x"ff8c0cc5",
			795 => x"00013c0c",
			796 => x"0a003808",
			797 => x"02012904",
			798 => x"00ad0cc5",
			799 => x"00290cc5",
			800 => x"ffe90cc5",
			801 => x"ffbd0cc5",
			802 => x"00014514",
			803 => x"01000704",
			804 => x"ffff0cc5",
			805 => x"0b001b08",
			806 => x"04002604",
			807 => x"ff330cc5",
			808 => x"fff50cc5",
			809 => x"04002304",
			810 => x"002f0cc5",
			811 => x"ffdf0cc5",
			812 => x"07003408",
			813 => x"09001b04",
			814 => x"ffb30cc5",
			815 => x"00730cc5",
			816 => x"ff900cc5",
			817 => x"02011c38",
			818 => x"01000d28",
			819 => x"0a003118",
			820 => x"06009f14",
			821 => x"00010a0c",
			822 => x"07002908",
			823 => x"08001804",
			824 => x"ff040db1",
			825 => x"009f0db1",
			826 => x"fee40db1",
			827 => x"0a002804",
			828 => x"002f0db1",
			829 => x"01270db1",
			830 => x"ff1a0db1",
			831 => x"09001f04",
			832 => x"febd0db1",
			833 => x"08001f04",
			834 => x"ff740db1",
			835 => x"0200de04",
			836 => x"fff50db1",
			837 => x"00ea0db1",
			838 => x"01001f0c",
			839 => x"0a003d04",
			840 => x"feac0db1",
			841 => x"06009604",
			842 => x"ffec0db1",
			843 => x"005c0db1",
			844 => x"00540db1",
			845 => x"07003734",
			846 => x"00013a1c",
			847 => x"0b001510",
			848 => x"0d00130c",
			849 => x"00012f04",
			850 => x"00b20db1",
			851 => x"0f00c204",
			852 => x"ff5c0db1",
			853 => x"00520db1",
			854 => x"ff2f0db1",
			855 => x"08001f04",
			856 => x"013d0db1",
			857 => x"00013204",
			858 => x"00750db1",
			859 => x"00240db1",
			860 => x"0f00d914",
			861 => x"0600b310",
			862 => x"08001908",
			863 => x"05002b04",
			864 => x"ffd60db1",
			865 => x"fedf0db1",
			866 => x"09001c04",
			867 => x"ffab0db1",
			868 => x"00960db1",
			869 => x"ff380db1",
			870 => x"00d10db1",
			871 => x"02013904",
			872 => x"fede0db1",
			873 => x"0600bb04",
			874 => x"00810db1",
			875 => x"ffa70db1",
			876 => x"0200e914",
			877 => x"04000808",
			878 => x"04000704",
			879 => x"ffe40e55",
			880 => x"004c0e55",
			881 => x"05003604",
			882 => x"ff1f0e55",
			883 => x"00008904",
			884 => x"00350e55",
			885 => x"ffbb0e55",
			886 => x"01001138",
			887 => x"03002104",
			888 => x"ff7f0e55",
			889 => x"0600af20",
			890 => x"01000910",
			891 => x"04001d08",
			892 => x"09001904",
			893 => x"00b40e55",
			894 => x"001b0e55",
			895 => x"0c001404",
			896 => x"00490e55",
			897 => x"ff590e55",
			898 => x"02011d08",
			899 => x"01000d04",
			900 => x"00570e55",
			901 => x"ff620e55",
			902 => x"05002d04",
			903 => x"fffa0e55",
			904 => x"00eb0e55",
			905 => x"01000904",
			906 => x"00620e55",
			907 => x"0f00d908",
			908 => x"04002304",
			909 => x"ff350e55",
			910 => x"fff70e55",
			911 => x"0f00e004",
			912 => x"00530e55",
			913 => x"ffe20e55",
			914 => x"01002104",
			915 => x"ff390e55",
			916 => x"002b0e55",
			917 => x"00010e1c",
			918 => x"07002b18",
			919 => x"08001804",
			920 => x"ffa90f19",
			921 => x"0f008b10",
			922 => x"04000804",
			923 => x"002f0f19",
			924 => x"09001f04",
			925 => x"ffa40f19",
			926 => x"09002004",
			927 => x"00160f19",
			928 => x"ffee0f19",
			929 => x"005c0f19",
			930 => x"ff8a0f19",
			931 => x"0d001630",
			932 => x"07002b10",
			933 => x"0e007704",
			934 => x"00520f19",
			935 => x"04001804",
			936 => x"00080f19",
			937 => x"0600a004",
			938 => x"ffeb0f19",
			939 => x"ff720f19",
			940 => x"0a003214",
			941 => x"0e009810",
			942 => x"04001d08",
			943 => x"0b001404",
			944 => x"00130f19",
			945 => x"00a30f19",
			946 => x"08001c04",
			947 => x"ffeb0f19",
			948 => x"00700f19",
			949 => x"ffd50f19",
			950 => x"04002708",
			951 => x"0e008504",
			952 => x"00120f19",
			953 => x"ff970f19",
			954 => x"00330f19",
			955 => x"00011804",
			956 => x"005b0f19",
			957 => x"05002c04",
			958 => x"ff640f19",
			959 => x"0500380c",
			960 => x"02012504",
			961 => x"ffcf0f19",
			962 => x"04002304",
			963 => x"00810f19",
			964 => x"fffc0f19",
			965 => x"ff920f19",
			966 => x"0e00972c",
			967 => x"0a003e28",
			968 => x"09001504",
			969 => x"012c0f75",
			970 => x"03002104",
			971 => x"fe8b0f75",
			972 => x"0c001910",
			973 => x"08002008",
			974 => x"0a003604",
			975 => x"003e0f75",
			976 => x"ff020f75",
			977 => x"01000e04",
			978 => x"00090f75",
			979 => x"fe810f75",
			980 => x"0d001508",
			981 => x"01000a04",
			982 => x"fe300f75",
			983 => x"011e0f75",
			984 => x"09002004",
			985 => x"01b60f75",
			986 => x"003e0f75",
			987 => x"fea40f75",
			988 => x"fea40f75",
			989 => x"0b001528",
			990 => x"0600ae1c",
			991 => x"05003118",
			992 => x"02012f14",
			993 => x"0600a710",
			994 => x"09001908",
			995 => x"0b001204",
			996 => x"ff9d1059",
			997 => x"00c61059",
			998 => x"07002e04",
			999 => x"ff571059",
			1000 => x"01351059",
			1001 => x"01071059",
			1002 => x"ff031059",
			1003 => x"fe9f1059",
			1004 => x"0600b704",
			1005 => x"fe621059",
			1006 => x"08001c04",
			1007 => x"00f81059",
			1008 => x"fecc1059",
			1009 => x"00012b28",
			1010 => x"01000d1c",
			1011 => x"01000908",
			1012 => x"09001b04",
			1013 => x"00ce1059",
			1014 => x"fe8e1059",
			1015 => x"07002d08",
			1016 => x"0200d104",
			1017 => x"ff1c1059",
			1018 => x"01591059",
			1019 => x"07002f04",
			1020 => x"fe9b1059",
			1021 => x"00010704",
			1022 => x"ff491059",
			1023 => x"014c1059",
			1024 => x"0a003d04",
			1025 => x"fe6f1059",
			1026 => x"0600a004",
			1027 => x"ffb61059",
			1028 => x"00ba1059",
			1029 => x"03002604",
			1030 => x"ffa01059",
			1031 => x"0e008a08",
			1032 => x"01000a04",
			1033 => x"00171059",
			1034 => x"019d1059",
			1035 => x"03002e08",
			1036 => x"0e009404",
			1037 => x"01031059",
			1038 => x"ff071059",
			1039 => x"0a003608",
			1040 => x"05003404",
			1041 => x"ffbb1059",
			1042 => x"fe6d1059",
			1043 => x"01001404",
			1044 => x"00dd1059",
			1045 => x"ff061059",
			1046 => x"00010e24",
			1047 => x"0700291c",
			1048 => x"0b001510",
			1049 => x"04000804",
			1050 => x"0031115d",
			1051 => x"01000508",
			1052 => x"05002404",
			1053 => x"0031115d",
			1054 => x"ffcd115d",
			1055 => x"ff6e115d",
			1056 => x"07002604",
			1057 => x"ffcb115d",
			1058 => x"0c001704",
			1059 => x"0084115d",
			1060 => x"ffe4115d",
			1061 => x"09001a04",
			1062 => x"fff5115d",
			1063 => x"ff2d115d",
			1064 => x"0f00c028",
			1065 => x"09001908",
			1066 => x"07002904",
			1067 => x"002a115d",
			1068 => x"00ab115d",
			1069 => x"01000a08",
			1070 => x"0f00b404",
			1071 => x"002b115d",
			1072 => x"ff55115d",
			1073 => x"0400260c",
			1074 => x"01000d04",
			1075 => x"00c9115d",
			1076 => x"0f00ba04",
			1077 => x"ff9c115d",
			1078 => x"005b115d",
			1079 => x"03003404",
			1080 => x"ff76115d",
			1081 => x"03003804",
			1082 => x"005c115d",
			1083 => x"ffee115d",
			1084 => x"0f00c714",
			1085 => x"0400230c",
			1086 => x"0d001104",
			1087 => x"0015115d",
			1088 => x"0b001704",
			1089 => x"ff25115d",
			1090 => x"ffec115d",
			1091 => x"03003104",
			1092 => x"005b115d",
			1093 => x"ffd4115d",
			1094 => x"0e009314",
			1095 => x"05002a08",
			1096 => x"01000a04",
			1097 => x"0046115d",
			1098 => x"ff61115d",
			1099 => x"0600af08",
			1100 => x"0d001304",
			1101 => x"001f115d",
			1102 => x"00c4115d",
			1103 => x"000e115d",
			1104 => x"07003004",
			1105 => x"002c115d",
			1106 => x"09002204",
			1107 => x"ff47115d",
			1108 => x"0600b404",
			1109 => x"003e115d",
			1110 => x"ffdf115d",
			1111 => x"0200eb14",
			1112 => x"0d001404",
			1113 => x"fe6a1211",
			1114 => x"0c00170c",
			1115 => x"08001f08",
			1116 => x"07002604",
			1117 => x"ff171211",
			1118 => x"01b71211",
			1119 => x"fea91211",
			1120 => x"fe7f1211",
			1121 => x"07003844",
			1122 => x"0b001528",
			1123 => x"01000710",
			1124 => x"0c001408",
			1125 => x"00013004",
			1126 => x"01a91211",
			1127 => x"00741211",
			1128 => x"0e008204",
			1129 => x"ff1d1211",
			1130 => x"01001211",
			1131 => x"0600a80c",
			1132 => x"04002008",
			1133 => x"03002404",
			1134 => x"ff2f1211",
			1135 => x"00bd1211",
			1136 => x"feb41211",
			1137 => x"04001a08",
			1138 => x"00014604",
			1139 => x"fe961211",
			1140 => x"00bc1211",
			1141 => x"fe171211",
			1142 => x"0d001408",
			1143 => x"08001904",
			1144 => x"00191211",
			1145 => x"01701211",
			1146 => x"01000904",
			1147 => x"fe771211",
			1148 => x"00012a08",
			1149 => x"01000b04",
			1150 => x"010a1211",
			1151 => x"ff061211",
			1152 => x"0e009004",
			1153 => x"00fc1211",
			1154 => x"ff991211",
			1155 => x"fe821211",
			1156 => x"0d001230",
			1157 => x"0b00141c",
			1158 => x"03002410",
			1159 => x"0a00210c",
			1160 => x"03001104",
			1161 => x"005f1335",
			1162 => x"04001404",
			1163 => x"ff571335",
			1164 => x"ffe51335",
			1165 => x"00e31335",
			1166 => x"0f00bb04",
			1167 => x"00181335",
			1168 => x"0a003104",
			1169 => x"ff0d1335",
			1170 => x"ffe01335",
			1171 => x"0d001004",
			1172 => x"ffa41335",
			1173 => x"0600a10c",
			1174 => x"0a002a08",
			1175 => x"03002104",
			1176 => x"ffd01335",
			1177 => x"009c1335",
			1178 => x"ff551335",
			1179 => x"010f1335",
			1180 => x"04001e2c",
			1181 => x"0e00851c",
			1182 => x"0e007514",
			1183 => x"08001908",
			1184 => x"0b001504",
			1185 => x"00be1335",
			1186 => x"fff21335",
			1187 => x"05002308",
			1188 => x"07002804",
			1189 => x"ffbd1335",
			1190 => x"005b1335",
			1191 => x"ff4d1335",
			1192 => x"05002304",
			1193 => x"ffc71335",
			1194 => x"fed81335",
			1195 => x"09001d0c",
			1196 => x"0600ae04",
			1197 => x"00961335",
			1198 => x"0f00df04",
			1199 => x"fecb1335",
			1200 => x"00221335",
			1201 => x"00c71335",
			1202 => x"0a002f14",
			1203 => x"01000e0c",
			1204 => x"01000904",
			1205 => x"ffc81335",
			1206 => x"07002604",
			1207 => x"ffaa1335",
			1208 => x"01101335",
			1209 => x"0c001a04",
			1210 => x"ff441335",
			1211 => x"fff91335",
			1212 => x"0c00180c",
			1213 => x"08001804",
			1214 => x"00201335",
			1215 => x"00013204",
			1216 => x"fedc1335",
			1217 => x"ffb91335",
			1218 => x"05003208",
			1219 => x"0e009004",
			1220 => x"00d61335",
			1221 => x"ffc51335",
			1222 => x"0a003408",
			1223 => x"0a003204",
			1224 => x"ff1a1335",
			1225 => x"ffd51335",
			1226 => x"0e008904",
			1227 => x"ffa31335",
			1228 => x"00601335",
			1229 => x"0001112c",
			1230 => x"0c001504",
			1231 => x"ff711401",
			1232 => x"05002b14",
			1233 => x"0f008b04",
			1234 => x"ffd01401",
			1235 => x"09001d0c",
			1236 => x"05002204",
			1237 => x"fff21401",
			1238 => x"0e008404",
			1239 => x"00811401",
			1240 => x"fffa1401",
			1241 => x"ffdf1401",
			1242 => x"0e006f10",
			1243 => x"0d00150c",
			1244 => x"04002f08",
			1245 => x"03002904",
			1246 => x"fff91401",
			1247 => x"004b1401",
			1248 => x"ffea1401",
			1249 => x"ffd41401",
			1250 => x"ff8c1401",
			1251 => x"06009b08",
			1252 => x"01000b04",
			1253 => x"008f1401",
			1254 => x"00041401",
			1255 => x"02011d0c",
			1256 => x"02010f04",
			1257 => x"001c1401",
			1258 => x"0c001404",
			1259 => x"00021401",
			1260 => x"ff661401",
			1261 => x"0600a814",
			1262 => x"0100090c",
			1263 => x"0c001404",
			1264 => x"004f1401",
			1265 => x"02012c04",
			1266 => x"ff911401",
			1267 => x"000c1401",
			1268 => x"05003804",
			1269 => x"009c1401",
			1270 => x"fff61401",
			1271 => x"01000704",
			1272 => x"00521401",
			1273 => x"00014508",
			1274 => x"05003404",
			1275 => x"ff5b1401",
			1276 => x"fff41401",
			1277 => x"07003204",
			1278 => x"00491401",
			1279 => x"ffbc1401",
			1280 => x"04002644",
			1281 => x"04002540",
			1282 => x"09001f2c",
			1283 => x"01000d20",
			1284 => x"09001b10",
			1285 => x"0600a908",
			1286 => x"0d001404",
			1287 => x"005a14bd",
			1288 => x"ff2114bd",
			1289 => x"01000804",
			1290 => x"fffb14bd",
			1291 => x"fec814bd",
			1292 => x"0e007c08",
			1293 => x"0a002c04",
			1294 => x"001414bd",
			1295 => x"ff1d14bd",
			1296 => x"0a003204",
			1297 => x"00db14bd",
			1298 => x"ff9714bd",
			1299 => x"02012608",
			1300 => x"03001d04",
			1301 => x"004f14bd",
			1302 => x"fed414bd",
			1303 => x"003514bd",
			1304 => x"0a003610",
			1305 => x"0600a60c",
			1306 => x"07003104",
			1307 => x"ff8314bd",
			1308 => x"0f00a904",
			1309 => x"ffe914bd",
			1310 => x"009514bd",
			1311 => x"fec314bd",
			1312 => x"005c14bd",
			1313 => x"011214bd",
			1314 => x"04002804",
			1315 => x"feec14bd",
			1316 => x"00012e0c",
			1317 => x"01000a08",
			1318 => x"01000904",
			1319 => x"ff6714bd",
			1320 => x"00b514bd",
			1321 => x"fee114bd",
			1322 => x"05003b08",
			1323 => x"0e009304",
			1324 => x"00de14bd",
			1325 => x"ff8b14bd",
			1326 => x"ff5614bd",
			1327 => x"0f00c058",
			1328 => x"00010e34",
			1329 => x"04001c1c",
			1330 => x"04001a10",
			1331 => x"04000808",
			1332 => x"04000704",
			1333 => x"ffee15e1",
			1334 => x"003215e1",
			1335 => x"0f00ac04",
			1336 => x"ffae15e1",
			1337 => x"000115e1",
			1338 => x"07002704",
			1339 => x"fff615e1",
			1340 => x"07002e04",
			1341 => x"005715e1",
			1342 => x"fff715e1",
			1343 => x"09001f08",
			1344 => x"0e007b04",
			1345 => x"ff8415e1",
			1346 => x"fffa15e1",
			1347 => x"0b00180c",
			1348 => x"0b001704",
			1349 => x"ffeb15e1",
			1350 => x"09002004",
			1351 => x"003b15e1",
			1352 => x"fffc15e1",
			1353 => x"ffd915e1",
			1354 => x"04002614",
			1355 => x"0a002804",
			1356 => x"fffa15e1",
			1357 => x"01000604",
			1358 => x"000315e1",
			1359 => x"01000d04",
			1360 => x"009f15e1",
			1361 => x"0d001a04",
			1362 => x"002215e1",
			1363 => x"ffec15e1",
			1364 => x"03003408",
			1365 => x"0e008a04",
			1366 => x"ffa415e1",
			1367 => x"000115e1",
			1368 => x"03003804",
			1369 => x"004215e1",
			1370 => x"ffe915e1",
			1371 => x"0f00c714",
			1372 => x"0d001208",
			1373 => x"0a002d04",
			1374 => x"002b15e1",
			1375 => x"ffaf15e1",
			1376 => x"05003604",
			1377 => x"ff5d15e1",
			1378 => x"05003b04",
			1379 => x"001515e1",
			1380 => x"ffea15e1",
			1381 => x"01000704",
			1382 => x"006a15e1",
			1383 => x"0c001810",
			1384 => x"0001570c",
			1385 => x"0600ae04",
			1386 => x"fff215e1",
			1387 => x"04001604",
			1388 => x"fff315e1",
			1389 => x"ff6215e1",
			1390 => x"001c15e1",
			1391 => x"0001470c",
			1392 => x"05003808",
			1393 => x"0600b404",
			1394 => x"008815e1",
			1395 => x"fff715e1",
			1396 => x"ffe215e1",
			1397 => x"03002d04",
			1398 => x"001815e1",
			1399 => x"ffaf15e1",
			1400 => x"0700374c",
			1401 => x"0e009648",
			1402 => x"0e008128",
			1403 => x"09001914",
			1404 => x"04001b0c",
			1405 => x"0a002508",
			1406 => x"05001104",
			1407 => x"011a168d",
			1408 => x"ff17168d",
			1409 => x"0151168d",
			1410 => x"03002604",
			1411 => x"ff1d168d",
			1412 => x"0027168d",
			1413 => x"01000604",
			1414 => x"fe81168d",
			1415 => x"04002108",
			1416 => x"05002604",
			1417 => x"0045168d",
			1418 => x"ff44168d",
			1419 => x"0a003604",
			1420 => x"0107168d",
			1421 => x"ff5a168d",
			1422 => x"00012a0c",
			1423 => x"00011608",
			1424 => x"0f00b204",
			1425 => x"ff67168d",
			1426 => x"00d3168d",
			1427 => x"fe89168d",
			1428 => x"0600a808",
			1429 => x"02012904",
			1430 => x"0172168d",
			1431 => x"001b168d",
			1432 => x"01000704",
			1433 => x"0110168d",
			1434 => x"05002c04",
			1435 => x"ff03168d",
			1436 => x"0089168d",
			1437 => x"feb2168d",
			1438 => x"02013904",
			1439 => x"fe97168d",
			1440 => x"02013b04",
			1441 => x"00fe168d",
			1442 => x"ff6a168d",
			1443 => x"0f008b10",
			1444 => x"09001504",
			1445 => x"00691741",
			1446 => x"0c001708",
			1447 => x"09001e04",
			1448 => x"fe661741",
			1449 => x"00d51741",
			1450 => x"fe631741",
			1451 => x"09002348",
			1452 => x"0600a830",
			1453 => x"01000918",
			1454 => x"0c001408",
			1455 => x"00012204",
			1456 => x"008e1741",
			1457 => x"02b01741",
			1458 => x"03002708",
			1459 => x"05002304",
			1460 => x"fe451741",
			1461 => x"012d1741",
			1462 => x"00011404",
			1463 => x"ff461741",
			1464 => x"fe241741",
			1465 => x"00012a10",
			1466 => x"01000d08",
			1467 => x"0c001604",
			1468 => x"00571741",
			1469 => x"02c91741",
			1470 => x"0a002c04",
			1471 => x"ffa61741",
			1472 => x"fe991741",
			1473 => x"0d001704",
			1474 => x"03001741",
			1475 => x"01c31741",
			1476 => x"0f00c708",
			1477 => x"07003404",
			1478 => x"fdbe1741",
			1479 => x"ff271741",
			1480 => x"0b001304",
			1481 => x"fe421741",
			1482 => x"01000704",
			1483 => x"02f11741",
			1484 => x"02013104",
			1485 => x"fef51741",
			1486 => x"015e1741",
			1487 => x"fe651741",
			1488 => x"0d001230",
			1489 => x"0b00141c",
			1490 => x"03002410",
			1491 => x"0a00210c",
			1492 => x"03001104",
			1493 => x"005a1885",
			1494 => x"04001404",
			1495 => x"ff5f1885",
			1496 => x"ffe61885",
			1497 => x"00d51885",
			1498 => x"0f00bb04",
			1499 => x"00161885",
			1500 => x"0a003104",
			1501 => x"ff181885",
			1502 => x"ffe11885",
			1503 => x"04002110",
			1504 => x"03002408",
			1505 => x"09001904",
			1506 => x"00191885",
			1507 => x"ff7b1885",
			1508 => x"05002c04",
			1509 => x"01081885",
			1510 => x"00641885",
			1511 => x"ff731885",
			1512 => x"04001e2c",
			1513 => x"0e00851c",
			1514 => x"0e007514",
			1515 => x"08001908",
			1516 => x"0b001504",
			1517 => x"00b71885",
			1518 => x"fff31885",
			1519 => x"05002308",
			1520 => x"0a002504",
			1521 => x"ffb91885",
			1522 => x"00601885",
			1523 => x"ff551885",
			1524 => x"05002304",
			1525 => x"ffcc1885",
			1526 => x"fee51885",
			1527 => x"09001d0c",
			1528 => x"0600ae04",
			1529 => x"008d1885",
			1530 => x"0f00df04",
			1531 => x"fed41885",
			1532 => x"00201885",
			1533 => x"00c01885",
			1534 => x"05003220",
			1535 => x"0600930c",
			1536 => x"07002808",
			1537 => x"01000a04",
			1538 => x"00711885",
			1539 => x"ffc41885",
			1540 => x"ff191885",
			1541 => x"0700320c",
			1542 => x"08001904",
			1543 => x"00271885",
			1544 => x"0f00bd04",
			1545 => x"00651885",
			1546 => x"012f1885",
			1547 => x"03002c04",
			1548 => x"ff2c1885",
			1549 => x"00461885",
			1550 => x"05003610",
			1551 => x"0f00c808",
			1552 => x"01001004",
			1553 => x"fec61885",
			1554 => x"ffee1885",
			1555 => x"0e009604",
			1556 => x"00a71885",
			1557 => x"ff9a1885",
			1558 => x"05003708",
			1559 => x"08002404",
			1560 => x"00f51885",
			1561 => x"ffa51885",
			1562 => x"00011808",
			1563 => x"0f009c04",
			1564 => x"ff731885",
			1565 => x"00b31885",
			1566 => x"0b001804",
			1567 => x"ff1c1885",
			1568 => x"ffdd1885",
			1569 => x"0b001208",
			1570 => x"0c001004",
			1571 => x"ffc11939",
			1572 => x"fe8d1939",
			1573 => x"04001618",
			1574 => x"01000504",
			1575 => x"fedb1939",
			1576 => x"0c001710",
			1577 => x"0e00960c",
			1578 => x"06004404",
			1579 => x"ffcc1939",
			1580 => x"01000a04",
			1581 => x"01a21939",
			1582 => x"00c91939",
			1583 => x"ff831939",
			1584 => x"fefa1939",
			1585 => x"0a003b34",
			1586 => x"0600b11c",
			1587 => x"0f00c710",
			1588 => x"0600a808",
			1589 => x"03002404",
			1590 => x"ff401939",
			1591 => x"00521939",
			1592 => x"05003604",
			1593 => x"fe451939",
			1594 => x"ffc01939",
			1595 => x"0c001504",
			1596 => x"fe441939",
			1597 => x"00014204",
			1598 => x"015e1939",
			1599 => x"00411939",
			1600 => x"0f00d90c",
			1601 => x"0e009504",
			1602 => x"fe571939",
			1603 => x"02013904",
			1604 => x"febd1939",
			1605 => x"011e1939",
			1606 => x"00015808",
			1607 => x"0600c304",
			1608 => x"01871939",
			1609 => x"ff5f1939",
			1610 => x"ff091939",
			1611 => x"05003d04",
			1612 => x"fffd1939",
			1613 => x"fe811939",
			1614 => x"0b00154c",
			1615 => x"09001924",
			1616 => x"0600a81c",
			1617 => x"04002018",
			1618 => x"00011910",
			1619 => x"08001808",
			1620 => x"0e006f04",
			1621 => x"feea1a75",
			1622 => x"ffdb1a75",
			1623 => x"01000804",
			1624 => x"01011a75",
			1625 => x"ff551a75",
			1626 => x"0600a004",
			1627 => x"015d1a75",
			1628 => x"00931a75",
			1629 => x"ff461a75",
			1630 => x"08001904",
			1631 => x"ffbf1a75",
			1632 => x"fedd1a75",
			1633 => x"02012b1c",
			1634 => x"0e00750c",
			1635 => x"05002608",
			1636 => x"05002204",
			1637 => x"ffa41a75",
			1638 => x"00f41a75",
			1639 => x"ff191a75",
			1640 => x"0e008104",
			1641 => x"fe7d1a75",
			1642 => x"0600a404",
			1643 => x"00df1a75",
			1644 => x"0a003104",
			1645 => x"fe981a75",
			1646 => x"00811a75",
			1647 => x"03002904",
			1648 => x"00db1a75",
			1649 => x"05002e04",
			1650 => x"fee01a75",
			1651 => x"005f1a75",
			1652 => x"0f00bb2c",
			1653 => x"01000d20",
			1654 => x"01000904",
			1655 => x"fed81a75",
			1656 => x"05003610",
			1657 => x"07002c08",
			1658 => x"0d001504",
			1659 => x"01081a75",
			1660 => x"ff3b1a75",
			1661 => x"0b001804",
			1662 => x"ff351a75",
			1663 => x"006e1a75",
			1664 => x"0a003d08",
			1665 => x"04003304",
			1666 => x"01511a75",
			1667 => x"ffd41a75",
			1668 => x"ff721a75",
			1669 => x"03003404",
			1670 => x"feb01a75",
			1671 => x"03003804",
			1672 => x"00931a75",
			1673 => x"ffa11a75",
			1674 => x"0600b414",
			1675 => x"0b001604",
			1676 => x"013c1a75",
			1677 => x"01000c04",
			1678 => x"ffae1a75",
			1679 => x"0d001804",
			1680 => x"016a1a75",
			1681 => x"05003404",
			1682 => x"ff501a75",
			1683 => x"00af1a75",
			1684 => x"0f00d90c",
			1685 => x"0a003604",
			1686 => x"feaf1a75",
			1687 => x"0600b704",
			1688 => x"00b31a75",
			1689 => x"ff731a75",
			1690 => x"04002104",
			1691 => x"01241a75",
			1692 => x"ff9f1a75",
			1693 => x"07003378",
			1694 => x"0b00153c",
			1695 => x"09001920",
			1696 => x"0b001418",
			1697 => x"06009d0c",
			1698 => x"06004404",
			1699 => x"ffa91b99",
			1700 => x"00011004",
			1701 => x"00191b99",
			1702 => x"00b61b99",
			1703 => x"07002d08",
			1704 => x"03002404",
			1705 => x"ffe51b99",
			1706 => x"ff331b99",
			1707 => x"002b1b99",
			1708 => x"00011e04",
			1709 => x"ffda1b99",
			1710 => x"00b31b99",
			1711 => x"02012b14",
			1712 => x"07002e0c",
			1713 => x"0e007508",
			1714 => x"06007b04",
			1715 => x"ff9c1b99",
			1716 => x"00341b99",
			1717 => x"ff141b99",
			1718 => x"04001a04",
			1719 => x"ffd51b99",
			1720 => x"006a1b99",
			1721 => x"03002904",
			1722 => x"008e1b99",
			1723 => x"ffbe1b99",
			1724 => x"0a003120",
			1725 => x"01000d18",
			1726 => x"0a00280c",
			1727 => x"0d001204",
			1728 => x"007d1b99",
			1729 => x"0b001704",
			1730 => x"ff641b99",
			1731 => x"00451b99",
			1732 => x"0b001908",
			1733 => x"0000f304",
			1734 => x"00251b99",
			1735 => x"010e1b99",
			1736 => x"ffc71b99",
			1737 => x"05002c04",
			1738 => x"ff321b99",
			1739 => x"00601b99",
			1740 => x"08001d0c",
			1741 => x"04002e04",
			1742 => x"ff331b99",
			1743 => x"05004704",
			1744 => x"003b1b99",
			1745 => x"ffd41b99",
			1746 => x"0f00ba0c",
			1747 => x"01000b04",
			1748 => x"00591b99",
			1749 => x"03003404",
			1750 => x"ff6f1b99",
			1751 => x"00111b99",
			1752 => x"00ab1b99",
			1753 => x"0a003604",
			1754 => x"ff2c1b99",
			1755 => x"0001370c",
			1756 => x"05003a04",
			1757 => x"00c41b99",
			1758 => x"0e008d04",
			1759 => x"ffb31b99",
			1760 => x"00011b99",
			1761 => x"02013904",
			1762 => x"ff7b1b99",
			1763 => x"02013e04",
			1764 => x"00521b99",
			1765 => x"fff11b99",
			1766 => x"0400080c",
			1767 => x"04000704",
			1768 => x"ff261c55",
			1769 => x"03001004",
			1770 => x"0b901c55",
			1771 => x"ff731c55",
			1772 => x"09002350",
			1773 => x"03002720",
			1774 => x"08001d18",
			1775 => x"0600ae10",
			1776 => x"0e008108",
			1777 => x"06009f04",
			1778 => x"00491c55",
			1779 => x"ff031c55",
			1780 => x"07002e04",
			1781 => x"01631c55",
			1782 => x"ff9b1c55",
			1783 => x"04001704",
			1784 => x"00741c55",
			1785 => x"fe761c55",
			1786 => x"03002604",
			1787 => x"fde21c55",
			1788 => x"00151c55",
			1789 => x"0201211c",
			1790 => x"0e007d10",
			1791 => x"01000b08",
			1792 => x"08001d04",
			1793 => x"00361c55",
			1794 => x"02651c55",
			1795 => x"0a002d04",
			1796 => x"ffcd1c55",
			1797 => x"fe721c55",
			1798 => x"0a003708",
			1799 => x"07002f04",
			1800 => x"fe351c55",
			1801 => x"ff091c55",
			1802 => x"fff71c55",
			1803 => x"07002b04",
			1804 => x"fe711c55",
			1805 => x"0600a808",
			1806 => x"02012d04",
			1807 => x"01bf1c55",
			1808 => x"fff91c55",
			1809 => x"03002f04",
			1810 => x"00bf1c55",
			1811 => x"ff441c55",
			1812 => x"fe871c55",
			1813 => x"02011f58",
			1814 => x"01000d4c",
			1815 => x"0a002f30",
			1816 => x"0a00281c",
			1817 => x"0d001210",
			1818 => x"08001808",
			1819 => x"07002904",
			1820 => x"ff2e1d59",
			1821 => x"00a91d59",
			1822 => x"0f004b04",
			1823 => x"ffa71d59",
			1824 => x"00eb1d59",
			1825 => x"08001b04",
			1826 => x"feb31d59",
			1827 => x"09001a04",
			1828 => x"00941d59",
			1829 => x"ff501d59",
			1830 => x"0e007e0c",
			1831 => x"0d001508",
			1832 => x"0c001804",
			1833 => x"01701d59",
			1834 => x"ffdd1d59",
			1835 => x"ffe71d59",
			1836 => x"0f00b804",
			1837 => x"ffe51d59",
			1838 => x"fedb1d59",
			1839 => x"08001f14",
			1840 => x"0f00b60c",
			1841 => x"0d001804",
			1842 => x"fea01d59",
			1843 => x"05005c04",
			1844 => x"00791d59",
			1845 => x"fffc1d59",
			1846 => x"00011f04",
			1847 => x"ffc61d59",
			1848 => x"005a1d59",
			1849 => x"0200ef04",
			1850 => x"ffe51d59",
			1851 => x"00be1d59",
			1852 => x"0a003d04",
			1853 => x"fe9e1d59",
			1854 => x"0e008804",
			1855 => x"ffe31d59",
			1856 => x"00601d59",
			1857 => x"0f00bc04",
			1858 => x"01341d59",
			1859 => x"0e007e04",
			1860 => x"ff201d59",
			1861 => x"0d001814",
			1862 => x"0600a504",
			1863 => x"00f11d59",
			1864 => x"0c001408",
			1865 => x"07002f04",
			1866 => x"feb11d59",
			1867 => x"006f1d59",
			1868 => x"07002e04",
			1869 => x"00bd1d59",
			1870 => x"00091d59",
			1871 => x"03002704",
			1872 => x"febf1d59",
			1873 => x"08002204",
			1874 => x"00ab1d59",
			1875 => x"0f00c004",
			1876 => x"007e1d59",
			1877 => x"fec71d59",
			1878 => x"0e009780",
			1879 => x"00013154",
			1880 => x"0600a03c",
			1881 => x"0a002f20",
			1882 => x"0a002810",
			1883 => x"07002d08",
			1884 => x"0e007604",
			1885 => x"001c1e5f",
			1886 => x"fedd1e5f",
			1887 => x"08001d04",
			1888 => x"010a1e5f",
			1889 => x"ffdc1e5f",
			1890 => x"05002a08",
			1891 => x"07002c04",
			1892 => x"015a1e5f",
			1893 => x"ffd21e5f",
			1894 => x"0d001504",
			1895 => x"00931e5f",
			1896 => x"ff401e5f",
			1897 => x"01000b10",
			1898 => x"08001d08",
			1899 => x"0f00a904",
			1900 => x"ff0d1e5f",
			1901 => x"001f1e5f",
			1902 => x"06008304",
			1903 => x"ffdc1e5f",
			1904 => x"00ee1e5f",
			1905 => x"07002f04",
			1906 => x"fec61e5f",
			1907 => x"03003104",
			1908 => x"00321e5f",
			1909 => x"ffbd1e5f",
			1910 => x"0b001704",
			1911 => x"fec41e5f",
			1912 => x"04002608",
			1913 => x"0600a704",
			1914 => x"00f21e5f",
			1915 => x"fff61e5f",
			1916 => x"0e008a04",
			1917 => x"ff121e5f",
			1918 => x"04002d04",
			1919 => x"00861e5f",
			1920 => x"fff71e5f",
			1921 => x"0600a910",
			1922 => x"00013b0c",
			1923 => x"01000a08",
			1924 => x"02012904",
			1925 => x"00b51e5f",
			1926 => x"ffe01e5f",
			1927 => x"01201e5f",
			1928 => x"ff891e5f",
			1929 => x"01000704",
			1930 => x"00a61e5f",
			1931 => x"05002c08",
			1932 => x"03002404",
			1933 => x"ffbc1e5f",
			1934 => x"fed01e5f",
			1935 => x"08002208",
			1936 => x"01000c04",
			1937 => x"00061e5f",
			1938 => x"00e61e5f",
			1939 => x"04002804",
			1940 => x"ff1e1e5f",
			1941 => x"00571e5f",
			1942 => x"ff0b1e5f",
			1943 => x"0e00971c",
			1944 => x"0f004b04",
			1945 => x"fee31e99",
			1946 => x"09001704",
			1947 => x"01141e99",
			1948 => x"03002104",
			1949 => x"fec61e99",
			1950 => x"08001504",
			1951 => x"fed61e99",
			1952 => x"07002604",
			1953 => x"fee21e99",
			1954 => x"0f00c004",
			1955 => x"00511e99",
			1956 => x"fffa1e99",
			1957 => x"fedd1e99",
			1958 => x"0f008b10",
			1959 => x"09001504",
			1960 => x"00621ef5",
			1961 => x"0c001708",
			1962 => x"09001e04",
			1963 => x"fe641ef5",
			1964 => x"00df1ef5",
			1965 => x"fe621ef5",
			1966 => x"0900231c",
			1967 => x"0e009718",
			1968 => x"0d000f04",
			1969 => x"022d1ef5",
			1970 => x"04001504",
			1971 => x"fe4b1ef5",
			1972 => x"0b001308",
			1973 => x"0600a004",
			1974 => x"01791ef5",
			1975 => x"fe1d1ef5",
			1976 => x"00012a04",
			1977 => x"00ae1ef5",
			1978 => x"017b1ef5",
			1979 => x"fe721ef5",
			1980 => x"fe641ef5",
			1981 => x"0e009720",
			1982 => x"0f004b04",
			1983 => x"ff271f39",
			1984 => x"09001704",
			1985 => x"00bf1f39",
			1986 => x"03002104",
			1987 => x"ff051f39",
			1988 => x"08001504",
			1989 => x"ff1c1f39",
			1990 => x"0a003108",
			1991 => x"01000d04",
			1992 => x"005c1f39",
			1993 => x"ff611f39",
			1994 => x"01000804",
			1995 => x"feb81f39",
			1996 => x"00211f39",
			1997 => x"ff151f39",
			1998 => x"0400262c",
			1999 => x"04002528",
			2000 => x"08002218",
			2001 => x"0a003614",
			2002 => x"05003210",
			2003 => x"0c001808",
			2004 => x"01000d04",
			2005 => x"00081fc5",
			2006 => x"ff3a1fc5",
			2007 => x"04001a04",
			2008 => x"ff031fc5",
			2009 => x"00c91fc5",
			2010 => x"ff101fc5",
			2011 => x"010d1fc5",
			2012 => x"04001b0c",
			2013 => x"07003104",
			2014 => x"ff981fc5",
			2015 => x"07003304",
			2016 => x"00891fc5",
			2017 => x"ffed1fc5",
			2018 => x"fec41fc5",
			2019 => x"01301fc5",
			2020 => x"04002e0c",
			2021 => x"0b001804",
			2022 => x"fed21fc5",
			2023 => x"0b001a04",
			2024 => x"00c61fc5",
			2025 => x"fef71fc5",
			2026 => x"0400320c",
			2027 => x"0f009c04",
			2028 => x"ff7a1fc5",
			2029 => x"03003504",
			2030 => x"01141fc5",
			2031 => x"fff31fc5",
			2032 => x"ff111fc5",
			2033 => x"02010518",
			2034 => x"0f008b10",
			2035 => x"09001504",
			2036 => x"ffe32049",
			2037 => x"0c001708",
			2038 => x"0c001604",
			2039 => x"fe5d2049",
			2040 => x"feef2049",
			2041 => x"fe5a2049",
			2042 => x"07002b04",
			2043 => x"01822049",
			2044 => x"fe5c2049",
			2045 => x"09002328",
			2046 => x"0600bb24",
			2047 => x"0600a814",
			2048 => x"0b001810",
			2049 => x"09001908",
			2050 => x"0f00c004",
			2051 => x"04d02049",
			2052 => x"01db2049",
			2053 => x"02011d04",
			2054 => x"00612049",
			2055 => x"02f22049",
			2056 => x"04e62049",
			2057 => x"02012804",
			2058 => x"fe402049",
			2059 => x"01000704",
			2060 => x"04a52049",
			2061 => x"09001c04",
			2062 => x"ff1e2049",
			2063 => x"02982049",
			2064 => x"fe5e2049",
			2065 => x"fe5b2049",
			2066 => x"0200e914",
			2067 => x"01000a04",
			2068 => x"fe5f20ed",
			2069 => x"0c00170c",
			2070 => x"01000e08",
			2071 => x"07002604",
			2072 => x"fec120ed",
			2073 => x"025520ed",
			2074 => x"fe9120ed",
			2075 => x"fe7920ed",
			2076 => x"0d001834",
			2077 => x"0600af20",
			2078 => x"0f00c614",
			2079 => x"0f00c410",
			2080 => x"09001908",
			2081 => x"0a002504",
			2082 => x"001820ed",
			2083 => x"015d20ed",
			2084 => x"01000604",
			2085 => x"fec720ed",
			2086 => x"007920ed",
			2087 => x"feb920ed",
			2088 => x"0c001504",
			2089 => x"fe7a20ed",
			2090 => x"0d001304",
			2091 => x"016320ed",
			2092 => x"021420ed",
			2093 => x"0201340c",
			2094 => x"07003204",
			2095 => x"fdfb20ed",
			2096 => x"0d001404",
			2097 => x"ff2120ed",
			2098 => x"003620ed",
			2099 => x"0f00d904",
			2100 => x"fffe20ed",
			2101 => x"016020ed",
			2102 => x"0c001904",
			2103 => x"fe6d20ed",
			2104 => x"09002204",
			2105 => x"014b20ed",
			2106 => x"fe7220ed",
			2107 => x"0200e914",
			2108 => x"01000a04",
			2109 => x"fe632181",
			2110 => x"0c00170c",
			2111 => x"01000e08",
			2112 => x"07002604",
			2113 => x"fecd2181",
			2114 => x"020a2181",
			2115 => x"fe992181",
			2116 => x"fe7d2181",
			2117 => x"0d00182c",
			2118 => x"0e007404",
			2119 => x"01872181",
			2120 => x"02011d10",
			2121 => x"0a00310c",
			2122 => x"0600a108",
			2123 => x"06009904",
			2124 => x"ffd82181",
			2125 => x"00f22181",
			2126 => x"fe5f2181",
			2127 => x"fe1e2181",
			2128 => x"07002b08",
			2129 => x"0c001404",
			2130 => x"00692181",
			2131 => x"feaa2181",
			2132 => x"0600af08",
			2133 => x"0e008804",
			2134 => x"00f32181",
			2135 => x"01cb2181",
			2136 => x"00014404",
			2137 => x"feeb2181",
			2138 => x"00702181",
			2139 => x"0c001904",
			2140 => x"fe8c2181",
			2141 => x"09002204",
			2142 => x"01322181",
			2143 => x"fe762181",
			2144 => x"0400080c",
			2145 => x"04000704",
			2146 => x"ff5521f5",
			2147 => x"09001d04",
			2148 => x"022121f5",
			2149 => x"ffa121f5",
			2150 => x"0a003e2c",
			2151 => x"0e004d04",
			2152 => x"fea221f5",
			2153 => x"0e007810",
			2154 => x"0001110c",
			2155 => x"0c001504",
			2156 => x"fe7e21f5",
			2157 => x"0d001504",
			2158 => x"011921f5",
			2159 => x"ff3c21f5",
			2160 => x"019a21f5",
			2161 => x"0e007c08",
			2162 => x"0c001504",
			2163 => x"008521f5",
			2164 => x"fe4e21f5",
			2165 => x"0b001408",
			2166 => x"03002604",
			2167 => x"006221f5",
			2168 => x"fed021f5",
			2169 => x"07002d04",
			2170 => x"00f321f5",
			2171 => x"000a21f5",
			2172 => x"fe9821f5",
			2173 => x"0200eb14",
			2174 => x"0d001404",
			2175 => x"fe662281",
			2176 => x"0c00170c",
			2177 => x"08001f08",
			2178 => x"07002604",
			2179 => x"ff0f2281",
			2180 => x"01e42281",
			2181 => x"fea12281",
			2182 => x"fe7c2281",
			2183 => x"07003830",
			2184 => x"0b001820",
			2185 => x"0800221c",
			2186 => x"0f00b50c",
			2187 => x"01000a08",
			2188 => x"0c001504",
			2189 => x"00782281",
			2190 => x"01ad2281",
			2191 => x"ffaf2281",
			2192 => x"02011c08",
			2193 => x"03002704",
			2194 => x"ff792281",
			2195 => x"fe212281",
			2196 => x"05002e04",
			2197 => x"ffee2281",
			2198 => x"00e42281",
			2199 => x"fe8b2281",
			2200 => x"0100140c",
			2201 => x"05003404",
			2202 => x"00522281",
			2203 => x"04002d04",
			2204 => x"01c62281",
			2205 => x"fedb2281",
			2206 => x"fe8e2281",
			2207 => x"fe7d2281",
			2208 => x"09001504",
			2209 => x"025c22d5",
			2210 => x"03002104",
			2211 => x"fe6a22d5",
			2212 => x"04003220",
			2213 => x"0100131c",
			2214 => x"0600ae10",
			2215 => x"09001908",
			2216 => x"00013c04",
			2217 => x"014b22d5",
			2218 => x"fe7a22d5",
			2219 => x"01000904",
			2220 => x"ff9c22d5",
			2221 => x"008422d5",
			2222 => x"00013604",
			2223 => x"fde222d5",
			2224 => x"0f00d904",
			2225 => x"ffe922d5",
			2226 => x"012d22d5",
			2227 => x"fe7022d5",
			2228 => x"fe6d22d5",
			2229 => x"00010a18",
			2230 => x"0f008b10",
			2231 => x"09001504",
			2232 => x"ffd52369",
			2233 => x"0c001708",
			2234 => x"0c001604",
			2235 => x"fe582369",
			2236 => x"fecc2369",
			2237 => x"fe552369",
			2238 => x"07002c04",
			2239 => x"03c82369",
			2240 => x"fe592369",
			2241 => x"09002330",
			2242 => x"0e00972c",
			2243 => x"0c00181c",
			2244 => x"03002c10",
			2245 => x"02012f08",
			2246 => x"0a002304",
			2247 => x"00f72369",
			2248 => x"06f42369",
			2249 => x"0e008b04",
			2250 => x"ff022369",
			2251 => x"05c12369",
			2252 => x"04002608",
			2253 => x"0e008204",
			2254 => x"05042369",
			2255 => x"ffcb2369",
			2256 => x"fe592369",
			2257 => x"0800230c",
			2258 => x"02011e04",
			2259 => x"03972369",
			2260 => x"01000c04",
			2261 => x"06e52369",
			2262 => x"099e2369",
			2263 => x"01552369",
			2264 => x"fe602369",
			2265 => x"fe562369",
			2266 => x"00010e04",
			2267 => x"ff8d240d",
			2268 => x"0a003128",
			2269 => x"0d001820",
			2270 => x"07002c14",
			2271 => x"0600a008",
			2272 => x"0a002804",
			2273 => x"ffe8240d",
			2274 => x"006d240d",
			2275 => x"03002608",
			2276 => x"0f00c904",
			2277 => x"0040240d",
			2278 => x"ffda240d",
			2279 => x"ffa3240d",
			2280 => x"0f00d204",
			2281 => x"007d240d",
			2282 => x"0f00d904",
			2283 => x"ffd8240d",
			2284 => x"0041240d",
			2285 => x"00013404",
			2286 => x"ffc0240d",
			2287 => x"0012240d",
			2288 => x"0b001814",
			2289 => x"0f00c80c",
			2290 => x"0e008208",
			2291 => x"0e007f04",
			2292 => x"ffe5240d",
			2293 => x"0014240d",
			2294 => x"ff97240d",
			2295 => x"0e009304",
			2296 => x"0032240d",
			2297 => x"ffce240d",
			2298 => x"0d001a08",
			2299 => x"0e008e04",
			2300 => x"0066240d",
			2301 => x"fffe240d",
			2302 => x"04002308",
			2303 => x"00013904",
			2304 => x"0027240d",
			2305 => x"fff0240d",
			2306 => x"ffbe240d",
			2307 => x"0200ef10",
			2308 => x"0c00170c",
			2309 => x"0c001604",
			2310 => x"fe5324a1",
			2311 => x"01000a04",
			2312 => x"fe8f24a1",
			2313 => x"01ce24a1",
			2314 => x"fe6b24a1",
			2315 => x"0d001b34",
			2316 => x"0a003e30",
			2317 => x"0f00c014",
			2318 => x"02011f0c",
			2319 => x"01000d08",
			2320 => x"08001b04",
			2321 => x"005d24a1",
			2322 => x"014a24a1",
			2323 => x"feeb24a1",
			2324 => x"01000904",
			2325 => x"007624a1",
			2326 => x"022024a1",
			2327 => x"02012b10",
			2328 => x"0b001508",
			2329 => x"03002604",
			2330 => x"ff3e24a1",
			2331 => x"fded24a1",
			2332 => x"08001f04",
			2333 => x"01c924a1",
			2334 => x"feb324a1",
			2335 => x"00013b04",
			2336 => x"018f24a1",
			2337 => x"0f00c804",
			2338 => x"febe24a1",
			2339 => x"00a224a1",
			2340 => x"fe5324a1",
			2341 => x"01001204",
			2342 => x"006924a1",
			2343 => x"fe6b24a1",
			2344 => x"0f008b14",
			2345 => x"09001504",
			2346 => x"01892545",
			2347 => x"0c00170c",
			2348 => x"08001d04",
			2349 => x"fe6b2545",
			2350 => x"0d001504",
			2351 => x"04132545",
			2352 => x"fea72545",
			2353 => x"fe672545",
			2354 => x"08002338",
			2355 => x"03003530",
			2356 => x"0c00181c",
			2357 => x"0a002f10",
			2358 => x"0600a008",
			2359 => x"0a002104",
			2360 => x"ff622545",
			2361 => x"01892545",
			2362 => x"00013104",
			2363 => x"fea92545",
			2364 => x"00aa2545",
			2365 => x"02012104",
			2366 => x"fe2c2545",
			2367 => x"0a003404",
			2368 => x"00b12545",
			2369 => x"fec22545",
			2370 => x"00012a08",
			2371 => x"05002f04",
			2372 => x"fe4d2545",
			2373 => x"00dc2545",
			2374 => x"01000c04",
			2375 => x"00a02545",
			2376 => x"0f00ce04",
			2377 => x"025e2545",
			2378 => x"01892545",
			2379 => x"08001d04",
			2380 => x"fe262545",
			2381 => x"ff952545",
			2382 => x"01001204",
			2383 => x"000e2545",
			2384 => x"fe582545",
			2385 => x"04002630",
			2386 => x"0400252c",
			2387 => x"08002328",
			2388 => x"0600af18",
			2389 => x"08001508",
			2390 => x"09001704",
			2391 => x"00a425f9",
			2392 => x"fe8325f9",
			2393 => x"0f00c708",
			2394 => x"01000d04",
			2395 => x"004e25f9",
			2396 => x"ff5a25f9",
			2397 => x"0c001504",
			2398 => x"fed725f9",
			2399 => x"010f25f9",
			2400 => x"01000904",
			2401 => x"008f25f9",
			2402 => x"00014504",
			2403 => x"fe5c25f9",
			2404 => x"05002a04",
			2405 => x"ff7c25f9",
			2406 => x"002725f9",
			2407 => x"fe9825f9",
			2408 => x"018825f9",
			2409 => x"04002b14",
			2410 => x"0b001808",
			2411 => x"05003404",
			2412 => x"ffaa25f9",
			2413 => x"fe7e25f9",
			2414 => x"05003904",
			2415 => x"fec725f9",
			2416 => x"05003a04",
			2417 => x"012c25f9",
			2418 => x"ff7e25f9",
			2419 => x"0f009c04",
			2420 => x"fec125f9",
			2421 => x"0a003d10",
			2422 => x"0500410c",
			2423 => x"00012e04",
			2424 => x"fea625f9",
			2425 => x"04002f04",
			2426 => x"015b25f9",
			2427 => x"ffbe25f9",
			2428 => x"018a25f9",
			2429 => x"feee25f9",
			2430 => x"0001111c",
			2431 => x"04000808",
			2432 => x"06003304",
			2433 => x"fff226a5",
			2434 => x"003726a5",
			2435 => x"06009c0c",
			2436 => x"05004204",
			2437 => x"ff8e26a5",
			2438 => x"05004404",
			2439 => x"001e26a5",
			2440 => x"ffda26a5",
			2441 => x"00010604",
			2442 => x"fff426a5",
			2443 => x"002026a5",
			2444 => x"0e007804",
			2445 => x"007226a5",
			2446 => x"07002b08",
			2447 => x"01000904",
			2448 => x"ff9726a5",
			2449 => x"fffa26a5",
			2450 => x"0d00161c",
			2451 => x"0a003110",
			2452 => x"0b001508",
			2453 => x"00013804",
			2454 => x"ffbc26a5",
			2455 => x"003a26a5",
			2456 => x"00013b04",
			2457 => x"007d26a5",
			2458 => x"001926a5",
			2459 => x"01000804",
			2460 => x"ff9c26a5",
			2461 => x"02011e04",
			2462 => x"ffc126a5",
			2463 => x"003f26a5",
			2464 => x"0a002f04",
			2465 => x"ff7a26a5",
			2466 => x"08002308",
			2467 => x"04002604",
			2468 => x"007d26a5",
			2469 => x"ffcd26a5",
			2470 => x"03003504",
			2471 => x"ffa126a5",
			2472 => x"001626a5",
			2473 => x"03003534",
			2474 => x"09001508",
			2475 => x"00006504",
			2476 => x"febe2711",
			2477 => x"033f2711",
			2478 => x"03002104",
			2479 => x"fe672711",
			2480 => x"08002320",
			2481 => x"0b001710",
			2482 => x"09001e08",
			2483 => x"0c001804",
			2484 => x"000e2711",
			2485 => x"01912711",
			2486 => x"01000c04",
			2487 => x"00342711",
			2488 => x"fdf92711",
			2489 => x"01000908",
			2490 => x"05002b04",
			2491 => x"01572711",
			2492 => x"fddc2711",
			2493 => x"05002c04",
			2494 => x"ff812711",
			2495 => x"01562711",
			2496 => x"07003204",
			2497 => x"00ce2711",
			2498 => x"fe5d2711",
			2499 => x"fe422711",
			2500 => x"0200e914",
			2501 => x"09001504",
			2502 => x"004a27ad",
			2503 => x"0c00170c",
			2504 => x"0b001708",
			2505 => x"0200d104",
			2506 => x"fe5e27ad",
			2507 => x"001027ad",
			2508 => x"015027ad",
			2509 => x"fe5d27ad",
			2510 => x"09002338",
			2511 => x"0e009430",
			2512 => x"02011d18",
			2513 => x"06009f10",
			2514 => x"0a003108",
			2515 => x"0c001504",
			2516 => x"01a627ad",
			2517 => x"03eb27ad",
			2518 => x"04002b04",
			2519 => x"fe3c27ad",
			2520 => x"010727ad",
			2521 => x"07002f04",
			2522 => x"fe3627ad",
			2523 => x"ffd627ad",
			2524 => x"07002b08",
			2525 => x"08001804",
			2526 => x"020b27ad",
			2527 => x"fe3c27ad",
			2528 => x"00013a08",
			2529 => x"03002604",
			2530 => x"013527ad",
			2531 => x"038c27ad",
			2532 => x"0f00c704",
			2533 => x"ff8427ad",
			2534 => x"026327ad",
			2535 => x"0f00cd04",
			2536 => x"005d27ad",
			2537 => x"fe6327ad",
			2538 => x"fe5f27ad",
			2539 => x"04000808",
			2540 => x"06003504",
			2541 => x"fed32859",
			2542 => x"08ea2859",
			2543 => x"0200eb18",
			2544 => x"01000a04",
			2545 => x"fe5c2859",
			2546 => x"0c001710",
			2547 => x"01000b04",
			2548 => x"02af2859",
			2549 => x"08001c08",
			2550 => x"05002304",
			2551 => x"fed02859",
			2552 => x"01812859",
			2553 => x"fe7f2859",
			2554 => x"fe762859",
			2555 => x"09001914",
			2556 => x"0600a208",
			2557 => x"03002304",
			2558 => x"00da2859",
			2559 => x"022d2859",
			2560 => x"0c001508",
			2561 => x"04001804",
			2562 => x"00392859",
			2563 => x"fe3b2859",
			2564 => x"00ff2859",
			2565 => x"08001910",
			2566 => x"07002c08",
			2567 => x"0f00bf04",
			2568 => x"ff722859",
			2569 => x"fde72859",
			2570 => x"05002a04",
			2571 => x"00c12859",
			2572 => x"ff582859",
			2573 => x"01001410",
			2574 => x"00012a08",
			2575 => x"02010f04",
			2576 => x"00c52859",
			2577 => x"fec02859",
			2578 => x"03002604",
			2579 => x"ff8f2859",
			2580 => x"00f22859",
			2581 => x"fe662859",
			2582 => x"04002654",
			2583 => x"05002e3c",
			2584 => x"01000d30",
			2585 => x"04001c1c",
			2586 => x"0c001610",
			2587 => x"0d001208",
			2588 => x"01000804",
			2589 => x"00ad2945",
			2590 => x"ff752945",
			2591 => x"0e007504",
			2592 => x"00932945",
			2593 => x"fefe2945",
			2594 => x"04001a08",
			2595 => x"05002504",
			2596 => x"00892945",
			2597 => x"ff3c2945",
			2598 => x"01302945",
			2599 => x"01000b10",
			2600 => x"04001e08",
			2601 => x"0b001504",
			2602 => x"feca2945",
			2603 => x"000b2945",
			2604 => x"08001904",
			2605 => x"ff942945",
			2606 => x"006d2945",
			2607 => x"008e2945",
			2608 => x"03002704",
			2609 => x"fecd2945",
			2610 => x"0f00bf04",
			2611 => x"ffaa2945",
			2612 => x"005f2945",
			2613 => x"08002314",
			2614 => x"08001c08",
			2615 => x"0f00bc04",
			2616 => x"00a72945",
			2617 => x"fef72945",
			2618 => x"00011304",
			2619 => x"ffcc2945",
			2620 => x"07003304",
			2621 => x"01432945",
			2622 => x"00612945",
			2623 => x"ff2e2945",
			2624 => x"04002b0c",
			2625 => x"05003904",
			2626 => x"ff212945",
			2627 => x"05003a04",
			2628 => x"006a2945",
			2629 => x"ff5d2945",
			2630 => x"00012e0c",
			2631 => x"01000a08",
			2632 => x"01000904",
			2633 => x"ff7f2945",
			2634 => x"00a82945",
			2635 => x"ff2a2945",
			2636 => x"04002f08",
			2637 => x"0600b104",
			2638 => x"00c02945",
			2639 => x"fff62945",
			2640 => x"ffb62945",
			2641 => x"08002358",
			2642 => x"0b001520",
			2643 => x"0600ae14",
			2644 => x"05003110",
			2645 => x"02012f0c",
			2646 => x"0600a708",
			2647 => x"0c001404",
			2648 => x"00a42a09",
			2649 => x"ffbc2a09",
			2650 => x"00f42a09",
			2651 => x"ff102a09",
			2652 => x"fea82a09",
			2653 => x"0600b704",
			2654 => x"fe6b2a09",
			2655 => x"0d001204",
			2656 => x"00ed2a09",
			2657 => x"fed22a09",
			2658 => x"02011e24",
			2659 => x"01000d18",
			2660 => x"01000908",
			2661 => x"09001b04",
			2662 => x"00c02a09",
			2663 => x"fe962a09",
			2664 => x"07002d08",
			2665 => x"0200d104",
			2666 => x"ff262a09",
			2667 => x"01462a09",
			2668 => x"07002f04",
			2669 => x"fea82a09",
			2670 => x"00cf2a09",
			2671 => x"0a003d04",
			2672 => x"fe7d2a09",
			2673 => x"0d001b04",
			2674 => x"009f2a09",
			2675 => x"fff02a09",
			2676 => x"03002704",
			2677 => x"ffde2a09",
			2678 => x"0a003104",
			2679 => x"018f2a09",
			2680 => x"01000c04",
			2681 => x"ff412a09",
			2682 => x"08002004",
			2683 => x"01592a09",
			2684 => x"00882a09",
			2685 => x"0c001c04",
			2686 => x"fe8d2a09",
			2687 => x"0d001b04",
			2688 => x"01182a09",
			2689 => x"ff1d2a09",
			2690 => x"02011c38",
			2691 => x"01000d28",
			2692 => x"0a003118",
			2693 => x"06009f14",
			2694 => x"00010a0c",
			2695 => x"07002908",
			2696 => x"08001804",
			2697 => x"fef82aed",
			2698 => x"00ae2aed",
			2699 => x"feda2aed",
			2700 => x"0a002804",
			2701 => x"00352aed",
			2702 => x"01322aed",
			2703 => x"ff0f2aed",
			2704 => x"09001f04",
			2705 => x"feb32aed",
			2706 => x"08001f04",
			2707 => x"ff6e2aed",
			2708 => x"0200de04",
			2709 => x"fff52aed",
			2710 => x"00f92aed",
			2711 => x"01001f0c",
			2712 => x"0a003d04",
			2713 => x"fea42aed",
			2714 => x"06009604",
			2715 => x"ffeb2aed",
			2716 => x"00602aed",
			2717 => x"00562aed",
			2718 => x"07003730",
			2719 => x"00013a18",
			2720 => x"03002404",
			2721 => x"ffa52aed",
			2722 => x"07002b04",
			2723 => x"ff862aed",
			2724 => x"0600a808",
			2725 => x"05003804",
			2726 => x"011d2aed",
			2727 => x"fff02aed",
			2728 => x"05002904",
			2729 => x"ff2e2aed",
			2730 => x"00842aed",
			2731 => x"0f00d914",
			2732 => x"0600b310",
			2733 => x"0f00c708",
			2734 => x"07002c04",
			2735 => x"00152aed",
			2736 => x"fefa2aed",
			2737 => x"0d001204",
			2738 => x"fefe2aed",
			2739 => x"00a32aed",
			2740 => x"ff2a2aed",
			2741 => x"00e12aed",
			2742 => x"02013904",
			2743 => x"fed22aed",
			2744 => x"00014a04",
			2745 => x"00862aed",
			2746 => x"ffa42aed",
			2747 => x"01000720",
			2748 => x"0e008118",
			2749 => x"0c001408",
			2750 => x"00011104",
			2751 => x"ff7f2bd9",
			2752 => x"00a02bd9",
			2753 => x"0100060c",
			2754 => x"07002808",
			2755 => x"0200af04",
			2756 => x"ffd72bd9",
			2757 => x"004a2bd9",
			2758 => x"feee2bd9",
			2759 => x"003c2bd9",
			2760 => x"05002d04",
			2761 => x"00f12bd9",
			2762 => x"ffc92bd9",
			2763 => x"0600af40",
			2764 => x"01000a1c",
			2765 => x"07002d18",
			2766 => x"05002608",
			2767 => x"0f004b04",
			2768 => x"ffc42bd9",
			2769 => x"00af2bd9",
			2770 => x"08001908",
			2771 => x"07002904",
			2772 => x"00042bd9",
			2773 => x"ff132bd9",
			2774 => x"08001c04",
			2775 => x"00732bd9",
			2776 => x"ff832bd9",
			2777 => x"fedf2bd9",
			2778 => x"00012d18",
			2779 => x"01000d0c",
			2780 => x"04002608",
			2781 => x"0c001604",
			2782 => x"ff972bd9",
			2783 => x"009e2bd9",
			2784 => x"ff602bd9",
			2785 => x"01001d08",
			2786 => x"0e008a04",
			2787 => x"ff012bd9",
			2788 => x"001c2bd9",
			2789 => x"00362bd9",
			2790 => x"01001408",
			2791 => x"05002e04",
			2792 => x"00042bd9",
			2793 => x"00e52bd9",
			2794 => x"ff7c2bd9",
			2795 => x"0a003610",
			2796 => x"0d001204",
			2797 => x"ffd92bd9",
			2798 => x"01001204",
			2799 => x"feed2bd9",
			2800 => x"01001504",
			2801 => x"00062bd9",
			2802 => x"fff32bd9",
			2803 => x"05003804",
			2804 => x"00962bd9",
			2805 => x"ff8f2bd9",
			2806 => x"04002348",
			2807 => x"01000d30",
			2808 => x"03002108",
			2809 => x"09001504",
			2810 => x"002b2cbd",
			2811 => x"ff6e2cbd",
			2812 => x"04001810",
			2813 => x"04001508",
			2814 => x"0e008f04",
			2815 => x"00112cbd",
			2816 => x"ffcc2cbd",
			2817 => x"00010c04",
			2818 => x"ffdf2cbd",
			2819 => x"00bd2cbd",
			2820 => x"04001a08",
			2821 => x"05002604",
			2822 => x"00252cbd",
			2823 => x"ff702cbd",
			2824 => x"01000b08",
			2825 => x"01000704",
			2826 => x"004a2cbd",
			2827 => x"ffcf2cbd",
			2828 => x"06009c04",
			2829 => x"ffdc2cbd",
			2830 => x"00b92cbd",
			2831 => x"05002d08",
			2832 => x"07001f04",
			2833 => x"001b2cbd",
			2834 => x"ff602cbd",
			2835 => x"00013204",
			2836 => x"ffad2cbd",
			2837 => x"00014708",
			2838 => x"0e009004",
			2839 => x"00882cbd",
			2840 => x"fff02cbd",
			2841 => x"ffc82cbd",
			2842 => x"04002508",
			2843 => x"07003204",
			2844 => x"00042cbd",
			2845 => x"ff532cbd",
			2846 => x"04002604",
			2847 => x"00662cbd",
			2848 => x"04002b10",
			2849 => x"0300340c",
			2850 => x"0f00ca04",
			2851 => x"ff762cbd",
			2852 => x"0f00cf04",
			2853 => x"001a2cbd",
			2854 => x"ffcf2cbd",
			2855 => x"00042cbd",
			2856 => x"0400320c",
			2857 => x"0c001804",
			2858 => x"ffdb2cbd",
			2859 => x"0200ef04",
			2860 => x"ffed2cbd",
			2861 => x"00592cbd",
			2862 => x"ffbf2cbd",
			2863 => x"0900191c",
			2864 => x"0f00c314",
			2865 => x"0001190c",
			2866 => x"0a002508",
			2867 => x"04000804",
			2868 => x"002e2db1",
			2869 => x"ff742db1",
			2870 => x"003b2db1",
			2871 => x"04001f04",
			2872 => x"00c92db1",
			2873 => x"00212db1",
			2874 => x"0c001404",
			2875 => x"ff712db1",
			2876 => x"003f2db1",
			2877 => x"00013130",
			2878 => x"02010f24",
			2879 => x"0f00b21c",
			2880 => x"0e006f0c",
			2881 => x"0f008b08",
			2882 => x"00008604",
			2883 => x"00022db1",
			2884 => x"ff8b2db1",
			2885 => x"006c2db1",
			2886 => x"04002208",
			2887 => x"04001804",
			2888 => x"000e2db1",
			2889 => x"ff492db1",
			2890 => x"0e007504",
			2891 => x"ffc02db1",
			2892 => x"00402db1",
			2893 => x"00010e04",
			2894 => x"ffe52db1",
			2895 => x"00ab2db1",
			2896 => x"0b001804",
			2897 => x"ff392db1",
			2898 => x"0f00bc04",
			2899 => x"00432db1",
			2900 => x"fff42db1",
			2901 => x"0600a90c",
			2902 => x"08001904",
			2903 => x"ffc02db1",
			2904 => x"05003704",
			2905 => x"00b32db1",
			2906 => x"ffeb2db1",
			2907 => x"03002708",
			2908 => x"07003004",
			2909 => x"00082db1",
			2910 => x"ff452db1",
			2911 => x"03002d0c",
			2912 => x"0b001904",
			2913 => x"009b2db1",
			2914 => x"05003404",
			2915 => x"ffb02db1",
			2916 => x"00072db1",
			2917 => x"00013708",
			2918 => x"0a003804",
			2919 => x"004c2db1",
			2920 => x"fffa2db1",
			2921 => x"02013204",
			2922 => x"ff632db1",
			2923 => x"fffb2db1",
			2924 => x"0e009348",
			2925 => x"00014a44",
			2926 => x"0600a830",
			2927 => x"0e00851c",
			2928 => x"0900190c",
			2929 => x"06004404",
			2930 => x"ff372e65",
			2931 => x"04002004",
			2932 => x"00ab2e65",
			2933 => x"ff6d2e65",
			2934 => x"03002408",
			2935 => x"0d001104",
			2936 => x"001e2e65",
			2937 => x"fed02e65",
			2938 => x"01000604",
			2939 => x"fecf2e65",
			2940 => x"00272e65",
			2941 => x"0f00bb0c",
			2942 => x"07003704",
			2943 => x"ff092e65",
			2944 => x"0a003904",
			2945 => x"00c82e65",
			2946 => x"fffa2e65",
			2947 => x"05003904",
			2948 => x"01472e65",
			2949 => x"000c2e65",
			2950 => x"02012804",
			2951 => x"feb72e65",
			2952 => x"09001a04",
			2953 => x"ff0c2e65",
			2954 => x"0f00c704",
			2955 => x"ff562e65",
			2956 => x"00014204",
			2957 => x"00e22e65",
			2958 => x"ffee2e65",
			2959 => x"00df2e65",
			2960 => x"0c001a08",
			2961 => x"05002204",
			2962 => x"00452e65",
			2963 => x"feb52e65",
			2964 => x"04002608",
			2965 => x"02013904",
			2966 => x"ffd22e65",
			2967 => x"00e12e65",
			2968 => x"ff4a2e65",
			2969 => x"0600af50",
			2970 => x"0f00c640",
			2971 => x"0f00c02c",
			2972 => x"02012020",
			2973 => x"01000d10",
			2974 => x"0a003108",
			2975 => x"0f004b04",
			2976 => x"fee42f41",
			2977 => x"00842f41",
			2978 => x"05004204",
			2979 => x"febb2f41",
			2980 => x"00552f41",
			2981 => x"03003408",
			2982 => x"01001a04",
			2983 => x"fe872f41",
			2984 => x"006c2f41",
			2985 => x"05003e04",
			2986 => x"00c32f41",
			2987 => x"ff702f41",
			2988 => x"01000904",
			2989 => x"00482f41",
			2990 => x"0d001a04",
			2991 => x"017e2f41",
			2992 => x"ff812f41",
			2993 => x"0d001104",
			2994 => x"00792f41",
			2995 => x"01000a04",
			2996 => x"fe6f2f41",
			2997 => x"02012b08",
			2998 => x"04002704",
			2999 => x"fefa2f41",
			3000 => x"003e2f41",
			3001 => x"01072f41",
			3002 => x"0c001504",
			3003 => x"fef12f41",
			3004 => x"09001f08",
			3005 => x"0d001304",
			3006 => x"00a82f41",
			3007 => x"015e2f41",
			3008 => x"ffdd2f41",
			3009 => x"01000904",
			3010 => x"00802f41",
			3011 => x"0c001808",
			3012 => x"0f00df04",
			3013 => x"fe962f41",
			3014 => x"00392f41",
			3015 => x"0a003208",
			3016 => x"00014504",
			3017 => x"ffa82f41",
			3018 => x"00e22f41",
			3019 => x"03003304",
			3020 => x"feb42f41",
			3021 => x"03003404",
			3022 => x"00e92f41",
			3023 => x"ffb22f41",
			3024 => x"0000f324",
			3025 => x"0400080c",
			3026 => x"04000704",
			3027 => x"ffdf3035",
			3028 => x"06002404",
			3029 => x"fffb3035",
			3030 => x"005f3035",
			3031 => x"09001f08",
			3032 => x"0d001704",
			3033 => x"ff0c3035",
			3034 => x"00113035",
			3035 => x"0d00150c",
			3036 => x"09002008",
			3037 => x"0b001704",
			3038 => x"fff83035",
			3039 => x"00533035",
			3040 => x"ffea3035",
			3041 => x"ffbe3035",
			3042 => x"0600a938",
			3043 => x"07002b10",
			3044 => x"06009404",
			3045 => x"008a3035",
			3046 => x"0c001408",
			3047 => x"01000704",
			3048 => x"00693035",
			3049 => x"ff933035",
			3050 => x"ff0c3035",
			3051 => x"08001f10",
			3052 => x"04002004",
			3053 => x"00ff3035",
			3054 => x"02012b08",
			3055 => x"00011804",
			3056 => x"00573035",
			3057 => x"ff8b3035",
			3058 => x"00643035",
			3059 => x"0e00830c",
			3060 => x"0e007e08",
			3061 => x"0e007804",
			3062 => x"fff43035",
			3063 => x"000e3035",
			3064 => x"ff4f3035",
			3065 => x"0600a204",
			3066 => x"ffcd3035",
			3067 => x"04002c04",
			3068 => x"00a63035",
			3069 => x"ffce3035",
			3070 => x"02012804",
			3071 => x"ff263035",
			3072 => x"07002c04",
			3073 => x"ff503035",
			3074 => x"0700340c",
			3075 => x"03002d08",
			3076 => x"01000904",
			3077 => x"00e43035",
			3078 => x"00213035",
			3079 => x"ffd93035",
			3080 => x"00013704",
			3081 => x"00733035",
			3082 => x"03003104",
			3083 => x"ff2b3035",
			3084 => x"ffe43035",
			3085 => x"03002108",
			3086 => x"0d000e04",
			3087 => x"fffb30f1",
			3088 => x"ff9230f1",
			3089 => x"05002614",
			3090 => x"07002f10",
			3091 => x"0c001508",
			3092 => x"05002404",
			3093 => x"ffd330f1",
			3094 => x"001030f1",
			3095 => x"0000cc04",
			3096 => x"fff530f1",
			3097 => x"00ad30f1",
			3098 => x"ffb530f1",
			3099 => x"0f00c72c",
			3100 => x"01000914",
			3101 => x"01000304",
			3102 => x"003430f1",
			3103 => x"0d001508",
			3104 => x"0c001404",
			3105 => x"fff130f1",
			3106 => x"ff4330f1",
			3107 => x"0c001a04",
			3108 => x"002b30f1",
			3109 => x"fffb30f1",
			3110 => x"0d001308",
			3111 => x"0000d104",
			3112 => x"fff230f1",
			3113 => x"006c30f1",
			3114 => x"05003608",
			3115 => x"08001d04",
			3116 => x"000830f1",
			3117 => x"ff9330f1",
			3118 => x"04002604",
			3119 => x"004e30f1",
			3120 => x"ffd830f1",
			3121 => x"0700340c",
			3122 => x"09001c08",
			3123 => x"0f00ca04",
			3124 => x"002e30f1",
			3125 => x"ffbb30f1",
			3126 => x"008630f1",
			3127 => x"0a003604",
			3128 => x"ff9a30f1",
			3129 => x"05003804",
			3130 => x"004130f1",
			3131 => x"ffe030f1",
			3132 => x"0f00c044",
			3133 => x"02012038",
			3134 => x"0a002f20",
			3135 => x"0000f314",
			3136 => x"04000808",
			3137 => x"04000704",
			3138 => x"fff731fd",
			3139 => x"002e31fd",
			3140 => x"0c001604",
			3141 => x"ff9731fd",
			3142 => x"0c001704",
			3143 => x"002e31fd",
			3144 => x"ffda31fd",
			3145 => x"0f00b508",
			3146 => x"0c001504",
			3147 => x"001331fd",
			3148 => x"008d31fd",
			3149 => x"ffe731fd",
			3150 => x"02011d14",
			3151 => x"05004208",
			3152 => x"07003704",
			3153 => x"ff6931fd",
			3154 => x"001331fd",
			3155 => x"05004708",
			3156 => x"01000a04",
			3157 => x"003431fd",
			3158 => x"fff531fd",
			3159 => x"ffdc31fd",
			3160 => x"001131fd",
			3161 => x"0d001a08",
			3162 => x"01000a04",
			3163 => x"001931fd",
			3164 => x"00a131fd",
			3165 => x"ffde31fd",
			3166 => x"0f00c610",
			3167 => x"0a002a04",
			3168 => x"002931fd",
			3169 => x"04002504",
			3170 => x"ff5e31fd",
			3171 => x"05003b04",
			3172 => x"001531fd",
			3173 => x"ffea31fd",
			3174 => x"0600ae0c",
			3175 => x"0c001504",
			3176 => x"ffca31fd",
			3177 => x"0b001604",
			3178 => x"007e31fd",
			3179 => x"fffd31fd",
			3180 => x"09001d14",
			3181 => x"0f00de0c",
			3182 => x"03002d08",
			3183 => x"04001704",
			3184 => x"fffe31fd",
			3185 => x"ff6c31fd",
			3186 => x"000c31fd",
			3187 => x"0f00e404",
			3188 => x"002d31fd",
			3189 => x"ffed31fd",
			3190 => x"04002308",
			3191 => x"0c001b04",
			3192 => x"009431fd",
			3193 => x"ffcc31fd",
			3194 => x"0a003604",
			3195 => x"ff9531fd",
			3196 => x"0a003704",
			3197 => x"003531fd",
			3198 => x"ffd931fd",
			3199 => x"0400262c",
			3200 => x"04002528",
			3201 => x"08002324",
			3202 => x"07003620",
			3203 => x"05002f10",
			3204 => x"0d001808",
			3205 => x"04002004",
			3206 => x"002f32a9",
			3207 => x"ff8032a9",
			3208 => x"0a002d04",
			3209 => x"fe8132a9",
			3210 => x"008e32a9",
			3211 => x"05003208",
			3212 => x"0e008304",
			3213 => x"013932a9",
			3214 => x"006532a9",
			3215 => x"07002e04",
			3216 => x"fedd32a9",
			3217 => x"006f32a9",
			3218 => x"febe32a9",
			3219 => x"feb632a9",
			3220 => x"016032a9",
			3221 => x"04002804",
			3222 => x"fe9e32a9",
			3223 => x"08001d10",
			3224 => x"0700320c",
			3225 => x"0c001904",
			3226 => x"fea432a9",
			3227 => x"05004704",
			3228 => x"00ab32a9",
			3229 => x"ff7532a9",
			3230 => x"00b032a9",
			3231 => x"0e008c14",
			3232 => x"0d001608",
			3233 => x"0a003d04",
			3234 => x"016132a9",
			3235 => x"ff7c32a9",
			3236 => x"03003404",
			3237 => x"fed332a9",
			3238 => x"05004004",
			3239 => x"012432a9",
			3240 => x"ff7432a9",
			3241 => x"fefd32a9",
			3242 => x"0700365c",
			3243 => x"0b001724",
			3244 => x"08001f20",
			3245 => x"0b001208",
			3246 => x"0c001004",
			3247 => x"00193375",
			3248 => x"ff2f3375",
			3249 => x"0e008a0c",
			3250 => x"0600ab08",
			3251 => x"05002c04",
			3252 => x"00553375",
			3253 => x"ff8b3375",
			3254 => x"ff533375",
			3255 => x"01000904",
			3256 => x"00d93375",
			3257 => x"04001604",
			3258 => x"00623375",
			3259 => x"ff823375",
			3260 => x"ff223375",
			3261 => x"01000910",
			3262 => x"05002b0c",
			3263 => x"0d001304",
			3264 => x"ffb93375",
			3265 => x"01000604",
			3266 => x"00813375",
			3267 => x"fffa3375",
			3268 => x"ff333375",
			3269 => x"05002c0c",
			3270 => x"08001c08",
			3271 => x"03001d04",
			3272 => x"fffa3375",
			3273 => x"00673375",
			3274 => x"ff683375",
			3275 => x"0900210c",
			3276 => x"00012a08",
			3277 => x"09001f04",
			3278 => x"ffa43375",
			3279 => x"006c3375",
			3280 => x"00fb3375",
			3281 => x"0b001b08",
			3282 => x"0d001804",
			3283 => x"fffe3375",
			3284 => x"ff7e3375",
			3285 => x"0c001d04",
			3286 => x"00583375",
			3287 => x"fff73375",
			3288 => x"0e008b08",
			3289 => x"0d001b04",
			3290 => x"003a3375",
			3291 => x"fff13375",
			3292 => x"ff1a3375",
			3293 => x"07003378",
			3294 => x"0b001540",
			3295 => x"09001920",
			3296 => x"0b001418",
			3297 => x"06009d0c",
			3298 => x"06004404",
			3299 => x"ffac34a1",
			3300 => x"00011004",
			3301 => x"001834a1",
			3302 => x"00b034a1",
			3303 => x"07002d08",
			3304 => x"03002404",
			3305 => x"ffe634a1",
			3306 => x"ff3e34a1",
			3307 => x"002834a1",
			3308 => x"0e008304",
			3309 => x"00c034a1",
			3310 => x"000434a1",
			3311 => x"02012b14",
			3312 => x"07002e0c",
			3313 => x"0e007508",
			3314 => x"06007b04",
			3315 => x"ffa034a1",
			3316 => x"003234a1",
			3317 => x"ff1e34a1",
			3318 => x"04001a04",
			3319 => x"ffd634a1",
			3320 => x"006434a1",
			3321 => x"01000a08",
			3322 => x"03002904",
			3323 => x"009434a1",
			3324 => x"000234a1",
			3325 => x"ffb634a1",
			3326 => x"0a00311c",
			3327 => x"01000d14",
			3328 => x"0a00280c",
			3329 => x"0d001204",
			3330 => x"007734a1",
			3331 => x"05002404",
			3332 => x"003934a1",
			3333 => x"ff5f34a1",
			3334 => x"0b001904",
			3335 => x"00f634a1",
			3336 => x"ffca34a1",
			3337 => x"05002c04",
			3338 => x"ff3a34a1",
			3339 => x"005934a1",
			3340 => x"08001d0c",
			3341 => x"04002e04",
			3342 => x"ff3d34a1",
			3343 => x"05004704",
			3344 => x"003a34a1",
			3345 => x"ffd634a1",
			3346 => x"0f00ba0c",
			3347 => x"01000b04",
			3348 => x"005434a1",
			3349 => x"03003404",
			3350 => x"ff7434a1",
			3351 => x"001034a1",
			3352 => x"00a334a1",
			3353 => x"0a003608",
			3354 => x"04002804",
			3355 => x"ff2b34a1",
			3356 => x"ffe234a1",
			3357 => x"0001370c",
			3358 => x"05003a04",
			3359 => x"00bc34a1",
			3360 => x"0e008d04",
			3361 => x"ffb534a1",
			3362 => x"000134a1",
			3363 => x"02013904",
			3364 => x"ff8034a1",
			3365 => x"02013e04",
			3366 => x"004f34a1",
			3367 => x"fff134a1",
			3368 => x"0b001208",
			3369 => x"0c001004",
			3370 => x"ffc83555",
			3371 => x"fe963555",
			3372 => x"04001618",
			3373 => x"01000504",
			3374 => x"feeb3555",
			3375 => x"0c001710",
			3376 => x"0e00960c",
			3377 => x"06004404",
			3378 => x"ffcf3555",
			3379 => x"01000a04",
			3380 => x"018b3555",
			3381 => x"00b33555",
			3382 => x"ff893555",
			3383 => x"ff083555",
			3384 => x"0a003b34",
			3385 => x"0600b11c",
			3386 => x"0f00c710",
			3387 => x"0600a808",
			3388 => x"03002404",
			3389 => x"ff533555",
			3390 => x"004b3555",
			3391 => x"05003604",
			3392 => x"fe513555",
			3393 => x"ffc23555",
			3394 => x"0c001504",
			3395 => x"fe553555",
			3396 => x"00014204",
			3397 => x"01473555",
			3398 => x"00393555",
			3399 => x"0f00d90c",
			3400 => x"0e009504",
			3401 => x"fe613555",
			3402 => x"02013904",
			3403 => x"fec73555",
			3404 => x"00f93555",
			3405 => x"00015808",
			3406 => x"0600c304",
			3407 => x"01783555",
			3408 => x"ff663555",
			3409 => x"ff153555",
			3410 => x"05003d04",
			3411 => x"fff93555",
			3412 => x"fe893555",
			3413 => x"0c00185c",
			3414 => x"0c00174c",
			3415 => x"0b001530",
			3416 => x"08001818",
			3417 => x"00011108",
			3418 => x"09001a04",
			3419 => x"ff553679",
			3420 => x"00263679",
			3421 => x"09001908",
			3422 => x"0c001404",
			3423 => x"00d33679",
			3424 => x"00183679",
			3425 => x"05002c04",
			3426 => x"fff03679",
			3427 => x"ff873679",
			3428 => x"09001c10",
			3429 => x"0e007808",
			3430 => x"0d001104",
			3431 => x"004b3679",
			3432 => x"ffe93679",
			3433 => x"00015204",
			3434 => x"ff403679",
			3435 => x"00173679",
			3436 => x"07002d04",
			3437 => x"ffaa3679",
			3438 => x"00743679",
			3439 => x"0a002f10",
			3440 => x"0d00150c",
			3441 => x"01000704",
			3442 => x"ffed3679",
			3443 => x"03002104",
			3444 => x"fff63679",
			3445 => x"00f13679",
			3446 => x"ffa03679",
			3447 => x"03002f04",
			3448 => x"ff6a3679",
			3449 => x"09001d04",
			3450 => x"ffe13679",
			3451 => x"00243679",
			3452 => x"01000604",
			3453 => x"00213679",
			3454 => x"05002d04",
			3455 => x"ff043679",
			3456 => x"03002f04",
			3457 => x"003d3679",
			3458 => x"ff7e3679",
			3459 => x"0b001a2c",
			3460 => x"08001c18",
			3461 => x"0100060c",
			3462 => x"0d001304",
			3463 => x"ffc73679",
			3464 => x"05002d04",
			3465 => x"008a3679",
			3466 => x"fff63679",
			3467 => x"05004604",
			3468 => x"ff593679",
			3469 => x"07002c04",
			3470 => x"ffe93679",
			3471 => x"002e3679",
			3472 => x"05002c04",
			3473 => x"ffa43679",
			3474 => x"0100140c",
			3475 => x"00012d08",
			3476 => x"05003804",
			3477 => x"ffca3679",
			3478 => x"00623679",
			3479 => x"00e93679",
			3480 => x"ffb13679",
			3481 => x"03003504",
			3482 => x"ff543679",
			3483 => x"0a003b04",
			3484 => x"00453679",
			3485 => x"ffe93679",
			3486 => x"0600a840",
			3487 => x"00013a3c",
			3488 => x"00013134",
			3489 => x"09001914",
			3490 => x"0b001208",
			3491 => x"0c001104",
			3492 => x"00033755",
			3493 => x"ffb83755",
			3494 => x"08001504",
			3495 => x"ffeb3755",
			3496 => x"0a002504",
			3497 => x"00073755",
			3498 => x"008b3755",
			3499 => x"01000910",
			3500 => x"08001d08",
			3501 => x"0a002404",
			3502 => x"000e3755",
			3503 => x"ff683755",
			3504 => x"07002e04",
			3505 => x"fff93755",
			3506 => x"001f3755",
			3507 => x"01000d08",
			3508 => x"0c001504",
			3509 => x"ffc33755",
			3510 => x"00583755",
			3511 => x"00012904",
			3512 => x"ff7b3755",
			3513 => x"00253755",
			3514 => x"08001f04",
			3515 => x"00903755",
			3516 => x"00193755",
			3517 => x"ff9b3755",
			3518 => x"0f00c708",
			3519 => x"0a002f04",
			3520 => x"000e3755",
			3521 => x"ff513755",
			3522 => x"0600ae08",
			3523 => x"0d001304",
			3524 => x"ffea3755",
			3525 => x"00953755",
			3526 => x"02013810",
			3527 => x"0c001804",
			3528 => x"ff4f3755",
			3529 => x"03002f08",
			3530 => x"0f00cf04",
			3531 => x"003e3755",
			3532 => x"fffa3755",
			3533 => x"ffd23755",
			3534 => x"05002804",
			3535 => x"00543755",
			3536 => x"0f00d304",
			3537 => x"00393755",
			3538 => x"0f00db04",
			3539 => x"ff7c3755",
			3540 => x"00113755",
			3541 => x"0f008b04",
			3542 => x"fe6737e1",
			3543 => x"07003840",
			3544 => x"0d001218",
			3545 => x"04002214",
			3546 => x"01000504",
			3547 => x"020437e1",
			3548 => x"0b001308",
			3549 => x"0600a004",
			3550 => x"013b37e1",
			3551 => x"fe6c37e1",
			3552 => x"03002304",
			3553 => x"ff3d37e1",
			3554 => x"019d37e1",
			3555 => x"fe7137e1",
			3556 => x"0c001508",
			3557 => x"05002704",
			3558 => x"fe1937e1",
			3559 => x"ffa637e1",
			3560 => x"01000810",
			3561 => x"05002b08",
			3562 => x"00011304",
			3563 => x"fedd37e1",
			3564 => x"00fc37e1",
			3565 => x"09001d04",
			3566 => x"fe6137e1",
			3567 => x"fdb637e1",
			3568 => x"01000d08",
			3569 => x"03003104",
			3570 => x"013137e1",
			3571 => x"ff9c37e1",
			3572 => x"05002c04",
			3573 => x"fdcd37e1",
			3574 => x"009537e1",
			3575 => x"fe6d37e1",
			3576 => x"0f008b04",
			3577 => x"fe66387f",
			3578 => x"07003848",
			3579 => x"0d001218",
			3580 => x"04002214",
			3581 => x"0f00bc08",
			3582 => x"03002104",
			3583 => x"0093387f",
			3584 => x"025b387f",
			3585 => x"0e008b08",
			3586 => x"0600a804",
			3587 => x"0088387f",
			3588 => x"fecd387f",
			3589 => x"027c387f",
			3590 => x"fe6b387f",
			3591 => x"01000810",
			3592 => x"05002b08",
			3593 => x"0600a704",
			3594 => x"ff38387f",
			3595 => x"018d387f",
			3596 => x"09001d04",
			3597 => x"fe56387f",
			3598 => x"fd94387f",
			3599 => x"05002c10",
			3600 => x"08001d08",
			3601 => x"0600ab04",
			3602 => x"013f387f",
			3603 => x"fed6387f",
			3604 => x"05002904",
			3605 => x"fe37387f",
			3606 => x"fcc7387f",
			3607 => x"00012d08",
			3608 => x"01000b04",
			3609 => x"00fa387f",
			3610 => x"feff387f",
			3611 => x"0d001a04",
			3612 => x"01b6387f",
			3613 => x"ff65387f",
			3614 => x"fe69387f",
			3615 => x"0f008b10",
			3616 => x"09001504",
			3617 => x"011a38d9",
			3618 => x"0c001708",
			3619 => x"09001e04",
			3620 => x"fe6b38d9",
			3621 => x"019138d9",
			3622 => x"fe6638d9",
			3623 => x"0900231c",
			3624 => x"0e006f04",
			3625 => x"020c38d9",
			3626 => x"03002108",
			3627 => x"00012204",
			3628 => x"fe4d38d9",
			3629 => x"ff6038d9",
			3630 => x"0f00a004",
			3631 => x"fe5638d9",
			3632 => x"0e009708",
			3633 => x"05002404",
			3634 => x"021a38d9",
			3635 => x"00cf38d9",
			3636 => x"fe7a38d9",
			3637 => x"fe6a38d9",
			3638 => x"03001008",
			3639 => x"06002d04",
			3640 => x"ff183945",
			3641 => x"04203945",
			3642 => x"05003a20",
			3643 => x"08001508",
			3644 => x"07002104",
			3645 => x"000c3945",
			3646 => x"fe563945",
			3647 => x"01000204",
			3648 => x"01a33945",
			3649 => x"08002410",
			3650 => x"05003608",
			3651 => x"08002004",
			3652 => x"00213945",
			3653 => x"ff513945",
			3654 => x"0b001704",
			3655 => x"fed83945",
			3656 => x"01a03945",
			3657 => x"fe903945",
			3658 => x"0b001708",
			3659 => x"0d001404",
			3660 => x"fec63945",
			3661 => x"01033945",
			3662 => x"04002704",
			3663 => x"004b3945",
			3664 => x"fe563945",
			3665 => x"09002038",
			3666 => x"0000f318",
			3667 => x"04000808",
			3668 => x"05000f04",
			3669 => x"feb239c9",
			3670 => x"07ca39c9",
			3671 => x"01000a04",
			3672 => x"fe5b39c9",
			3673 => x"0c001604",
			3674 => x"fe7239c9",
			3675 => x"0c001704",
			3676 => x"027139c9",
			3677 => x"fe7e39c9",
			3678 => x"0e00961c",
			3679 => x"00014514",
			3680 => x"0600ae10",
			3681 => x"05002708",
			3682 => x"0a002104",
			3683 => x"ff8d39c9",
			3684 => x"019839c9",
			3685 => x"01000904",
			3686 => x"ffed39c9",
			3687 => x"00c439c9",
			3688 => x"ff1639c9",
			3689 => x"0b001504",
			3690 => x"007439c9",
			3691 => x"01f839c9",
			3692 => x"fe6d39c9",
			3693 => x"0600a304",
			3694 => x"fe6439c9",
			3695 => x"01001204",
			3696 => x"00a839c9",
			3697 => x"fe5539c9",
			3698 => x"0200ef10",
			3699 => x"0c00170c",
			3700 => x"0c001604",
			3701 => x"fe4f3a35",
			3702 => x"01000a04",
			3703 => x"fe893a35",
			3704 => x"02133a35",
			3705 => x"fe693a35",
			3706 => x"09002324",
			3707 => x"09001704",
			3708 => x"019e3a35",
			3709 => x"03002104",
			3710 => x"fe5e3a35",
			3711 => x"07002b10",
			3712 => x"0600a008",
			3713 => x"09001904",
			3714 => x"017f3a35",
			3715 => x"ff6e3a35",
			3716 => x"0c001404",
			3717 => x"fec83a35",
			3718 => x"fe123a35",
			3719 => x"01000404",
			3720 => x"02513a35",
			3721 => x"00012a04",
			3722 => x"ffde3a35",
			3723 => x"00ab3a35",
			3724 => x"fe753a35",
			3725 => x"0f008b10",
			3726 => x"09001504",
			3727 => x"00133aa9",
			3728 => x"0c001708",
			3729 => x"0b001704",
			3730 => x"fe633aa9",
			3731 => x"01293aa9",
			3732 => x"fe603aa9",
			3733 => x"09002328",
			3734 => x"0e009724",
			3735 => x"0200eb08",
			3736 => x"0f008e04",
			3737 => x"02c03aa9",
			3738 => x"fe5d3aa9",
			3739 => x"0c001810",
			3740 => x"0a003208",
			3741 => x"01000d04",
			3742 => x"01993aa9",
			3743 => x"fffd3aa9",
			3744 => x"01000a04",
			3745 => x"fe513aa9",
			3746 => x"00233aa9",
			3747 => x"08002308",
			3748 => x"03002c04",
			3749 => x"01353aa9",
			3750 => x"029c3aa9",
			3751 => x"002f3aa9",
			3752 => x"fe6f3aa9",
			3753 => x"fe623aa9",
			3754 => x"04002644",
			3755 => x"05002e2c",
			3756 => x"01000d20",
			3757 => x"05002b14",
			3758 => x"07003310",
			3759 => x"0b001508",
			3760 => x"04001e04",
			3761 => x"ffdd3b7d",
			3762 => x"00813b7d",
			3763 => x"0a002804",
			3764 => x"fffe3b7d",
			3765 => x"013a3b7d",
			3766 => x"ff373b7d",
			3767 => x"0e008308",
			3768 => x"00012b04",
			3769 => x"fff63b7d",
			3770 => x"fed23b7d",
			3771 => x"00463b7d",
			3772 => x"03002704",
			3773 => x"fec23b7d",
			3774 => x"0f00bf04",
			3775 => x"ffa73b7d",
			3776 => x"00643b7d",
			3777 => x"08002314",
			3778 => x"08001c08",
			3779 => x"0f00bc04",
			3780 => x"00b93b7d",
			3781 => x"feec3b7d",
			3782 => x"00011304",
			3783 => x"ffca3b7d",
			3784 => x"07003304",
			3785 => x"014e3b7d",
			3786 => x"006e3b7d",
			3787 => x"ff293b7d",
			3788 => x"0c001914",
			3789 => x"04002e08",
			3790 => x"0a003604",
			3791 => x"ffb33b7d",
			3792 => x"fed53b7d",
			3793 => x"07002a04",
			3794 => x"ff9a3b7d",
			3795 => x"01000604",
			3796 => x"fff33b7d",
			3797 => x"00a53b7d",
			3798 => x"09002108",
			3799 => x"07002c04",
			3800 => x"ffc23b7d",
			3801 => x"00ad3b7d",
			3802 => x"0d001608",
			3803 => x"0c001c04",
			3804 => x"ffbf3b7d",
			3805 => x"00393b7d",
			3806 => x"ff233b7d",
			3807 => x"0200e914",
			3808 => x"09001504",
			3809 => x"003d3c09",
			3810 => x"0c00170c",
			3811 => x"0b001708",
			3812 => x"0200d104",
			3813 => x"fe5c3c09",
			3814 => x"00093c09",
			3815 => x"01713c09",
			3816 => x"fe5b3c09",
			3817 => x"0900222c",
			3818 => x"0e009428",
			3819 => x"0c001514",
			3820 => x"0600a50c",
			3821 => x"00011904",
			3822 => x"fedd3c09",
			3823 => x"0a002c04",
			3824 => x"04e43c09",
			3825 => x"01f93c09",
			3826 => x"0e008d04",
			3827 => x"fe333c09",
			3828 => x"006f3c09",
			3829 => x"05002504",
			3830 => x"046c3c09",
			3831 => x"08001908",
			3832 => x"0f00c604",
			3833 => x"ff513c09",
			3834 => x"02ff3c09",
			3835 => x"01000d04",
			3836 => x"03653c09",
			3837 => x"01ea3c09",
			3838 => x"fe573c09",
			3839 => x"0d001804",
			3840 => x"00f13c09",
			3841 => x"fe5c3c09",
			3842 => x"0200e914",
			3843 => x"04000808",
			3844 => x"04000704",
			3845 => x"ffe43c9d",
			3846 => x"004a3c9d",
			3847 => x"05003604",
			3848 => x"ff273c9d",
			3849 => x"00008904",
			3850 => x"00323c9d",
			3851 => x"ffbd3c9d",
			3852 => x"01001130",
			3853 => x"03002104",
			3854 => x"ff863c9d",
			3855 => x"0600af1c",
			3856 => x"0b001810",
			3857 => x"0a002f08",
			3858 => x"0600a004",
			3859 => x"008c3c9d",
			3860 => x"00153c9d",
			3861 => x"02011d04",
			3862 => x"ff703c9d",
			3863 => x"00243c9d",
			3864 => x"0e008208",
			3865 => x"08002004",
			3866 => x"00223c9d",
			3867 => x"ffcf3c9d",
			3868 => x"00ca3c9d",
			3869 => x"01000904",
			3870 => x"005b3c9d",
			3871 => x"02013704",
			3872 => x"ff303c9d",
			3873 => x"0f00d504",
			3874 => x"002d3c9d",
			3875 => x"ffb13c9d",
			3876 => x"01002104",
			3877 => x"ff433c9d",
			3878 => x"002a3c9d",
			3879 => x"0900204c",
			3880 => x"0c001828",
			3881 => x"0d001824",
			3882 => x"0600ae18",
			3883 => x"0a003410",
			3884 => x"0e008908",
			3885 => x"08001f04",
			3886 => x"00383d79",
			3887 => x"ff033d79",
			3888 => x"0e008d04",
			3889 => x"01383d79",
			3890 => x"ff993d79",
			3891 => x"0b001604",
			3892 => x"fecf3d79",
			3893 => x"ffee3d79",
			3894 => x"02013c08",
			3895 => x"02013404",
			3896 => x"fe883d79",
			3897 => x"ff8c3d79",
			3898 => x"00a33d79",
			3899 => x"fe913d79",
			3900 => x"08001d18",
			3901 => x"04001e08",
			3902 => x"04001a04",
			3903 => x"ff3d3d79",
			3904 => x"015b3d79",
			3905 => x"04002e08",
			3906 => x"05003504",
			3907 => x"ff783d79",
			3908 => x"fea13d79",
			3909 => x"04003504",
			3910 => x"00e23d79",
			3911 => x"ffb03d79",
			3912 => x"05002d04",
			3913 => x"ff0b3d79",
			3914 => x"04002804",
			3915 => x"01613d79",
			3916 => x"00593d79",
			3917 => x"03003110",
			3918 => x"0700320c",
			3919 => x"04001b08",
			3920 => x"04001a04",
			3921 => x"ff9f3d79",
			3922 => x"00a23d79",
			3923 => x"ff653d79",
			3924 => x"fe9c3d79",
			3925 => x"05003808",
			3926 => x"05003604",
			3927 => x"ffca3d79",
			3928 => x"01123d79",
			3929 => x"08002404",
			3930 => x"fee83d79",
			3931 => x"01001104",
			3932 => x"007e3d79",
			3933 => x"ffa93d79",
			3934 => x"0900203c",
			3935 => x"0e009638",
			3936 => x"0c00181c",
			3937 => x"0d001818",
			3938 => x"0600ae10",
			3939 => x"0a002f08",
			3940 => x"05002e04",
			3941 => x"002a3e25",
			3942 => x"01333e25",
			3943 => x"00012904",
			3944 => x"fe913e25",
			3945 => x"00423e25",
			3946 => x"00014104",
			3947 => x"fe943e25",
			3948 => x"00203e25",
			3949 => x"fe9e3e25",
			3950 => x"0e008114",
			3951 => x"01000b0c",
			3952 => x"08001d08",
			3953 => x"05004604",
			3954 => x"ff0b3e25",
			3955 => x"006c3e25",
			3956 => x"013b3e25",
			3957 => x"0c001a04",
			3958 => x"fec03e25",
			3959 => x"ffe43e25",
			3960 => x"01000c04",
			3961 => x"00173e25",
			3962 => x"017e3e25",
			3963 => x"fedc3e25",
			3964 => x"03003110",
			3965 => x"0700320c",
			3966 => x"04001b08",
			3967 => x"04001a04",
			3968 => x"ffa53e25",
			3969 => x"00953e25",
			3970 => x"ff6c3e25",
			3971 => x"fea33e25",
			3972 => x"0d001a08",
			3973 => x"00012e04",
			3974 => x"ff0f3e25",
			3975 => x"00d23e25",
			3976 => x"feef3e25",
			3977 => x"03001008",
			3978 => x"0e002b04",
			3979 => x"ff283eb9",
			3980 => x"03463eb9",
			3981 => x"0200e914",
			3982 => x"01000a04",
			3983 => x"fe773eb9",
			3984 => x"0c00170c",
			3985 => x"03002c08",
			3986 => x"08001b04",
			3987 => x"009c3eb9",
			3988 => x"fea43eb9",
			3989 => x"019a3eb9",
			3990 => x"fe9f3eb9",
			3991 => x"0e007508",
			3992 => x"0a003604",
			3993 => x"01663eb9",
			3994 => x"fe9f3eb9",
			3995 => x"07002b0c",
			3996 => x"09001908",
			3997 => x"0600a004",
			3998 => x"008b3eb9",
			3999 => x"ff093eb9",
			4000 => x"fe473eb9",
			4001 => x"0e008710",
			4002 => x"00012908",
			4003 => x"02010f04",
			4004 => x"00db3eb9",
			4005 => x"ff033eb9",
			4006 => x"0c001804",
			4007 => x"00773eb9",
			4008 => x"017c3eb9",
			4009 => x"01000704",
			4010 => x"00a93eb9",
			4011 => x"08001c04",
			4012 => x"fea93eb9",
			4013 => x"00013eb9",
			4014 => x"00010e24",
			4015 => x"09001c18",
			4016 => x"08001804",
			4017 => x"ff143f95",
			4018 => x"08001b0c",
			4019 => x"06004404",
			4020 => x"ffd43f95",
			4021 => x"0e006a04",
			4022 => x"00ee3f95",
			4023 => x"00123f95",
			4024 => x"06009204",
			4025 => x"ff5a3f95",
			4026 => x"00743f95",
			4027 => x"0d001208",
			4028 => x"04001e04",
			4029 => x"00673f95",
			4030 => x"ffeb3f95",
			4031 => x"fecd3f95",
			4032 => x"0600a828",
			4033 => x"03002408",
			4034 => x"0d001204",
			4035 => x"00763f95",
			4036 => x"ff2b3f95",
			4037 => x"0600a314",
			4038 => x"0a003108",
			4039 => x"04001e04",
			4040 => x"00033f95",
			4041 => x"00c33f95",
			4042 => x"00012a08",
			4043 => x"05004104",
			4044 => x"fef03f95",
			4045 => x"00553f95",
			4046 => x"00623f95",
			4047 => x"02012e08",
			4048 => x"05003a04",
			4049 => x"01103f95",
			4050 => x"ffc53f95",
			4051 => x"ff5a3f95",
			4052 => x"0f00c704",
			4053 => x"ff0c3f95",
			4054 => x"0300270c",
			4055 => x"01000b08",
			4056 => x"03002404",
			4057 => x"00663f95",
			4058 => x"ff7b3f95",
			4059 => x"feef3f95",
			4060 => x"0e009308",
			4061 => x"09001c04",
			4062 => x"ffd03f95",
			4063 => x"00f53f95",
			4064 => x"03002904",
			4065 => x"00a23f95",
			4066 => x"09002204",
			4067 => x"fefe3f95",
			4068 => x"002e3f95",
			4069 => x"0000f320",
			4070 => x"0400080c",
			4071 => x"04000704",
			4072 => x"ffe04069",
			4073 => x"06002404",
			4074 => x"fffb4069",
			4075 => x"005c4069",
			4076 => x"0500360c",
			4077 => x"0d001704",
			4078 => x"ff184069",
			4079 => x"0d001804",
			4080 => x"001b4069",
			4081 => x"ffe34069",
			4082 => x"05003904",
			4083 => x"00474069",
			4084 => x"ffb14069",
			4085 => x"0600a92c",
			4086 => x"07002b10",
			4087 => x"06009504",
			4088 => x"00784069",
			4089 => x"0c001408",
			4090 => x"08001804",
			4091 => x"004c4069",
			4092 => x"ffc74069",
			4093 => x"ff0f4069",
			4094 => x"05002a04",
			4095 => x"00e44069",
			4096 => x"0201190c",
			4097 => x"0c001904",
			4098 => x"ff5d4069",
			4099 => x"00011404",
			4100 => x"ffe34069",
			4101 => x"006d4069",
			4102 => x"00013b08",
			4103 => x"09002204",
			4104 => x"00914069",
			4105 => x"ffdc4069",
			4106 => x"ffbd4069",
			4107 => x"02012804",
			4108 => x"ff2d4069",
			4109 => x"07002c04",
			4110 => x"ff594069",
			4111 => x"0700340c",
			4112 => x"03002d08",
			4113 => x"01000904",
			4114 => x"00d84069",
			4115 => x"00214069",
			4116 => x"ffdd4069",
			4117 => x"05003404",
			4118 => x"ff334069",
			4119 => x"05003804",
			4120 => x"00944069",
			4121 => x"ff954069",
			4122 => x"03003530",
			4123 => x"09001508",
			4124 => x"04001204",
			4125 => x"05a540cd",
			4126 => x"015140cd",
			4127 => x"03002104",
			4128 => x"fe6a40cd",
			4129 => x"01001320",
			4130 => x"0b001710",
			4131 => x"09001e08",
			4132 => x"05002e04",
			4133 => x"fff340cd",
			4134 => x"00de40cd",
			4135 => x"01000c04",
			4136 => x"002a40cd",
			4137 => x"fe1040cd",
			4138 => x"01000908",
			4139 => x"05002b04",
			4140 => x"014140cd",
			4141 => x"fdef40cd",
			4142 => x"05003604",
			4143 => x"008940cd",
			4144 => x"01f640cd",
			4145 => x"fe6d40cd",
			4146 => x"fe4840cd",
			4147 => x"0201051c",
			4148 => x"0200e914",
			4149 => x"09001504",
			4150 => x"ffec4169",
			4151 => x"0c00170c",
			4152 => x"08001c04",
			4153 => x"fe594169",
			4154 => x"0c001604",
			4155 => x"fe614169",
			4156 => x"01cb4169",
			4157 => x"fe584169",
			4158 => x"07002b04",
			4159 => x"02134169",
			4160 => x"fe5b4169",
			4161 => x"09002330",
			4162 => x"0e00972c",
			4163 => x"0500270c",
			4164 => x"0d001104",
			4165 => x"07b14169",
			4166 => x"03002104",
			4167 => x"fe654169",
			4168 => x"045c4169",
			4169 => x"09001c10",
			4170 => x"00013a08",
			4171 => x"04002004",
			4172 => x"04f94169",
			4173 => x"fe544169",
			4174 => x"0c001404",
			4175 => x"ffd14169",
			4176 => x"fe4b4169",
			4177 => x"0d001808",
			4178 => x"0f00c704",
			4179 => x"03df4169",
			4180 => x"072c4169",
			4181 => x"09002104",
			4182 => x"03784169",
			4183 => x"000e4169",
			4184 => x"fe624169",
			4185 => x"fe594169",
			4186 => x"0000f310",
			4187 => x"0d001704",
			4188 => x"ff9b4235",
			4189 => x"0d001808",
			4190 => x"01000c04",
			4191 => x"ffef4235",
			4192 => x"00204235",
			4193 => x"ffe94235",
			4194 => x"0800223c",
			4195 => x"0b001418",
			4196 => x"0e007904",
			4197 => x"003a4235",
			4198 => x"07002d0c",
			4199 => x"01000504",
			4200 => x"00114235",
			4201 => x"01000a04",
			4202 => x"ff694235",
			4203 => x"ffff4235",
			4204 => x"01000a04",
			4205 => x"00304235",
			4206 => x"ffe04235",
			4207 => x"0f00c314",
			4208 => x"04001e08",
			4209 => x"0600a004",
			4210 => x"00134235",
			4211 => x"ff714235",
			4212 => x"07003608",
			4213 => x"0a003e04",
			4214 => x"00574235",
			4215 => x"ffe44235",
			4216 => x"ffd14235",
			4217 => x"0e00970c",
			4218 => x"09001f08",
			4219 => x"0a003104",
			4220 => x"008d4235",
			4221 => x"ffdc4235",
			4222 => x"00074235",
			4223 => x"ffd04235",
			4224 => x"04002b10",
			4225 => x"0f00b804",
			4226 => x"000d4235",
			4227 => x"00014804",
			4228 => x"ff964235",
			4229 => x"00014b04",
			4230 => x"00074235",
			4231 => x"fffa4235",
			4232 => x"0f00bb04",
			4233 => x"ffe54235",
			4234 => x"0f00be04",
			4235 => x"002e4235",
			4236 => x"fffc4235",
			4237 => x"03002e5c",
			4238 => x"00011928",
			4239 => x"0c001510",
			4240 => x"05001004",
			4241 => x"00244341",
			4242 => x"0a002804",
			4243 => x"ff544341",
			4244 => x"04001a04",
			4245 => x"000f4341",
			4246 => x"fffd4341",
			4247 => x"0a002f14",
			4248 => x"0000cc08",
			4249 => x"03002b04",
			4250 => x"ffa04341",
			4251 => x"00264341",
			4252 => x"08001d08",
			4253 => x"07003004",
			4254 => x"009d4341",
			4255 => x"fff74341",
			4256 => x"ffcc4341",
			4257 => x"ff934341",
			4258 => x"0d001624",
			4259 => x"0b001518",
			4260 => x"0600ae0c",
			4261 => x"02012f08",
			4262 => x"02012b04",
			4263 => x"001f4341",
			4264 => x"00a64341",
			4265 => x"ffb74341",
			4266 => x"0e009004",
			4267 => x"ff574341",
			4268 => x"09001904",
			4269 => x"ffd24341",
			4270 => x"00494341",
			4271 => x"0d001304",
			4272 => x"fff14341",
			4273 => x"04002004",
			4274 => x"00ca4341",
			4275 => x"00004341",
			4276 => x"05002d04",
			4277 => x"ff6d4341",
			4278 => x"04002608",
			4279 => x"07003804",
			4280 => x"00744341",
			4281 => x"fff74341",
			4282 => x"ffd64341",
			4283 => x"0c001b18",
			4284 => x"04002e10",
			4285 => x"0f00c908",
			4286 => x"08001804",
			4287 => x"00004341",
			4288 => x"ff494341",
			4289 => x"0f00d404",
			4290 => x"00244341",
			4291 => x"ffde4341",
			4292 => x"04003204",
			4293 => x"00464341",
			4294 => x"ffd54341",
			4295 => x"0d001a0c",
			4296 => x"0b001b08",
			4297 => x"00010a04",
			4298 => x"fff44341",
			4299 => x"00814341",
			4300 => x"ffe14341",
			4301 => x"01000d04",
			4302 => x"001b4341",
			4303 => x"ffba4341",
			4304 => x"03001008",
			4305 => x"06002d04",
			4306 => x"ff0b43dd",
			4307 => x"054243dd",
			4308 => x"05003a38",
			4309 => x"08001508",
			4310 => x"07002104",
			4311 => x"000243dd",
			4312 => x"fe4b43dd",
			4313 => x"08001810",
			4314 => x"00011104",
			4315 => x"fe6143dd",
			4316 => x"05002c08",
			4317 => x"0a002c04",
			4318 => x"019e43dd",
			4319 => x"00d743dd",
			4320 => x"ffeb43dd",
			4321 => x"0c001610",
			4322 => x"0a002a08",
			4323 => x"04001e04",
			4324 => x"ff8443dd",
			4325 => x"017843dd",
			4326 => x"04001a04",
			4327 => x"ffd843dd",
			4328 => x"fea043dd",
			4329 => x"05003608",
			4330 => x"08002004",
			4331 => x"005443dd",
			4332 => x"ff2c43dd",
			4333 => x"0b001704",
			4334 => x"fedc43dd",
			4335 => x"018543dd",
			4336 => x"0b001708",
			4337 => x"0d001404",
			4338 => x"febc43dd",
			4339 => x"011843dd",
			4340 => x"04002704",
			4341 => x"005543dd",
			4342 => x"fe4c43dd",
			4343 => x"09001504",
			4344 => x"01a64451",
			4345 => x"03002104",
			4346 => x"fe7c4451",
			4347 => x"05002414",
			4348 => x"0a002808",
			4349 => x"09001c04",
			4350 => x"01db4451",
			4351 => x"ff824451",
			4352 => x"09001b04",
			4353 => x"feed4451",
			4354 => x"08001f04",
			4355 => x"016a4451",
			4356 => x"ffa44451",
			4357 => x"0a003e1c",
			4358 => x"0600a90c",
			4359 => x"03002304",
			4360 => x"fe7e4451",
			4361 => x"0f00c604",
			4362 => x"002f4451",
			4363 => x"01444451",
			4364 => x"0f00c708",
			4365 => x"05003604",
			4366 => x"fe0f4451",
			4367 => x"ff4c4451",
			4368 => x"01000704",
			4369 => x"01464451",
			4370 => x"ffc14451",
			4371 => x"fe884451",
			4372 => x"00010e24",
			4373 => x"0700291c",
			4374 => x"0b001510",
			4375 => x"04000804",
			4376 => x"0033454d",
			4377 => x"01000508",
			4378 => x"05002404",
			4379 => x"0033454d",
			4380 => x"ffcb454d",
			4381 => x"ff68454d",
			4382 => x"07002604",
			4383 => x"ffc9454d",
			4384 => x"0c001704",
			4385 => x"0089454d",
			4386 => x"ffe4454d",
			4387 => x"09001a04",
			4388 => x"fff5454d",
			4389 => x"ff25454d",
			4390 => x"0f00c024",
			4391 => x"09001908",
			4392 => x"07002904",
			4393 => x"002b454d",
			4394 => x"00b7454d",
			4395 => x"01000a08",
			4396 => x"0f00b404",
			4397 => x"002e454d",
			4398 => x"ff4a454d",
			4399 => x"0f00ba0c",
			4400 => x"00011804",
			4401 => x"0052454d",
			4402 => x"0b001804",
			4403 => x"ff78454d",
			4404 => x"0023454d",
			4405 => x"09002104",
			4406 => x"00ca454d",
			4407 => x"ffdf454d",
			4408 => x"0f00c714",
			4409 => x"0400230c",
			4410 => x"0d001104",
			4411 => x"0018454d",
			4412 => x"0b001704",
			4413 => x"ff19454d",
			4414 => x"ffe8454d",
			4415 => x"03003104",
			4416 => x"005e454d",
			4417 => x"ffd2454d",
			4418 => x"0e009314",
			4419 => x"05002a08",
			4420 => x"01000a04",
			4421 => x"004b454d",
			4422 => x"ff5a454d",
			4423 => x"0600af08",
			4424 => x"0d001304",
			4425 => x"0022454d",
			4426 => x"00ce454d",
			4427 => x"0011454d",
			4428 => x"07003004",
			4429 => x"002e454d",
			4430 => x"09002204",
			4431 => x"ff3f454d",
			4432 => x"0600b404",
			4433 => x"0040454d",
			4434 => x"ffde454d",
			4435 => x"00010e1c",
			4436 => x"07002b18",
			4437 => x"08001804",
			4438 => x"ffa64611",
			4439 => x"0f008b10",
			4440 => x"04000804",
			4441 => x"002f4611",
			4442 => x"05003604",
			4443 => x"ffa14611",
			4444 => x"05003b04",
			4445 => x"001f4611",
			4446 => x"ffe64611",
			4447 => x"00604611",
			4448 => x"ff844611",
			4449 => x"0d001630",
			4450 => x"07002b10",
			4451 => x"0e007704",
			4452 => x"00554611",
			4453 => x"04001804",
			4454 => x"00094611",
			4455 => x"0600a004",
			4456 => x"ffea4611",
			4457 => x"ff6e4611",
			4458 => x"0a003214",
			4459 => x"0e009810",
			4460 => x"04001d08",
			4461 => x"0b001404",
			4462 => x"00144611",
			4463 => x"00ad4611",
			4464 => x"04001e04",
			4465 => x"ffce4611",
			4466 => x"00574611",
			4467 => x"ffd44611",
			4468 => x"04002708",
			4469 => x"0e008504",
			4470 => x"00114611",
			4471 => x"ff934611",
			4472 => x"00354611",
			4473 => x"00011804",
			4474 => x"005e4611",
			4475 => x"05002c04",
			4476 => x"ff5f4611",
			4477 => x"0500380c",
			4478 => x"02012504",
			4479 => x"ffcc4611",
			4480 => x"04002304",
			4481 => x"00854611",
			4482 => x"fffc4611",
			4483 => x"ff8d4611",
			4484 => x"0800225c",
			4485 => x"0c001630",
			4486 => x"04002028",
			4487 => x"0f00cc1c",
			4488 => x"00011910",
			4489 => x"0c001508",
			4490 => x"05001204",
			4491 => x"001e46f5",
			4492 => x"ff7b46f5",
			4493 => x"05002404",
			4494 => x"004746f5",
			4495 => x"ffe346f5",
			4496 => x"0a002c04",
			4497 => x"008d46f5",
			4498 => x"0e008104",
			4499 => x"fff346f5",
			4500 => x"002446f5",
			4501 => x"04001908",
			4502 => x"04001504",
			4503 => x"ffc946f5",
			4504 => x"006546f5",
			4505 => x"ff5d46f5",
			4506 => x"0b001504",
			4507 => x"ff5346f5",
			4508 => x"fff946f5",
			4509 => x"02012820",
			4510 => x"06009e18",
			4511 => x"0c00170c",
			4512 => x"0a002f08",
			4513 => x"07002604",
			4514 => x"ffe646f5",
			4515 => x"009046f5",
			4516 => x"ffc646f5",
			4517 => x"08001d04",
			4518 => x"ff8646f5",
			4519 => x"0d001604",
			4520 => x"006e46f5",
			4521 => x"ffbb46f5",
			4522 => x"04001a04",
			4523 => x"fff846f5",
			4524 => x"ff8546f5",
			4525 => x"0e009308",
			4526 => x"05003504",
			4527 => x"00b646f5",
			4528 => x"ffec46f5",
			4529 => x"ffc546f5",
			4530 => x"0600a80c",
			4531 => x"00012d08",
			4532 => x"0e008a04",
			4533 => x"ffa046f5",
			4534 => x"001846f5",
			4535 => x"006546f5",
			4536 => x"04002804",
			4537 => x"ff5846f5",
			4538 => x"04002904",
			4539 => x"001746f5",
			4540 => x"fff646f5",
			4541 => x"02011940",
			4542 => x"0f00b430",
			4543 => x"00011124",
			4544 => x"05002510",
			4545 => x"0c001508",
			4546 => x"03001004",
			4547 => x"004a4809",
			4548 => x"ff454809",
			4549 => x"0200c204",
			4550 => x"ffaa4809",
			4551 => x"00c94809",
			4552 => x"05003008",
			4553 => x"04002204",
			4554 => x"fef34809",
			4555 => x"000b4809",
			4556 => x"0a003608",
			4557 => x"0d001504",
			4558 => x"00a24809",
			4559 => x"ffb84809",
			4560 => x"ff7e4809",
			4561 => x"0e007a04",
			4562 => x"00e44809",
			4563 => x"06009a04",
			4564 => x"ff9a4809",
			4565 => x"002c4809",
			4566 => x"0b001808",
			4567 => x"08001904",
			4568 => x"ffd14809",
			4569 => x"fee24809",
			4570 => x"0600a604",
			4571 => x"00874809",
			4572 => x"fffb4809",
			4573 => x"00013b28",
			4574 => x"02012b20",
			4575 => x"0b001510",
			4576 => x"09001908",
			4577 => x"02012304",
			4578 => x"00f94809",
			4579 => x"ffa94809",
			4580 => x"01000904",
			4581 => x"feea4809",
			4582 => x"ffd64809",
			4583 => x"0e00900c",
			4584 => x"0f00bb04",
			4585 => x"ffe64809",
			4586 => x"08002304",
			4587 => x"00fa4809",
			4588 => x"00094809",
			4589 => x"ff8c4809",
			4590 => x"03002e04",
			4591 => x"00f34809",
			4592 => x"ffb14809",
			4593 => x"0f00c808",
			4594 => x"0c001604",
			4595 => x"fff74809",
			4596 => x"ff324809",
			4597 => x"0700340c",
			4598 => x"09001c08",
			4599 => x"05002804",
			4600 => x"00674809",
			4601 => x"fefe4809",
			4602 => x"00904809",
			4603 => x"03003104",
			4604 => x"ff194809",
			4605 => x"03003408",
			4606 => x"02013a04",
			4607 => x"00614809",
			4608 => x"fff34809",
			4609 => x"ffb64809",
			4610 => x"0201193c",
			4611 => x"0f00b430",
			4612 => x"00011124",
			4613 => x"05002510",
			4614 => x"0c001508",
			4615 => x"03001004",
			4616 => x"004e490d",
			4617 => x"ff3c490d",
			4618 => x"0200c204",
			4619 => x"ffa6490d",
			4620 => x"00d4490d",
			4621 => x"05003008",
			4622 => x"04002204",
			4623 => x"fee9490d",
			4624 => x"000d490d",
			4625 => x"0a003608",
			4626 => x"0d001504",
			4627 => x"00aa490d",
			4628 => x"ffb4490d",
			4629 => x"ff78490d",
			4630 => x"0e007a04",
			4631 => x"00ef490d",
			4632 => x"06009a04",
			4633 => x"ff94490d",
			4634 => x"0032490d",
			4635 => x"0b001804",
			4636 => x"fee7490d",
			4637 => x"0600a604",
			4638 => x"008c490d",
			4639 => x"fffb490d",
			4640 => x"00013b24",
			4641 => x"07002b08",
			4642 => x"05002b04",
			4643 => x"0032490d",
			4644 => x"ff3b490d",
			4645 => x"0e009018",
			4646 => x"0b001508",
			4647 => x"09001a04",
			4648 => x"00b6490d",
			4649 => x"ffc1490d",
			4650 => x"03003308",
			4651 => x"08002304",
			4652 => x"0115490d",
			4653 => x"ffb2490d",
			4654 => x"0f00bc04",
			4655 => x"003e490d",
			4656 => x"ff8b490d",
			4657 => x"ff72490d",
			4658 => x"0f00c808",
			4659 => x"0c001604",
			4660 => x"fff7490d",
			4661 => x"ff26490d",
			4662 => x"0700340c",
			4663 => x"09001c08",
			4664 => x"05002804",
			4665 => x"006e490d",
			4666 => x"fef5490d",
			4667 => x"009a490d",
			4668 => x"03003104",
			4669 => x"ff0f490d",
			4670 => x"03003408",
			4671 => x"02013a04",
			4672 => x"0068490d",
			4673 => x"fff3490d",
			4674 => x"ffb5490d",
			4675 => x"0600a84c",
			4676 => x"02011f3c",
			4677 => x"0a002f24",
			4678 => x"0e007e1c",
			4679 => x"0a00280c",
			4680 => x"09001504",
			4681 => x"003749f1",
			4682 => x"05002a04",
			4683 => x"ff9649f1",
			4684 => x"001349f1",
			4685 => x"0d001508",
			4686 => x"0c001804",
			4687 => x"00a849f1",
			4688 => x"fff949f1",
			4689 => x"0d001704",
			4690 => x"ffd049f1",
			4691 => x"001949f1",
			4692 => x"0e008204",
			4693 => x"ffad49f1",
			4694 => x"000d49f1",
			4695 => x"0500420c",
			4696 => x"0e008a08",
			4697 => x"04001f04",
			4698 => x"000349f1",
			4699 => x"ff6249f1",
			4700 => x"001149f1",
			4701 => x"05004708",
			4702 => x"07002904",
			4703 => x"fff749f1",
			4704 => x"002c49f1",
			4705 => x"ffe149f1",
			4706 => x"0e007d04",
			4707 => x"ffa649f1",
			4708 => x"00013b08",
			4709 => x"0a003804",
			4710 => x"00a649f1",
			4711 => x"fff649f1",
			4712 => x"ffd749f1",
			4713 => x"01000704",
			4714 => x"001a49f1",
			4715 => x"09001c08",
			4716 => x"0f00df04",
			4717 => x"ff4849f1",
			4718 => x"000349f1",
			4719 => x"09001f08",
			4720 => x"0a003104",
			4721 => x"006349f1",
			4722 => x"ffd249f1",
			4723 => x"04002508",
			4724 => x"0b001b04",
			4725 => x"ff7449f1",
			4726 => x"001349f1",
			4727 => x"00014104",
			4728 => x"ffcc49f1",
			4729 => x"04002904",
			4730 => x"005b49f1",
			4731 => x"ffea49f1",
			4732 => x"00010e04",
			4733 => x"ff954aa5",
			4734 => x"0a00312c",
			4735 => x"0a002808",
			4736 => x"0d001204",
			4737 => x"002e4aa5",
			4738 => x"ffc74aa5",
			4739 => x"0800201c",
			4740 => x"0b001410",
			4741 => x"03002608",
			4742 => x"0600b304",
			4743 => x"00494aa5",
			4744 => x"00034aa5",
			4745 => x"02012304",
			4746 => x"00034aa5",
			4747 => x"ffba4aa5",
			4748 => x"04002208",
			4749 => x"0600a304",
			4750 => x"000b4aa5",
			4751 => x"00994aa5",
			4752 => x"00014aa5",
			4753 => x"00013f04",
			4754 => x"ffd84aa5",
			4755 => x"00044aa5",
			4756 => x"0b001818",
			4757 => x"03002e0c",
			4758 => x"0c001708",
			4759 => x"0f00c204",
			4760 => x"000a4aa5",
			4761 => x"ffba4aa5",
			4762 => x"00354aa5",
			4763 => x"0e007e04",
			4764 => x"00074aa5",
			4765 => x"0f00c804",
			4766 => x"ff8b4aa5",
			4767 => x"fffd4aa5",
			4768 => x"0d001a08",
			4769 => x"0e008e04",
			4770 => x"00624aa5",
			4771 => x"fffe4aa5",
			4772 => x"04002308",
			4773 => x"00013904",
			4774 => x"00274aa5",
			4775 => x"fff14aa5",
			4776 => x"ffc04aa5",
			4777 => x"0400263c",
			4778 => x"04002538",
			4779 => x"04002330",
			4780 => x"0000f31c",
			4781 => x"0400080c",
			4782 => x"04000704",
			4783 => x"ffd74b71",
			4784 => x"01000804",
			4785 => x"007c4b71",
			4786 => x"fff94b71",
			4787 => x"0d001708",
			4788 => x"09001c04",
			4789 => x"ff1a4b71",
			4790 => x"ffca4b71",
			4791 => x"04001b04",
			4792 => x"00634b71",
			4793 => x"ffb44b71",
			4794 => x"0e007504",
			4795 => x"00c54b71",
			4796 => x"0e007c08",
			4797 => x"09001904",
			4798 => x"003a4b71",
			4799 => x"fed94b71",
			4800 => x"0b001404",
			4801 => x"ff9b4b71",
			4802 => x"00474b71",
			4803 => x"09001f04",
			4804 => x"001e4b71",
			4805 => x"ff094b71",
			4806 => x"00f54b71",
			4807 => x"04002b14",
			4808 => x"0500390c",
			4809 => x"0f00cb04",
			4810 => x"ff1a4b71",
			4811 => x"0f00d304",
			4812 => x"00334b71",
			4813 => x"ff9d4b71",
			4814 => x"05003a04",
			4815 => x"00584b71",
			4816 => x"ff854b71",
			4817 => x"04003214",
			4818 => x"0c001804",
			4819 => x"ffb44b71",
			4820 => x"0200ef04",
			4821 => x"ffde4b71",
			4822 => x"04002e08",
			4823 => x"00012e04",
			4824 => x"ff904b71",
			4825 => x"00874b71",
			4826 => x"00b14b71",
			4827 => x"ff794b71",
			4828 => x"00010e24",
			4829 => x"0400080c",
			4830 => x"04000704",
			4831 => x"ffe34c65",
			4832 => x"01000804",
			4833 => x"00524c65",
			4834 => x"fffc4c65",
			4835 => x"05003008",
			4836 => x"03002c04",
			4837 => x"ff5e4c65",
			4838 => x"ffe94c65",
			4839 => x"01000904",
			4840 => x"ffaf4c65",
			4841 => x"0c001908",
			4842 => x"07002604",
			4843 => x"ffe54c65",
			4844 => x"00794c65",
			4845 => x"ffcd4c65",
			4846 => x"0f00c024",
			4847 => x"0c001404",
			4848 => x"00ae4c65",
			4849 => x"01000a08",
			4850 => x"0f00b404",
			4851 => x"004e4c65",
			4852 => x"ff444c65",
			4853 => x"0400260c",
			4854 => x"01000d04",
			4855 => x"00e04c65",
			4856 => x"0f00bb04",
			4857 => x"ffa44c65",
			4858 => x"00684c65",
			4859 => x"0c001c04",
			4860 => x"ff844c65",
			4861 => x"00012e04",
			4862 => x"fff84c65",
			4863 => x"00584c65",
			4864 => x"02012b18",
			4865 => x"0a002a04",
			4866 => x"00104c65",
			4867 => x"0c001808",
			4868 => x"0f00c704",
			4869 => x"fef34c65",
			4870 => x"ffc84c65",
			4871 => x"0f00c204",
			4872 => x"ffd64c65",
			4873 => x"0f00c704",
			4874 => x"005e4c65",
			4875 => x"fffc4c65",
			4876 => x"00013a04",
			4877 => x"00b44c65",
			4878 => x"0e008808",
			4879 => x"08001b04",
			4880 => x"ff3f4c65",
			4881 => x"fff64c65",
			4882 => x"07003308",
			4883 => x"09001c04",
			4884 => x"00064c65",
			4885 => x"00944c65",
			4886 => x"0a003604",
			4887 => x"ff604c65",
			4888 => x"00044c65",
			4889 => x"0900191c",
			4890 => x"0600a814",
			4891 => x"0001190c",
			4892 => x"0a002508",
			4893 => x"04000804",
			4894 => x"00304d61",
			4895 => x"ff6e4d61",
			4896 => x"00394d61",
			4897 => x"04001f04",
			4898 => x"00cc4d61",
			4899 => x"00134d61",
			4900 => x"0c001404",
			4901 => x"ff7f4d61",
			4902 => x"002c4d61",
			4903 => x"0c00183c",
			4904 => x"0a002f2c",
			4905 => x"0c001618",
			4906 => x"07002c0c",
			4907 => x"08001c04",
			4908 => x"ff3f4d61",
			4909 => x"08001d04",
			4910 => x"001e4d61",
			4911 => x"ffde4d61",
			4912 => x"07002e04",
			4913 => x"007a4d61",
			4914 => x"0e009204",
			4915 => x"ff7e4d61",
			4916 => x"002d4d61",
			4917 => x"07002c0c",
			4918 => x"0c001708",
			4919 => x"07002604",
			4920 => x"ffde4d61",
			4921 => x"00c54d61",
			4922 => x"ffcb4d61",
			4923 => x"0e008804",
			4924 => x"ff694d61",
			4925 => x"003b4d61",
			4926 => x"04001b04",
			4927 => x"00284d61",
			4928 => x"0b001708",
			4929 => x"09001a04",
			4930 => x"fffb4d61",
			4931 => x"ff2b4d61",
			4932 => x"00174d61",
			4933 => x"08001c10",
			4934 => x"0b00170c",
			4935 => x"08001b08",
			4936 => x"0d001404",
			4937 => x"fff34d61",
			4938 => x"00504d61",
			4939 => x"ffd74d61",
			4940 => x"ff6c4d61",
			4941 => x"01001314",
			4942 => x"05002c04",
			4943 => x"ffae4d61",
			4944 => x"00012d08",
			4945 => x"01000d04",
			4946 => x"00584d61",
			4947 => x"ff914d61",
			4948 => x"0e009404",
			4949 => x"00cc4d61",
			4950 => x"ffe14d61",
			4951 => x"ffa24d61",
			4952 => x"0f008b0c",
			4953 => x"0c001708",
			4954 => x"0b001704",
			4955 => x"fe664e05",
			4956 => x"015d4e05",
			4957 => x"fe654e05",
			4958 => x"08002340",
			4959 => x"03003538",
			4960 => x"0c001620",
			4961 => x"09001910",
			4962 => x"0f00c308",
			4963 => x"00011104",
			4964 => x"ff654e05",
			4965 => x"01f44e05",
			4966 => x"0b001304",
			4967 => x"fe354e05",
			4968 => x"00de4e05",
			4969 => x"0a002c08",
			4970 => x"0a002704",
			4971 => x"fe224e05",
			4972 => x"00bd4e05",
			4973 => x"0e008904",
			4974 => x"fe294e05",
			4975 => x"ffa04e05",
			4976 => x"0e009010",
			4977 => x"02012a08",
			4978 => x"01000d04",
			4979 => x"01824e05",
			4980 => x"ffbd4e05",
			4981 => x"02012e04",
			4982 => x"030c4e05",
			4983 => x"016b4e05",
			4984 => x"00014404",
			4985 => x"fe2a4e05",
			4986 => x"01294e05",
			4987 => x"07003004",
			4988 => x"ff604e05",
			4989 => x"fe0e4e05",
			4990 => x"09002204",
			4991 => x"ffad4e05",
			4992 => x"fe654e05",
			4993 => x"0f00c058",
			4994 => x"00010e34",
			4995 => x"04001c1c",
			4996 => x"04001a10",
			4997 => x"04000808",
			4998 => x"04000704",
			4999 => x"ffef4f29",
			5000 => x"00314f29",
			5001 => x"0f00ac04",
			5002 => x"ffb14f29",
			5003 => x"00014f29",
			5004 => x"07002704",
			5005 => x"fff64f29",
			5006 => x"07002e04",
			5007 => x"00544f29",
			5008 => x"fff74f29",
			5009 => x"09001f08",
			5010 => x"0e007b04",
			5011 => x"ff894f29",
			5012 => x"fffb4f29",
			5013 => x"0b00180c",
			5014 => x"0b001704",
			5015 => x"ffeb4f29",
			5016 => x"09002004",
			5017 => x"00394f29",
			5018 => x"fffc4f29",
			5019 => x"ffda4f29",
			5020 => x"04002614",
			5021 => x"0a002804",
			5022 => x"fffa4f29",
			5023 => x"01000604",
			5024 => x"00054f29",
			5025 => x"01000d04",
			5026 => x"00984f29",
			5027 => x"0d001a04",
			5028 => x"001f4f29",
			5029 => x"ffed4f29",
			5030 => x"03003408",
			5031 => x"0e008a04",
			5032 => x"ffa84f29",
			5033 => x"00014f29",
			5034 => x"03003804",
			5035 => x"00424f29",
			5036 => x"ffea4f29",
			5037 => x"0f00c710",
			5038 => x"0d001208",
			5039 => x"0a002d04",
			5040 => x"00294f29",
			5041 => x"ffb24f29",
			5042 => x"0d001b04",
			5043 => x"ff6e4f29",
			5044 => x"000f4f29",
			5045 => x"01000704",
			5046 => x"00664f29",
			5047 => x"09001c0c",
			5048 => x"00015508",
			5049 => x"04001604",
			5050 => x"fff74f29",
			5051 => x"ff5c4f29",
			5052 => x"001f4f29",
			5053 => x"0600b40c",
			5054 => x"0d001804",
			5055 => x"00894f29",
			5056 => x"02012b04",
			5057 => x"00044f29",
			5058 => x"ffc44f29",
			5059 => x"0f00d908",
			5060 => x"0a003604",
			5061 => x"ff9d4f29",
			5062 => x"00094f29",
			5063 => x"02014204",
			5064 => x"00214f29",
			5065 => x"fff54f29",
			5066 => x"0f00c044",
			5067 => x"02012038",
			5068 => x"0a002f20",
			5069 => x"0c00181c",
			5070 => x"0b00120c",
			5071 => x"01000b08",
			5072 => x"01000504",
			5073 => x"00055035",
			5074 => x"ffae5035",
			5075 => x"00155035",
			5076 => x"0a002808",
			5077 => x"00010f04",
			5078 => x"00395035",
			5079 => x"ffa95035",
			5080 => x"0000f304",
			5081 => x"fff95035",
			5082 => x"00ad5035",
			5083 => x"ffbf5035",
			5084 => x"02011d14",
			5085 => x"04002e08",
			5086 => x"07003704",
			5087 => x"ff605035",
			5088 => x"00135035",
			5089 => x"05004708",
			5090 => x"0e006e04",
			5091 => x"ffee5035",
			5092 => x"003d5035",
			5093 => x"ffdc5035",
			5094 => x"00125035",
			5095 => x"0d001a08",
			5096 => x"01000a04",
			5097 => x"001a5035",
			5098 => x"00a65035",
			5099 => x"ffdd5035",
			5100 => x"0f00c610",
			5101 => x"0a002a04",
			5102 => x"00285035",
			5103 => x"04002504",
			5104 => x"ff555035",
			5105 => x"05003b04",
			5106 => x"00175035",
			5107 => x"ffe95035",
			5108 => x"0600ae0c",
			5109 => x"0c001504",
			5110 => x"ffc85035",
			5111 => x"0b001604",
			5112 => x"00845035",
			5113 => x"fffd5035",
			5114 => x"09001d14",
			5115 => x"0f00de0c",
			5116 => x"03002d08",
			5117 => x"04001704",
			5118 => x"fffe5035",
			5119 => x"ff655035",
			5120 => x"000c5035",
			5121 => x"0f00e404",
			5122 => x"002f5035",
			5123 => x"ffed5035",
			5124 => x"04002308",
			5125 => x"0c001b04",
			5126 => x"009a5035",
			5127 => x"ffcc5035",
			5128 => x"0a003604",
			5129 => x"ff925035",
			5130 => x"0a003704",
			5131 => x"00355035",
			5132 => x"ffd85035",
			5133 => x"0600a85c",
			5134 => x"01000928",
			5135 => x"0c001410",
			5136 => x"0400200c",
			5137 => x"08001504",
			5138 => x"ffe25151",
			5139 => x"00011104",
			5140 => x"ffff5151",
			5141 => x"008f5151",
			5142 => x"ffdb5151",
			5143 => x"04001c10",
			5144 => x"0300240c",
			5145 => x"09001904",
			5146 => x"00225151",
			5147 => x"09001b04",
			5148 => x"ff965151",
			5149 => x"00135151",
			5150 => x"004a5151",
			5151 => x"08001d04",
			5152 => x"ff3a5151",
			5153 => x"001a5151",
			5154 => x"00012a28",
			5155 => x"01000d1c",
			5156 => x"0c00160c",
			5157 => x"08001b04",
			5158 => x"ffb75151",
			5159 => x"09001a04",
			5160 => x"001b5151",
			5161 => x"ffea5151",
			5162 => x"0f008b08",
			5163 => x"05003604",
			5164 => x"ffd05151",
			5165 => x"00185151",
			5166 => x"07003004",
			5167 => x"00875151",
			5168 => x"fff15151",
			5169 => x"01001c08",
			5170 => x"0e008a04",
			5171 => x"ff5c5151",
			5172 => x"00145151",
			5173 => x"001a5151",
			5174 => x"00013708",
			5175 => x"0d001804",
			5176 => x"00c95151",
			5177 => x"00215151",
			5178 => x"fffa5151",
			5179 => x"0f00c708",
			5180 => x"0a002f04",
			5181 => x"000e5151",
			5182 => x"ff485151",
			5183 => x"0600ae08",
			5184 => x"0d001304",
			5185 => x"ffea5151",
			5186 => x"009c5151",
			5187 => x"02013810",
			5188 => x"0c001804",
			5189 => x"ff485151",
			5190 => x"03002f08",
			5191 => x"03002d04",
			5192 => x"00005151",
			5193 => x"00455151",
			5194 => x"ffd15151",
			5195 => x"04002108",
			5196 => x"0600bd04",
			5197 => x"00635151",
			5198 => x"ffc95151",
			5199 => x"0a003604",
			5200 => x"ff925151",
			5201 => x"00014d04",
			5202 => x"004a5151",
			5203 => x"ffe75151",
			5204 => x"0e00944c",
			5205 => x"00014c48",
			5206 => x"0600a834",
			5207 => x"0e008520",
			5208 => x"09001910",
			5209 => x"0b001408",
			5210 => x"06009d04",
			5211 => x"009c5205",
			5212 => x"ff8a5205",
			5213 => x"08001804",
			5214 => x"01475205",
			5215 => x"00145205",
			5216 => x"03002408",
			5217 => x"0d001104",
			5218 => x"00235205",
			5219 => x"fec15205",
			5220 => x"01000604",
			5221 => x"fec55205",
			5222 => x"002d5205",
			5223 => x"02011e0c",
			5224 => x"07003704",
			5225 => x"feef5205",
			5226 => x"0a003704",
			5227 => x"fff75205",
			5228 => x"00d85205",
			5229 => x"05003a04",
			5230 => x"015d5205",
			5231 => x"ffa55205",
			5232 => x"02012804",
			5233 => x"feac5205",
			5234 => x"09001a04",
			5235 => x"fefe5205",
			5236 => x"00013b04",
			5237 => x"00b45205",
			5238 => x"0e008d04",
			5239 => x"001c5205",
			5240 => x"ff5f5205",
			5241 => x"00ce5205",
			5242 => x"09002204",
			5243 => x"feca5205",
			5244 => x"0600b408",
			5245 => x"0600b204",
			5246 => x"fffa5205",
			5247 => x"00ab5205",
			5248 => x"ff815205",
			5249 => x"01000414",
			5250 => x"0a002a0c",
			5251 => x"09001908",
			5252 => x"0a002004",
			5253 => x"ffe15301",
			5254 => x"00335301",
			5255 => x"ff6a5301",
			5256 => x"04002104",
			5257 => x"00db5301",
			5258 => x"ffb35301",
			5259 => x"0600a944",
			5260 => x"01000a24",
			5261 => x"05002910",
			5262 => x"0e00810c",
			5263 => x"0a002808",
			5264 => x"04000804",
			5265 => x"00585301",
			5266 => x"ff5a5301",
			5267 => x"00695301",
			5268 => x"00a45301",
			5269 => x"06009e0c",
			5270 => x"00011308",
			5271 => x"08001b04",
			5272 => x"00215301",
			5273 => x"ff7c5301",
			5274 => x"00835301",
			5275 => x"0f00c304",
			5276 => x"fecc5301",
			5277 => x"ffe95301",
			5278 => x"00012d18",
			5279 => x"0a002f10",
			5280 => x"04001808",
			5281 => x"0c001204",
			5282 => x"fffb5301",
			5283 => x"ff695301",
			5284 => x"08001f04",
			5285 => x"00b35301",
			5286 => x"ffa15301",
			5287 => x"0e008a04",
			5288 => x"ff135301",
			5289 => x"00645301",
			5290 => x"0b001904",
			5291 => x"00e75301",
			5292 => x"00065301",
			5293 => x"01000704",
			5294 => x"003d5301",
			5295 => x"05002e10",
			5296 => x"0001570c",
			5297 => x"04001608",
			5298 => x"04001504",
			5299 => x"ff935301",
			5300 => x"001e5301",
			5301 => x"fed75301",
			5302 => x"001a5301",
			5303 => x"05003810",
			5304 => x"08002208",
			5305 => x"0f00cc04",
			5306 => x"00da5301",
			5307 => x"00145301",
			5308 => x"03002904",
			5309 => x"001e5301",
			5310 => x"ff555301",
			5311 => x"ff2c5301",
			5312 => x"07003668",
			5313 => x"0b001734",
			5314 => x"08001f30",
			5315 => x"09001c1c",
			5316 => x"0600960c",
			5317 => x"00011008",
			5318 => x"08001804",
			5319 => x"ff3653e5",
			5320 => x"005c53e5",
			5321 => x"00d053e5",
			5322 => x"02012b08",
			5323 => x"0d001104",
			5324 => x"ffd053e5",
			5325 => x"ff1a53e5",
			5326 => x"00013c04",
			5327 => x"00ac53e5",
			5328 => x"ff9153e5",
			5329 => x"0e007c0c",
			5330 => x"0a002404",
			5331 => x"004c53e5",
			5332 => x"05004604",
			5333 => x"ff3553e5",
			5334 => x"002f53e5",
			5335 => x"03002a04",
			5336 => x"00bd53e5",
			5337 => x"001953e5",
			5338 => x"ff1553e5",
			5339 => x"01000910",
			5340 => x"05002b0c",
			5341 => x"0d001304",
			5342 => x"ffb453e5",
			5343 => x"07002904",
			5344 => x"fff953e5",
			5345 => x"008253e5",
			5346 => x"ff2853e5",
			5347 => x"00012a18",
			5348 => x"01000b0c",
			5349 => x"08001d04",
			5350 => x"ffbf53e5",
			5351 => x"0b001a04",
			5352 => x"00b953e5",
			5353 => x"fff553e5",
			5354 => x"0b001804",
			5355 => x"ff4e53e5",
			5356 => x"0d001a04",
			5357 => x"003353e5",
			5358 => x"ffe953e5",
			5359 => x"09002108",
			5360 => x"01001004",
			5361 => x"010053e5",
			5362 => x"006253e5",
			5363 => x"ffeb53e5",
			5364 => x"0e008b08",
			5365 => x"0d001b04",
			5366 => x"003c53e5",
			5367 => x"fff053e5",
			5368 => x"ff1053e5",
			5369 => x"0100136c",
			5370 => x"0c00162c",
			5371 => x"0400201c",
			5372 => x"01000c18",
			5373 => x"0b001208",
			5374 => x"0d000e04",
			5375 => x"ffc654c1",
			5376 => x"fed254c1",
			5377 => x"0f00bf08",
			5378 => x"08001904",
			5379 => x"00c654c1",
			5380 => x"ff4854c1",
			5381 => x"07002c04",
			5382 => x"fea354c1",
			5383 => x"006754c1",
			5384 => x"feba54c1",
			5385 => x"0b00150c",
			5386 => x"07002808",
			5387 => x"07002204",
			5388 => x"ff8f54c1",
			5389 => x"004554c1",
			5390 => x"fe7b54c1",
			5391 => x"003954c1",
			5392 => x"0f00c62c",
			5393 => x"01000910",
			5394 => x"08001d04",
			5395 => x"fe7754c1",
			5396 => x"05003108",
			5397 => x"07002904",
			5398 => x"fffa54c1",
			5399 => x"011554c1",
			5400 => x"ffc454c1",
			5401 => x"08001c0c",
			5402 => x"07002d08",
			5403 => x"0a003d04",
			5404 => x"016f54c1",
			5405 => x"ff4954c1",
			5406 => x"fecd54c1",
			5407 => x"04001e08",
			5408 => x"0e007e04",
			5409 => x"004154c1",
			5410 => x"fea754c1",
			5411 => x"00012d04",
			5412 => x"ffd454c1",
			5413 => x"00f854c1",
			5414 => x"0e009008",
			5415 => x"04002004",
			5416 => x"009154c1",
			5417 => x"013654c1",
			5418 => x"0f00d908",
			5419 => x"0a003604",
			5420 => x"fe7f54c1",
			5421 => x"00ac54c1",
			5422 => x"00c354c1",
			5423 => x"fec154c1",
			5424 => x"01001374",
			5425 => x"0c001634",
			5426 => x"04002024",
			5427 => x"01000c20",
			5428 => x"06009f10",
			5429 => x"0d001208",
			5430 => x"0b001204",
			5431 => x"ff6d55af",
			5432 => x"012355af",
			5433 => x"09001904",
			5434 => x"008455af",
			5435 => x"ff3d55af",
			5436 => x"01000808",
			5437 => x"0f00c704",
			5438 => x"fead55af",
			5439 => x"007455af",
			5440 => x"05002704",
			5441 => x"ff1d55af",
			5442 => x"010e55af",
			5443 => x"feb055af",
			5444 => x"0b00150c",
			5445 => x"07002808",
			5446 => x"07002204",
			5447 => x"ff8a55af",
			5448 => x"004f55af",
			5449 => x"fe7355af",
			5450 => x"004055af",
			5451 => x"0f00c62c",
			5452 => x"0100090c",
			5453 => x"08001d04",
			5454 => x"fe6f55af",
			5455 => x"07002d04",
			5456 => x"ffc255af",
			5457 => x"011c55af",
			5458 => x"08001c10",
			5459 => x"0c001808",
			5460 => x"0000cc04",
			5461 => x"ffa955af",
			5462 => x"018c55af",
			5463 => x"05004604",
			5464 => x"feb455af",
			5465 => x"008955af",
			5466 => x"04001e08",
			5467 => x"0e007e04",
			5468 => x"004755af",
			5469 => x"fe9155af",
			5470 => x"01000b04",
			5471 => x"017155af",
			5472 => x"fffa55af",
			5473 => x"0e009008",
			5474 => x"0d001504",
			5475 => x"009755af",
			5476 => x"013655af",
			5477 => x"0a003608",
			5478 => x"0f00d804",
			5479 => x"fe8755af",
			5480 => x"002c55af",
			5481 => x"00aa55af",
			5482 => x"feba55af",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1943, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3615, initial_addr_3'length));
	end generate gen_rom_3;

	gen_rom_4: if SELECT_ROM = 4 generate
		bank <= (
			0 => x"03002418",
			1 => x"0600930c",
			2 => x"05002704",
			3 => x"ffc40095",
			4 => x"05002904",
			5 => x"00180095",
			6 => x"fff30095",
			7 => x"00013808",
			8 => x"0e008504",
			9 => x"00860095",
			10 => x"00040095",
			11 => x"ffd70095",
			12 => x"0b00171c",
			13 => x"01000d14",
			14 => x"0200fd0c",
			15 => x"0f009204",
			16 => x"ffe10095",
			17 => x"05002704",
			18 => x"fffc0095",
			19 => x"00330095",
			20 => x"03003304",
			21 => x"ff760095",
			22 => x"000c0095",
			23 => x"09001c04",
			24 => x"002a0095",
			25 => x"ffd70095",
			26 => x"02012d08",
			27 => x"09001e04",
			28 => x"00260095",
			29 => x"ffb20095",
			30 => x"08002004",
			31 => x"00700095",
			32 => x"0c001e04",
			33 => x"ffd50095",
			34 => x"03003104",
			35 => x"fffb0095",
			36 => x"001d0095",
			37 => x"0d001424",
			38 => x"00011918",
			39 => x"08001b0c",
			40 => x"0f009204",
			41 => x"ffdb0139",
			42 => x"07002d04",
			43 => x"00820139",
			44 => x"ffeb0139",
			45 => x"07002404",
			46 => x"00170139",
			47 => x"0a002104",
			48 => x"000a0139",
			49 => x"ffb70139",
			50 => x"0e009a08",
			51 => x"0a002504",
			52 => x"fffb0139",
			53 => x"ff3c0139",
			54 => x"00240139",
			55 => x"02012018",
			56 => x"09001b08",
			57 => x"04001a04",
			58 => x"ffed0139",
			59 => x"00430139",
			60 => x"03002904",
			61 => x"ff710139",
			62 => x"04002108",
			63 => x"04002004",
			64 => x"ffeb0139",
			65 => x"004e0139",
			66 => x"ffbe0139",
			67 => x"01000c04",
			68 => x"007a0139",
			69 => x"04002608",
			70 => x"05002c04",
			71 => x"00140139",
			72 => x"ff950139",
			73 => x"00014304",
			74 => x"ffe10139",
			75 => x"07003f04",
			76 => x"004e0139",
			77 => x"fff60139",
			78 => x"05002a2c",
			79 => x"0c001514",
			80 => x"00011108",
			81 => x"0000e504",
			82 => x"ffbd01f5",
			83 => x"00ef01f5",
			84 => x"0600a504",
			85 => x"ff4501f5",
			86 => x"0e009104",
			87 => x"00cc01f5",
			88 => x"ff8801f5",
			89 => x"0300220c",
			90 => x"0b001708",
			91 => x"0f00b404",
			92 => x"ff6601f5",
			93 => x"00d501f5",
			94 => x"ff2901f5",
			95 => x"0b001904",
			96 => x"fecf01f5",
			97 => x"09002104",
			98 => x"007401f5",
			99 => x"ffe001f5",
			100 => x"0b001614",
			101 => x"05002f10",
			102 => x"0a002d08",
			103 => x"07002a04",
			104 => x"003501f5",
			105 => x"ff5301f5",
			106 => x"02013104",
			107 => x"00b901f5",
			108 => x"ffd101f5",
			109 => x"ff4601f5",
			110 => x"01000a08",
			111 => x"0f00ba04",
			112 => x"ffa801f5",
			113 => x"010e01f5",
			114 => x"07002f0c",
			115 => x"01000b04",
			116 => x"ffcb01f5",
			117 => x"09001f04",
			118 => x"00b901f5",
			119 => x"ffed01f5",
			120 => x"07003704",
			121 => x"fefe01f5",
			122 => x"0d001a04",
			123 => x"00be01f5",
			124 => x"ffaa01f5",
			125 => x"0e008234",
			126 => x"06009e28",
			127 => x"0c001610",
			128 => x"0f009204",
			129 => x"ffd002a9",
			130 => x"00011908",
			131 => x"05002404",
			132 => x"000202a9",
			133 => x"005402a9",
			134 => x"ffdc02a9",
			135 => x"07002408",
			136 => x"0d001204",
			137 => x"001402a9",
			138 => x"fff602a9",
			139 => x"01000c04",
			140 => x"ffa102a9",
			141 => x"0a002f04",
			142 => x"ffed02a9",
			143 => x"01001004",
			144 => x"001f02a9",
			145 => x"fffa02a9",
			146 => x"05002d08",
			147 => x"0f00c304",
			148 => x"008702a9",
			149 => x"fff402a9",
			150 => x"ffe002a9",
			151 => x"09001f14",
			152 => x"0d00130c",
			153 => x"0f00cb04",
			154 => x"ffc102a9",
			155 => x"0f00da04",
			156 => x"004302a9",
			157 => x"ffed02a9",
			158 => x"05002304",
			159 => x"000602a9",
			160 => x"ff6c02a9",
			161 => x"08001f04",
			162 => x"005a02a9",
			163 => x"0c001d08",
			164 => x"02012504",
			165 => x"000802a9",
			166 => x"ffaa02a9",
			167 => x"09002604",
			168 => x"003602a9",
			169 => x"fff502a9",
			170 => x"0f009d14",
			171 => x"0d001208",
			172 => x"0f007d04",
			173 => x"fe63032d",
			174 => x"02f3032d",
			175 => x"09001e08",
			176 => x"0a003204",
			177 => x"fe60032d",
			178 => x"008a032d",
			179 => x"fe5d032d",
			180 => x"01001028",
			181 => x"0d001720",
			182 => x"03001f04",
			183 => x"03ca032d",
			184 => x"0d00120c",
			185 => x"05002304",
			186 => x"00ab032d",
			187 => x"09001804",
			188 => x"ffe1032d",
			189 => x"fe32032d",
			190 => x"0e008108",
			191 => x"04002104",
			192 => x"07ab032d",
			193 => x"fffd032d",
			194 => x"09001b04",
			195 => x"fe67032d",
			196 => x"01ba032d",
			197 => x"00012404",
			198 => x"0152032d",
			199 => x"0886032d",
			200 => x"04001e04",
			201 => x"ffa8032d",
			202 => x"fe5b032d",
			203 => x"0d001428",
			204 => x"00012720",
			205 => x"05002714",
			206 => x"0300210c",
			207 => x"0e006a04",
			208 => x"ff9103d1",
			209 => x"0000e904",
			210 => x"ffed03d1",
			211 => x"00fd03d1",
			212 => x"07002804",
			213 => x"fffd03d1",
			214 => x"fee303d1",
			215 => x"03002a08",
			216 => x"06006c04",
			217 => x"ffed03d1",
			218 => x"00f403d1",
			219 => x"ff7103d1",
			220 => x"03002304",
			221 => x"ffe603d1",
			222 => x"feab03d1",
			223 => x"02010f0c",
			224 => x"07002d08",
			225 => x"0e006e04",
			226 => x"ff1c03d1",
			227 => x"00a703d1",
			228 => x"fed203d1",
			229 => x"0e008104",
			230 => x"010503d1",
			231 => x"00012d0c",
			232 => x"0d001a04",
			233 => x"ff0303d1",
			234 => x"0600a304",
			235 => x"001e03d1",
			236 => x"fff003d1",
			237 => x"03002604",
			238 => x"011703d1",
			239 => x"09001e04",
			240 => x"fed003d1",
			241 => x"0c001904",
			242 => x"ffb703d1",
			243 => x"00b603d1",
			244 => x"0a00230c",
			245 => x"07002504",
			246 => x"ff260445",
			247 => x"0000e904",
			248 => x"ff8a0445",
			249 => x"015c0445",
			250 => x"08001604",
			251 => x"fec50445",
			252 => x"08001914",
			253 => x"0c001508",
			254 => x"09001904",
			255 => x"001e0445",
			256 => x"016d0445",
			257 => x"07002e08",
			258 => x"03002204",
			259 => x"002b0445",
			260 => x"fea40445",
			261 => x"01150445",
			262 => x"0c001404",
			263 => x"febb0445",
			264 => x"0a003810",
			265 => x"0b001908",
			266 => x"0f00c304",
			267 => x"00370445",
			268 => x"ff6f0445",
			269 => x"0d001a04",
			270 => x"01050445",
			271 => x"ff4a0445",
			272 => x"fed60445",
			273 => x"0f009d14",
			274 => x"0f009810",
			275 => x"09001e0c",
			276 => x"08001d04",
			277 => x"c6d304c9",
			278 => x"00008304",
			279 => x"c6e504c9",
			280 => x"ccfd04c9",
			281 => x"c6d204c9",
			282 => x"c89504c9",
			283 => x"0a002504",
			284 => x"f13204c9",
			285 => x"0300240c",
			286 => x"04001704",
			287 => x"c89504c9",
			288 => x"0a002a04",
			289 => x"e1ea04c9",
			290 => x"cf0f04c9",
			291 => x"08002018",
			292 => x"0c00180c",
			293 => x"03002a08",
			294 => x"0b001504",
			295 => x"c8c704c9",
			296 => x"ceec04c9",
			297 => x"c6d704c9",
			298 => x"0600b008",
			299 => x"0b001804",
			300 => x"d2a804c9",
			301 => x"c6f204c9",
			302 => x"df0804c9",
			303 => x"01001004",
			304 => x"c89504c9",
			305 => x"c6d304c9",
			306 => x"01000e40",
			307 => x"05002414",
			308 => x"0a00230c",
			309 => x"06009508",
			310 => x"01000904",
			311 => x"ffd0056d",
			312 => x"0002056d",
			313 => x"0055056d",
			314 => x"07002e04",
			315 => x"ff90056d",
			316 => x"0002056d",
			317 => x"04001808",
			318 => x"08001c04",
			319 => x"ffa7056d",
			320 => x"001d056d",
			321 => x"04002110",
			322 => x"0f00d60c",
			323 => x"0d001608",
			324 => x"01000704",
			325 => x"0006056d",
			326 => x"0086056d",
			327 => x"ffea056d",
			328 => x"ffe3056d",
			329 => x"0d001810",
			330 => x"0c001908",
			331 => x"04002d04",
			332 => x"ff7f056d",
			333 => x"0009056d",
			334 => x"0b001804",
			335 => x"0037056d",
			336 => x"ffdd056d",
			337 => x"003b056d",
			338 => x"0c001d0c",
			339 => x"03002408",
			340 => x"03002104",
			341 => x"ffee056d",
			342 => x"0012056d",
			343 => x"ff7c056d",
			344 => x"09002404",
			345 => x"0039056d",
			346 => x"ffde056d",
			347 => x"0f00b52c",
			348 => x"0a002f20",
			349 => x"0c00150c",
			350 => x"07002808",
			351 => x"07002404",
			352 => x"ffa70639",
			353 => x"009a0639",
			354 => x"ffb10639",
			355 => x"05002d0c",
			356 => x"03001e08",
			357 => x"03001d04",
			358 => x"ffe20639",
			359 => x"00140639",
			360 => x"ff110639",
			361 => x"03002904",
			362 => x"00250639",
			363 => x"ffc80639",
			364 => x"01000b04",
			365 => x"ff710639",
			366 => x"09002004",
			367 => x"00ba0639",
			368 => x"ffe90639",
			369 => x"01000a18",
			370 => x"04001808",
			371 => x"05002304",
			372 => x"006d0639",
			373 => x"ff480639",
			374 => x"01000504",
			375 => x"ffd80639",
			376 => x"02012104",
			377 => x"ffd20639",
			378 => x"0d001104",
			379 => x"ffe60639",
			380 => x"00f60639",
			381 => x"04001a08",
			382 => x"0c001504",
			383 => x"ffb20639",
			384 => x"00c30639",
			385 => x"04002610",
			386 => x"08001c04",
			387 => x"00280639",
			388 => x"0b001904",
			389 => x"ff050639",
			390 => x"02012704",
			391 => x"00570639",
			392 => x"ffb90639",
			393 => x"09002408",
			394 => x"0600ad04",
			395 => x"000c0639",
			396 => x"009a0639",
			397 => x"ffd80639",
			398 => x"0b001934",
			399 => x"0700322c",
			400 => x"02013724",
			401 => x"0e008718",
			402 => x"0e008210",
			403 => x"0b001608",
			404 => x"04001e04",
			405 => x"002d06dd",
			406 => x"ff4606dd",
			407 => x"05003804",
			408 => x"00ae06dd",
			409 => x"ff9406dd",
			410 => x"0600a704",
			411 => x"fefd06dd",
			412 => x"ffda06dd",
			413 => x"01000904",
			414 => x"fff706dd",
			415 => x"02012804",
			416 => x"000206dd",
			417 => x"011306dd",
			418 => x"0c001504",
			419 => x"ffda06dd",
			420 => x"ff1406dd",
			421 => x"00014a04",
			422 => x"fee106dd",
			423 => x"005406dd",
			424 => x"0d001a18",
			425 => x"0a003610",
			426 => x"0900240c",
			427 => x"09001e04",
			428 => x"ffe406dd",
			429 => x"0000f504",
			430 => x"fff406dd",
			431 => x"012306dd",
			432 => x"ffe206dd",
			433 => x"07003804",
			434 => x"ff7306dd",
			435 => x"007a06dd",
			436 => x"01000c04",
			437 => x"001c06dd",
			438 => x"ff6706dd",
			439 => x"0f009214",
			440 => x"09001e10",
			441 => x"0c001a0c",
			442 => x"0000be04",
			443 => x"fe650751",
			444 => x"0a002d04",
			445 => x"01070751",
			446 => x"fe970751",
			447 => x"02630751",
			448 => x"fe630751",
			449 => x"01001224",
			450 => x"06008804",
			451 => x"04c30751",
			452 => x"0000f904",
			453 => x"fe4b0751",
			454 => x"03002d10",
			455 => x"09001908",
			456 => x"00012704",
			457 => x"01560751",
			458 => x"fe350751",
			459 => x"01000704",
			460 => x"00550751",
			461 => x"022f0751",
			462 => x"00013a04",
			463 => x"fe5c0751",
			464 => x"0b001704",
			465 => x"fe640751",
			466 => x"01f90751",
			467 => x"fe640751",
			468 => x"0f006904",
			469 => x"fe7007a5",
			470 => x"05003f24",
			471 => x"01001220",
			472 => x"0600890c",
			473 => x"07002a08",
			474 => x"01000704",
			475 => x"043407a5",
			476 => x"021507a5",
			477 => x"fe8507a5",
			478 => x"0b001910",
			479 => x"07003208",
			480 => x"02013704",
			481 => x"009607a5",
			482 => x"fe4d07a5",
			483 => x"02013704",
			484 => x"fe4f07a5",
			485 => x"007507a5",
			486 => x"01b207a5",
			487 => x"fe7507a5",
			488 => x"fe6c07a5",
			489 => x"0f009810",
			490 => x"09001e0c",
			491 => x"08001d04",
			492 => x"fe5e0831",
			493 => x"0f004d04",
			494 => x"fe720831",
			495 => x"03b00831",
			496 => x"fe5c0831",
			497 => x"01001234",
			498 => x"03002414",
			499 => x"0000e904",
			500 => x"fe500831",
			501 => x"09001908",
			502 => x"0a002704",
			503 => x"043c0831",
			504 => x"fe5c0831",
			505 => x"04001704",
			506 => x"04430831",
			507 => x"08300831",
			508 => x"0d00140c",
			509 => x"01000b08",
			510 => x"05002504",
			511 => x"001e0831",
			512 => x"fe5c0831",
			513 => x"04bf0831",
			514 => x"00013b08",
			515 => x"07002f04",
			516 => x"07a90831",
			517 => x"fe570831",
			518 => x"0b001504",
			519 => x"fe800831",
			520 => x"08002004",
			521 => x"0a7e0831",
			522 => x"01bd0831",
			523 => x"fe5a0831",
			524 => x"04002e40",
			525 => x"0b001928",
			526 => x"0500351c",
			527 => x"09001f18",
			528 => x"0d001710",
			529 => x"00012708",
			530 => x"04002104",
			531 => x"007a08b5",
			532 => x"feec08b5",
			533 => x"0600af04",
			534 => x"ff2408b5",
			535 => x"003708b5",
			536 => x"0000e704",
			537 => x"ff8308b5",
			538 => x"00ec08b5",
			539 => x"fe8008b5",
			540 => x"0c001804",
			541 => x"fed508b5",
			542 => x"08001f04",
			543 => x"01c208b5",
			544 => x"ff2c08b5",
			545 => x"0a00360c",
			546 => x"09002408",
			547 => x"0f00c004",
			548 => x"ff5508b5",
			549 => x"01dc08b5",
			550 => x"fee708b5",
			551 => x"0c001d04",
			552 => x"fe8f08b5",
			553 => x"0c001e04",
			554 => x"010508b5",
			555 => x"ff8408b5",
			556 => x"fe9c08b5",
			557 => x"0f00be44",
			558 => x"07002a1c",
			559 => x"00011114",
			560 => x"04001e08",
			561 => x"0000be04",
			562 => x"ffbc0991",
			563 => x"00ca0991",
			564 => x"0c001a04",
			565 => x"ff8d0991",
			566 => x"0200a104",
			567 => x"fffa0991",
			568 => x"00310991",
			569 => x"0e007904",
			570 => x"ff590991",
			571 => x"00230991",
			572 => x"0400200c",
			573 => x"03001e08",
			574 => x"03001c04",
			575 => x"fffc0991",
			576 => x"000e0991",
			577 => x"fef30991",
			578 => x"02010b10",
			579 => x"0b001704",
			580 => x"ff900991",
			581 => x"01000e04",
			582 => x"ffe30991",
			583 => x"01001004",
			584 => x"001b0991",
			585 => x"fffb0991",
			586 => x"02011304",
			587 => x"009b0991",
			588 => x"04002804",
			589 => x"ff860991",
			590 => x"00150991",
			591 => x"0f00c30c",
			592 => x"04002108",
			593 => x"09001a04",
			594 => x"ffe00991",
			595 => x"00cd0991",
			596 => x"ff9a0991",
			597 => x"09001f10",
			598 => x"0300270c",
			599 => x"0f00cb04",
			600 => x"ff650991",
			601 => x"01000904",
			602 => x"ffd20991",
			603 => x"009d0991",
			604 => x"ff180991",
			605 => x"01001004",
			606 => x"00aa0991",
			607 => x"00013204",
			608 => x"001b0991",
			609 => x"02014804",
			610 => x"ff8e0991",
			611 => x"00110991",
			612 => x"0f00b53c",
			613 => x"05002820",
			614 => x"07002814",
			615 => x"0500240c",
			616 => x"04001308",
			617 => x"05001c04",
			618 => x"ffe10a75",
			619 => x"00360a75",
			620 => x"ff7b0a75",
			621 => x"0c001504",
			622 => x"00730a75",
			623 => x"ffe00a75",
			624 => x"0a002108",
			625 => x"04001304",
			626 => x"fff90a75",
			627 => x"00150a75",
			628 => x"ff140a75",
			629 => x"04002110",
			630 => x"0b001404",
			631 => x"ffc80a75",
			632 => x"0f009d08",
			633 => x"05002a04",
			634 => x"00330a75",
			635 => x"ffb90a75",
			636 => x"00c80a75",
			637 => x"0e005608",
			638 => x"0200a104",
			639 => x"ffe30a75",
			640 => x"00380a75",
			641 => x"ff5a0a75",
			642 => x"0d001728",
			643 => x"02011c08",
			644 => x"07002f04",
			645 => x"00d60a75",
			646 => x"ff7c0a75",
			647 => x"0600a910",
			648 => x"0100080c",
			649 => x"08001804",
			650 => x"ff830a75",
			651 => x"01000704",
			652 => x"fff40a75",
			653 => x"006c0a75",
			654 => x"ff120a75",
			655 => x"02013308",
			656 => x"0e009504",
			657 => x"009f0a75",
			658 => x"ffbd0a75",
			659 => x"07003004",
			660 => x"ff480a75",
			661 => x"00500a75",
			662 => x"05002c04",
			663 => x"00e40a75",
			664 => x"04002604",
			665 => x"ff4b0a75",
			666 => x"09002404",
			667 => x"00af0a75",
			668 => x"ffd50a75",
			669 => x"04001a24",
			670 => x"03002118",
			671 => x"07002504",
			672 => x"ff490b49",
			673 => x"08001c08",
			674 => x"0000e904",
			675 => x"ffe20b49",
			676 => x"011e0b49",
			677 => x"03001c08",
			678 => x"0a001b04",
			679 => x"ffef0b49",
			680 => x"00370b49",
			681 => x"ffc20b49",
			682 => x"0c001508",
			683 => x"09001904",
			684 => x"ff190b49",
			685 => x"00850b49",
			686 => x"fe9c0b49",
			687 => x"0a002818",
			688 => x"01000c10",
			689 => x"09001d0c",
			690 => x"05002404",
			691 => x"ffd00b49",
			692 => x"06006c04",
			693 => x"ffe50b49",
			694 => x"01460b49",
			695 => x"ff970b49",
			696 => x"0b001704",
			697 => x"ff4d0b49",
			698 => x"00690b49",
			699 => x"05002a0c",
			700 => x"0b001404",
			701 => x"00380b49",
			702 => x"0b001804",
			703 => x"fea60b49",
			704 => x"00810b49",
			705 => x"0a003614",
			706 => x"0d001408",
			707 => x"01000a04",
			708 => x"fed70b49",
			709 => x"00910b49",
			710 => x"01000a04",
			711 => x"01250b49",
			712 => x"07002f04",
			713 => x"007f0b49",
			714 => x"ff760b49",
			715 => x"08001908",
			716 => x"01000804",
			717 => x"ffbf0b49",
			718 => x"00930b49",
			719 => x"0f00e104",
			720 => x"feda0b49",
			721 => x"00350b49",
			722 => x"0a003440",
			723 => x"0c00192c",
			724 => x"04002128",
			725 => x"05002a10",
			726 => x"04001e0c",
			727 => x"0a002c08",
			728 => x"0b001704",
			729 => x"006f0bed",
			730 => x"ff380bed",
			731 => x"ff170bed",
			732 => x"fece0bed",
			733 => x"0f00c30c",
			734 => x"07002904",
			735 => x"ff6e0bed",
			736 => x"04002004",
			737 => x"006b0bed",
			738 => x"01360bed",
			739 => x"08001b08",
			740 => x"0e008404",
			741 => x"ffc40bed",
			742 => x"00b60bed",
			743 => x"ff060bed",
			744 => x"fed10bed",
			745 => x"0a00310c",
			746 => x"07003204",
			747 => x"ff2a0bed",
			748 => x"08002404",
			749 => x"00de0bed",
			750 => x"ffb10bed",
			751 => x"01001004",
			752 => x"01300bed",
			753 => x"ffc80bed",
			754 => x"04002904",
			755 => x"ff090bed",
			756 => x"04002e0c",
			757 => x"07002e04",
			758 => x"ffd40bed",
			759 => x"01001404",
			760 => x"00af0bed",
			761 => x"fff10bed",
			762 => x"ff640bed",
			763 => x"05002a40",
			764 => x"0a002828",
			765 => x"0f00b520",
			766 => x"0c00150c",
			767 => x"07002404",
			768 => x"ffc20cd9",
			769 => x"07002804",
			770 => x"007d0cd9",
			771 => x"ffe70cd9",
			772 => x"07002408",
			773 => x"00009b04",
			774 => x"fff80cd9",
			775 => x"00270cd9",
			776 => x"0a001c08",
			777 => x"03001a04",
			778 => x"fff90cd9",
			779 => x"000a0cd9",
			780 => x"ff6a0cd9",
			781 => x"04001704",
			782 => x"000b0cd9",
			783 => x"008d0cd9",
			784 => x"01000d0c",
			785 => x"05002208",
			786 => x"0b001504",
			787 => x"000b0cd9",
			788 => x"ffea0cd9",
			789 => x"ff240cd9",
			790 => x"03002604",
			791 => x"ffbf0cd9",
			792 => x"03002c04",
			793 => x"002e0cd9",
			794 => x"fffb0cd9",
			795 => x"0a003424",
			796 => x"0b001610",
			797 => x"01000b08",
			798 => x"0000f304",
			799 => x"00160cd9",
			800 => x"ff770cd9",
			801 => x"0a002d04",
			802 => x"ffc20cd9",
			803 => x"007a0cd9",
			804 => x"01000a04",
			805 => x"00e20cd9",
			806 => x"0b001704",
			807 => x"ffb10cd9",
			808 => x"07002f04",
			809 => x"006d0cd9",
			810 => x"0e009104",
			811 => x"ff9d0cd9",
			812 => x"00430cd9",
			813 => x"0c001d0c",
			814 => x"04002d04",
			815 => x"ff640cd9",
			816 => x"04003104",
			817 => x"001b0cd9",
			818 => x"ffd40cd9",
			819 => x"09002504",
			820 => x"00600cd9",
			821 => x"ffea0cd9",
			822 => x"0b001944",
			823 => x"09001d2c",
			824 => x"07003020",
			825 => x"0001371c",
			826 => x"0f00b510",
			827 => x"05002d08",
			828 => x"0c001504",
			829 => x"001d0d95",
			830 => x"ff180d95",
			831 => x"07002904",
			832 => x"ff840d95",
			833 => x"00dc0d95",
			834 => x"00012804",
			835 => x"01020d95",
			836 => x"0a002c04",
			837 => x"005f0d95",
			838 => x"ff5a0d95",
			839 => x"fed10d95",
			840 => x"03002708",
			841 => x"0600ac04",
			842 => x"fff50d95",
			843 => x"01110d95",
			844 => x"ff720d95",
			845 => x"05003308",
			846 => x"08001904",
			847 => x"00870d95",
			848 => x"feb00d95",
			849 => x"05003f0c",
			850 => x"01001008",
			851 => x"09001f04",
			852 => x"00bc0d95",
			853 => x"002c0d95",
			854 => x"ffc80d95",
			855 => x"ffa40d95",
			856 => x"09002418",
			857 => x"0a003608",
			858 => x"0f00c004",
			859 => x"ffe10d95",
			860 => x"00ff0d95",
			861 => x"01000c08",
			862 => x"01000a04",
			863 => x"fff50d95",
			864 => x"00610d95",
			865 => x"08002004",
			866 => x"fff90d95",
			867 => x"ff930d95",
			868 => x"ff7e0d95",
			869 => x"0000e50c",
			870 => x"07002708",
			871 => x"0e005504",
			872 => x"fe800e21",
			873 => x"01060e21",
			874 => x"fe740e21",
			875 => x"0200dc04",
			876 => x"04140e21",
			877 => x"01000e20",
			878 => x"0d001818",
			879 => x"0001270c",
			880 => x"07002f08",
			881 => x"01000b04",
			882 => x"007c0e21",
			883 => x"01dd0e21",
			884 => x"fe7b0e21",
			885 => x"0e008004",
			886 => x"fe5a0e21",
			887 => x"01000c04",
			888 => x"00b20e21",
			889 => x"fee70e21",
			890 => x"0200fa04",
			891 => x"ff360e21",
			892 => x"02420e21",
			893 => x"0300290c",
			894 => x"00012304",
			895 => x"ff410e21",
			896 => x"05002c04",
			897 => x"01570e21",
			898 => x"febf0e21",
			899 => x"0c001d04",
			900 => x"fe540e21",
			901 => x"0b001c04",
			902 => x"01bb0e21",
			903 => x"fe9a0e21",
			904 => x"0f00b634",
			905 => x"0e007c24",
			906 => x"0e007518",
			907 => x"00010714",
			908 => x"09001b08",
			909 => x"0f008c04",
			910 => x"ff890f05",
			911 => x"00dd0f05",
			912 => x"0e005908",
			913 => x"06006004",
			914 => x"ff740f05",
			915 => x"00990f05",
			916 => x"fefe0f05",
			917 => x"fee30f05",
			918 => x"01000c08",
			919 => x"01000704",
			920 => x"ffad0f05",
			921 => x"012c0f05",
			922 => x"ffc80f05",
			923 => x"01000d08",
			924 => x"04001804",
			925 => x"00060f05",
			926 => x"feb20f05",
			927 => x"02010f04",
			928 => x"ffd40f05",
			929 => x"00970f05",
			930 => x"0d001418",
			931 => x"0001270c",
			932 => x"0f00bb04",
			933 => x"ffcb0f05",
			934 => x"07002e04",
			935 => x"01340f05",
			936 => x"ffa30f05",
			937 => x"0f00cc04",
			938 => x"feb10f05",
			939 => x"0f00db04",
			940 => x"00cb0f05",
			941 => x"ff0f0f05",
			942 => x"01000c0c",
			943 => x"04001d04",
			944 => x"00470f05",
			945 => x"01000a04",
			946 => x"01610f05",
			947 => x"001e0f05",
			948 => x"0a002c04",
			949 => x"00cd0f05",
			950 => x"0e009008",
			951 => x"0f00ba04",
			952 => x"ffd10f05",
			953 => x"feba0f05",
			954 => x"04002608",
			955 => x"03002904",
			956 => x"006a0f05",
			957 => x"ff3c0f05",
			958 => x"0b001b04",
			959 => x"00e90f05",
			960 => x"ffb70f05",
			961 => x"0f00b638",
			962 => x"0e007c28",
			963 => x"05002710",
			964 => x"0e00750c",
			965 => x"04001008",
			966 => x"05001b04",
			967 => x"ffb20fe9",
			968 => x"00360fe9",
			969 => x"fec80fe9",
			970 => x"00100fe9",
			971 => x"04002314",
			972 => x"0d00160c",
			973 => x"05002f08",
			974 => x"0000be04",
			975 => x"ffc70fe9",
			976 => x"01260fe9",
			977 => x"ffd90fe9",
			978 => x"05002d04",
			979 => x"ff660fe9",
			980 => x"004f0fe9",
			981 => x"ff070fe9",
			982 => x"01000d08",
			983 => x"04001804",
			984 => x"000b0fe9",
			985 => x"fea60fe9",
			986 => x"02010f04",
			987 => x"ffc40fe9",
			988 => x"00c10fe9",
			989 => x"01000a14",
			990 => x"0d001410",
			991 => x"0300270c",
			992 => x"0600af08",
			993 => x"00012804",
			994 => x"00f70fe9",
			995 => x"fec10fe9",
			996 => x"00d70fe9",
			997 => x"fecf0fe9",
			998 => x"00e00fe9",
			999 => x"0b001918",
			1000 => x"01000d10",
			1001 => x"08001f0c",
			1002 => x"02010a04",
			1003 => x"00130fe9",
			1004 => x"02013804",
			1005 => x"fea40fe9",
			1006 => x"ff810fe9",
			1007 => x"00020fe9",
			1008 => x"08001f04",
			1009 => x"00d00fe9",
			1010 => x"fef50fe9",
			1011 => x"0d001a04",
			1012 => x"00be0fe9",
			1013 => x"00012708",
			1014 => x"0f00bd04",
			1015 => x"fff60fe9",
			1016 => x"00250fe9",
			1017 => x"ff350fe9",
			1018 => x"06009e2c",
			1019 => x"02010c24",
			1020 => x"07002d20",
			1021 => x"0e00751c",
			1022 => x"0c00150c",
			1023 => x"0a002808",
			1024 => x"0200a104",
			1025 => x"ffe510a5",
			1026 => x"006a10a5",
			1027 => x"ffcf10a5",
			1028 => x"0e005908",
			1029 => x"0f006804",
			1030 => x"ffd510a5",
			1031 => x"003c10a5",
			1032 => x"05002d04",
			1033 => x"ff8910a5",
			1034 => x"fffb10a5",
			1035 => x"007c10a5",
			1036 => x"ff9410a5",
			1037 => x"04002704",
			1038 => x"ff5f10a5",
			1039 => x"003b10a5",
			1040 => x"0d001414",
			1041 => x"00012808",
			1042 => x"00011304",
			1043 => x"ffda10a5",
			1044 => x"007010a5",
			1045 => x"0600af04",
			1046 => x"ff4810a5",
			1047 => x"0f00da04",
			1048 => x"006310a5",
			1049 => x"ffbe10a5",
			1050 => x"01000c08",
			1051 => x"0e009204",
			1052 => x"00b810a5",
			1053 => x"000d10a5",
			1054 => x"01000d04",
			1055 => x"ff9310a5",
			1056 => x"0201370c",
			1057 => x"0600b508",
			1058 => x"0a003604",
			1059 => x"007b10a5",
			1060 => x"ffe610a5",
			1061 => x"ffcf10a5",
			1062 => x"0f00e204",
			1063 => x"ffa210a5",
			1064 => x"002710a5",
			1065 => x"0a002824",
			1066 => x"05002410",
			1067 => x"0300210c",
			1068 => x"07002504",
			1069 => x"ff8b1191",
			1070 => x"0000e904",
			1071 => x"ffce1191",
			1072 => x"00db1191",
			1073 => x"ff291191",
			1074 => x"03002610",
			1075 => x"01000c0c",
			1076 => x"04001e08",
			1077 => x"04001a04",
			1078 => x"002b1191",
			1079 => x"01021191",
			1080 => x"ffee1191",
			1081 => x"ffd11191",
			1082 => x"ffa61191",
			1083 => x"0b001728",
			1084 => x"01000b14",
			1085 => x"0000f208",
			1086 => x"0f009d04",
			1087 => x"ffc91191",
			1088 => x"004a1191",
			1089 => x"0b001608",
			1090 => x"01000504",
			1091 => x"ffe51191",
			1092 => x"fed91191",
			1093 => x"ffe11191",
			1094 => x"0b001404",
			1095 => x"ff761191",
			1096 => x"0d001508",
			1097 => x"07002f04",
			1098 => x"00e61191",
			1099 => x"ffce1191",
			1100 => x"04001b04",
			1101 => x"00521191",
			1102 => x"ff661191",
			1103 => x"0a003418",
			1104 => x"05002904",
			1105 => x"ff881191",
			1106 => x"0d001908",
			1107 => x"06006104",
			1108 => x"fff81191",
			1109 => x"00b21191",
			1110 => x"0f00d404",
			1111 => x"ffb51191",
			1112 => x"0e00a204",
			1113 => x"001c1191",
			1114 => x"fffc1191",
			1115 => x"0c001d0c",
			1116 => x"08001908",
			1117 => x"01000804",
			1118 => x"fff01191",
			1119 => x"00441191",
			1120 => x"ff431191",
			1121 => x"0b001b04",
			1122 => x"006f1191",
			1123 => x"ffda1191",
			1124 => x"0d001748",
			1125 => x"0a00230c",
			1126 => x"07002504",
			1127 => x"ffc71255",
			1128 => x"0000e904",
			1129 => x"fff41255",
			1130 => x"00921255",
			1131 => x"0c001930",
			1132 => x"08001b18",
			1133 => x"0d00120c",
			1134 => x"0f00cc08",
			1135 => x"0000e904",
			1136 => x"00201255",
			1137 => x"ff581255",
			1138 => x"00401255",
			1139 => x"05002e08",
			1140 => x"08001804",
			1141 => x"ffe91255",
			1142 => x"00871255",
			1143 => x"ffb21255",
			1144 => x"0001290c",
			1145 => x"05002704",
			1146 => x"ff781255",
			1147 => x"07002f04",
			1148 => x"00701255",
			1149 => x"ffc11255",
			1150 => x"0f00d204",
			1151 => x"ff2a1255",
			1152 => x"0600c104",
			1153 => x"00151255",
			1154 => x"ffd21255",
			1155 => x"05002f04",
			1156 => x"ffca1255",
			1157 => x"04002704",
			1158 => x"00851255",
			1159 => x"ffe71255",
			1160 => x"01000f10",
			1161 => x"0001240c",
			1162 => x"07002b08",
			1163 => x"07002a04",
			1164 => x"fffb1255",
			1165 => x"00101255",
			1166 => x"ffc61255",
			1167 => x"00ae1255",
			1168 => x"03002408",
			1169 => x"09002204",
			1170 => x"003d1255",
			1171 => x"ffe81255",
			1172 => x"ff971255",
			1173 => x"0e006610",
			1174 => x"08001f04",
			1175 => x"fe6c1311",
			1176 => x"08002008",
			1177 => x"0000a804",
			1178 => x"ff441311",
			1179 => x"01561311",
			1180 => x"fea81311",
			1181 => x"0300272c",
			1182 => x"0c001514",
			1183 => x"0a002c10",
			1184 => x"0f00c30c",
			1185 => x"00011108",
			1186 => x"0000d304",
			1187 => x"ff1d1311",
			1188 => x"01f81311",
			1189 => x"ff421311",
			1190 => x"025c1311",
			1191 => x"fea71311",
			1192 => x"00011108",
			1193 => x"04001504",
			1194 => x"002e1311",
			1195 => x"fe341311",
			1196 => x"0d00170c",
			1197 => x"02011904",
			1198 => x"00ed1311",
			1199 => x"07002d04",
			1200 => x"fe561311",
			1201 => x"003e1311",
			1202 => x"01e31311",
			1203 => x"0b001608",
			1204 => x"0000f304",
			1205 => x"012a1311",
			1206 => x"fe5b1311",
			1207 => x"07002f08",
			1208 => x"05003904",
			1209 => x"016f1311",
			1210 => x"fea61311",
			1211 => x"08001c04",
			1212 => x"010a1311",
			1213 => x"0b001a08",
			1214 => x"09002204",
			1215 => x"fe581311",
			1216 => x"ff2f1311",
			1217 => x"09002404",
			1218 => x"01821311",
			1219 => x"fe961311",
			1220 => x"0b00194c",
			1221 => x"0a002308",
			1222 => x"0e006a04",
			1223 => x"ffce13cd",
			1224 => x"007213cd",
			1225 => x"0e008224",
			1226 => x"0500270c",
			1227 => x"0d001408",
			1228 => x"03002104",
			1229 => x"000e13cd",
			1230 => x"ff8113cd",
			1231 => x"001513cd",
			1232 => x"0400210c",
			1233 => x"0f00c308",
			1234 => x"05002f04",
			1235 => x"006313cd",
			1236 => x"ffe913cd",
			1237 => x"ffde13cd",
			1238 => x"05003404",
			1239 => x"ff9c13cd",
			1240 => x"01000b04",
			1241 => x"ffd313cd",
			1242 => x"003c13cd",
			1243 => x"0d00130c",
			1244 => x"0f00cc04",
			1245 => x"ffa913cd",
			1246 => x"03002704",
			1247 => x"005d13cd",
			1248 => x"ffe213cd",
			1249 => x"0500330c",
			1250 => x"01000d04",
			1251 => x"ff4813cd",
			1252 => x"0f00d104",
			1253 => x"002213cd",
			1254 => x"ffd613cd",
			1255 => x"0c001904",
			1256 => x"ffbd13cd",
			1257 => x"004413cd",
			1258 => x"09002410",
			1259 => x"0a003608",
			1260 => x"0f00c004",
			1261 => x"fff513cd",
			1262 => x"008d13cd",
			1263 => x"01000c04",
			1264 => x"001413cd",
			1265 => x"ffd913cd",
			1266 => x"ffcf13cd",
			1267 => x"0000e50c",
			1268 => x"0f006904",
			1269 => x"fe671471",
			1270 => x"0e005a04",
			1271 => x"02dc1471",
			1272 => x"fe651471",
			1273 => x"03002720",
			1274 => x"0d00171c",
			1275 => x"00011908",
			1276 => x"0a002804",
			1277 => x"02581471",
			1278 => x"006e1471",
			1279 => x"0e007b04",
			1280 => x"fe2d1471",
			1281 => x"0600af08",
			1282 => x"00013504",
			1283 => x"011f1471",
			1284 => x"fe221471",
			1285 => x"0f00da04",
			1286 => x"027d1471",
			1287 => x"fe931471",
			1288 => x"02c21471",
			1289 => x"09002424",
			1290 => x"0b001710",
			1291 => x"0001270c",
			1292 => x"0a003108",
			1293 => x"0b001404",
			1294 => x"fe6f1471",
			1295 => x"01fb1471",
			1296 => x"fe691471",
			1297 => x"fe4c1471",
			1298 => x"0100100c",
			1299 => x"0a003404",
			1300 => x"01f81471",
			1301 => x"0d001704",
			1302 => x"fe521471",
			1303 => x"015f1471",
			1304 => x"04002804",
			1305 => x"fe691471",
			1306 => x"00d81471",
			1307 => x"fe6a1471",
			1308 => x"0a002828",
			1309 => x"0f00b520",
			1310 => x"07002814",
			1311 => x"07002304",
			1312 => x"ff78154d",
			1313 => x"0c001504",
			1314 => x"00fa154d",
			1315 => x"01000b04",
			1316 => x"ff9b154d",
			1317 => x"08001f04",
			1318 => x"0044154d",
			1319 => x"fffa154d",
			1320 => x"03001e08",
			1321 => x"05001c04",
			1322 => x"fff7154d",
			1323 => x"0034154d",
			1324 => x"ff31154d",
			1325 => x"0d001204",
			1326 => x"ffea154d",
			1327 => x"00f0154d",
			1328 => x"0d001724",
			1329 => x"0500351c",
			1330 => x"00015818",
			1331 => x"01000d10",
			1332 => x"05002508",
			1333 => x"0f00c304",
			1334 => x"ff8c154d",
			1335 => x"0057154d",
			1336 => x"0f00b204",
			1337 => x"fffe154d",
			1338 => x"fee9154d",
			1339 => x"0600a304",
			1340 => x"006e154d",
			1341 => x"ffab154d",
			1342 => x"0077154d",
			1343 => x"05003804",
			1344 => x"00bd154d",
			1345 => x"ff9b154d",
			1346 => x"01000c08",
			1347 => x"0e007b04",
			1348 => x"ffce154d",
			1349 => x"00e9154d",
			1350 => x"05002704",
			1351 => x"0073154d",
			1352 => x"07002e08",
			1353 => x"0000c604",
			1354 => x"fff4154d",
			1355 => x"006b154d",
			1356 => x"0c001e08",
			1357 => x"07003a04",
			1358 => x"ff17154d",
			1359 => x"fff9154d",
			1360 => x"0d001a04",
			1361 => x"0075154d",
			1362 => x"ffdc154d",
			1363 => x"0400215c",
			1364 => x"04001d38",
			1365 => x"0d001728",
			1366 => x"0c001514",
			1367 => x"01000c10",
			1368 => x"09001908",
			1369 => x"0a002304",
			1370 => x"00771629",
			1371 => x"feaf1629",
			1372 => x"08001c04",
			1373 => x"01a41629",
			1374 => x"ff651629",
			1375 => x"fea41629",
			1376 => x"07003410",
			1377 => x"03002108",
			1378 => x"0e007504",
			1379 => x"ff231629",
			1380 => x"01451629",
			1381 => x"01000c04",
			1382 => x"febc1629",
			1383 => x"009f1629",
			1384 => x"00ec1629",
			1385 => x"0d001808",
			1386 => x"08001d04",
			1387 => x"ffcc1629",
			1388 => x"01c71629",
			1389 => x"0c001b04",
			1390 => x"00061629",
			1391 => x"ff4c1629",
			1392 => x"0201311c",
			1393 => x"0b001710",
			1394 => x"09001d0c",
			1395 => x"0a002804",
			1396 => x"01a01629",
			1397 => x"08001804",
			1398 => x"feba1629",
			1399 => x"00b71629",
			1400 => x"fe8a1629",
			1401 => x"07003208",
			1402 => x"09002004",
			1403 => x"018b1629",
			1404 => x"ffc81629",
			1405 => x"ffd61629",
			1406 => x"0b001b04",
			1407 => x"fe961629",
			1408 => x"002e1629",
			1409 => x"09001e04",
			1410 => x"fe6d1629",
			1411 => x"08001d08",
			1412 => x"0e007604",
			1413 => x"fee11629",
			1414 => x"01611629",
			1415 => x"00015304",
			1416 => x"fe7b1629",
			1417 => x"011b1629",
			1418 => x"01000e60",
			1419 => x"0d001438",
			1420 => x"01000920",
			1421 => x"0b001718",
			1422 => x"0a00230c",
			1423 => x"0e007508",
			1424 => x"04001804",
			1425 => x"ffdf1715",
			1426 => x"00051715",
			1427 => x"00291715",
			1428 => x"0200db08",
			1429 => x"0000d204",
			1430 => x"fff41715",
			1431 => x"001b1715",
			1432 => x"ff7a1715",
			1433 => x"04001904",
			1434 => x"002e1715",
			1435 => x"ffdf1715",
			1436 => x"0e008f14",
			1437 => x"0500290c",
			1438 => x"0b001608",
			1439 => x"09001904",
			1440 => x"ffee1715",
			1441 => x"008a1715",
			1442 => x"ffe31715",
			1443 => x"00012704",
			1444 => x"000d1715",
			1445 => x"ffd31715",
			1446 => x"ffca1715",
			1447 => x"01000a10",
			1448 => x"06009c0c",
			1449 => x"0000f208",
			1450 => x"0000dd04",
			1451 => x"fff21715",
			1452 => x"001e1715",
			1453 => x"ffc61715",
			1454 => x"009b1715",
			1455 => x"04002008",
			1456 => x"08001c04",
			1457 => x"00231715",
			1458 => x"ff951715",
			1459 => x"01000b04",
			1460 => x"ffd01715",
			1461 => x"0e008108",
			1462 => x"07002f04",
			1463 => x"00631715",
			1464 => x"ffee1715",
			1465 => x"fff71715",
			1466 => x"02014814",
			1467 => x"04001808",
			1468 => x"04001604",
			1469 => x"fff81715",
			1470 => x"001a1715",
			1471 => x"03002408",
			1472 => x"03002304",
			1473 => x"fff21715",
			1474 => x"000f1715",
			1475 => x"ff7f1715",
			1476 => x"00221715",
			1477 => x"0b001950",
			1478 => x"0a002308",
			1479 => x"0e006a04",
			1480 => x"ffcc17d9",
			1481 => x"007517d9",
			1482 => x"0e008224",
			1483 => x"0500270c",
			1484 => x"0d001408",
			1485 => x"03002104",
			1486 => x"000e17d9",
			1487 => x"ff7917d9",
			1488 => x"001517d9",
			1489 => x"0400210c",
			1490 => x"05002f08",
			1491 => x"0f00c304",
			1492 => x"006817d9",
			1493 => x"ffdd17d9",
			1494 => x"ffe617d9",
			1495 => x"05003404",
			1496 => x"ff9817d9",
			1497 => x"01000b04",
			1498 => x"ffd117d9",
			1499 => x"003d17d9",
			1500 => x"0c001408",
			1501 => x"0600b004",
			1502 => x"004817d9",
			1503 => x"ffde17d9",
			1504 => x"0700300c",
			1505 => x"03002904",
			1506 => x"ff4717d9",
			1507 => x"05003004",
			1508 => x"001117d9",
			1509 => x"fff417d9",
			1510 => x"05002708",
			1511 => x"0e009204",
			1512 => x"006117d9",
			1513 => x"fff817d9",
			1514 => x"0f00c704",
			1515 => x"001b17d9",
			1516 => x"ff9917d9",
			1517 => x"09002410",
			1518 => x"0a003608",
			1519 => x"0f00c004",
			1520 => x"fff517d9",
			1521 => x"009117d9",
			1522 => x"01000c04",
			1523 => x"001517d9",
			1524 => x"ffd817d9",
			1525 => x"ffcd17d9",
			1526 => x"0a003850",
			1527 => x"01000f3c",
			1528 => x"05003530",
			1529 => x"0300271c",
			1530 => x"0b001710",
			1531 => x"0600a108",
			1532 => x"00011904",
			1533 => x"0073187d",
			1534 => x"fec0187d",
			1535 => x"0d001404",
			1536 => x"0064187d",
			1537 => x"01f6187d",
			1538 => x"0d001304",
			1539 => x"0192187d",
			1540 => x"0d001904",
			1541 => x"fe11187d",
			1542 => x"000f187d",
			1543 => x"09001c04",
			1544 => x"fe62187d",
			1545 => x"00012908",
			1546 => x"07002e04",
			1547 => x"01a1187d",
			1548 => x"ff7d187d",
			1549 => x"07003204",
			1550 => x"fe5b187d",
			1551 => x"0078187d",
			1552 => x"05003908",
			1553 => x"08001d04",
			1554 => x"02c6187d",
			1555 => x"00d0187d",
			1556 => x"feb7187d",
			1557 => x"05003c0c",
			1558 => x"05002608",
			1559 => x"0a002704",
			1560 => x"feed187d",
			1561 => x"00e5187d",
			1562 => x"fe6c187d",
			1563 => x"03003304",
			1564 => x"00fe187d",
			1565 => x"ffb6187d",
			1566 => x"fe73187d",
			1567 => x"06009f38",
			1568 => x"0700281c",
			1569 => x"07002304",
			1570 => x"ffc51981",
			1571 => x"0a002810",
			1572 => x"0c001504",
			1573 => x"00611981",
			1574 => x"01000b04",
			1575 => x"ffd91981",
			1576 => x"08001f04",
			1577 => x"00271981",
			1578 => x"fff51981",
			1579 => x"0c001a04",
			1580 => x"ffc51981",
			1581 => x"00161981",
			1582 => x"03002308",
			1583 => x"0e007604",
			1584 => x"ffe61981",
			1585 => x"002a1981",
			1586 => x"0e00800c",
			1587 => x"0c001a04",
			1588 => x"ff4f1981",
			1589 => x"0c001b04",
			1590 => x"000d1981",
			1591 => x"fff71981",
			1592 => x"0e008104",
			1593 => x"000b1981",
			1594 => x"fffb1981",
			1595 => x"0f00da44",
			1596 => x"05002d1c",
			1597 => x"09001908",
			1598 => x"00012a04",
			1599 => x"00011981",
			1600 => x"ffd81981",
			1601 => x"0f00c308",
			1602 => x"0200f704",
			1603 => x"fff81981",
			1604 => x"00ab1981",
			1605 => x"0f00cb08",
			1606 => x"00013404",
			1607 => x"00121981",
			1608 => x"ff9e1981",
			1609 => x"006f1981",
			1610 => x"0c001910",
			1611 => x"0d00180c",
			1612 => x"0c001608",
			1613 => x"0f00c204",
			1614 => x"00171981",
			1615 => x"fff71981",
			1616 => x"ff7b1981",
			1617 => x"00161981",
			1618 => x"0a00360c",
			1619 => x"00013b04",
			1620 => x"ffe01981",
			1621 => x"0b001c04",
			1622 => x"008e1981",
			1623 => x"fffa1981",
			1624 => x"0b001d04",
			1625 => x"ffbf1981",
			1626 => x"04002904",
			1627 => x"00171981",
			1628 => x"fffb1981",
			1629 => x"04002604",
			1630 => x"ffa21981",
			1631 => x"00151981",
			1632 => x"03002444",
			1633 => x"01000714",
			1634 => x"01000204",
			1635 => x"00741a95",
			1636 => x"04001c0c",
			1637 => x"05002208",
			1638 => x"05001f04",
			1639 => x"ffb11a95",
			1640 => x"005b1a95",
			1641 => x"ff1f1a95",
			1642 => x"003b1a95",
			1643 => x"01000a14",
			1644 => x"0400170c",
			1645 => x"04001308",
			1646 => x"07002504",
			1647 => x"ffed1a95",
			1648 => x"00491a95",
			1649 => x"ffb21a95",
			1650 => x"0000f404",
			1651 => x"fff01a95",
			1652 => x"012c1a95",
			1653 => x"0600a218",
			1654 => x"0700280c",
			1655 => x"0c001204",
			1656 => x"ffcd1a95",
			1657 => x"09001c04",
			1658 => x"00961a95",
			1659 => x"ffe91a95",
			1660 => x"03001e08",
			1661 => x"0a001b04",
			1662 => x"fffa1a95",
			1663 => x"001d1a95",
			1664 => x"ff151a95",
			1665 => x"008c1a95",
			1666 => x"0500352c",
			1667 => x"0600af1c",
			1668 => x"02012218",
			1669 => x"0a002f0c",
			1670 => x"0600a108",
			1671 => x"0000f204",
			1672 => x"00511a95",
			1673 => x"fed81a95",
			1674 => x"009c1a95",
			1675 => x"01000b04",
			1676 => x"ff5c1a95",
			1677 => x"0e008104",
			1678 => x"00dd1a95",
			1679 => x"ffb81a95",
			1680 => x"fecd1a95",
			1681 => x"03002704",
			1682 => x"00b41a95",
			1683 => x"04002308",
			1684 => x"0c001d04",
			1685 => x"ff111a95",
			1686 => x"000b1a95",
			1687 => x"00581a95",
			1688 => x"00011d04",
			1689 => x"ff791a95",
			1690 => x"0c001804",
			1691 => x"ffc11a95",
			1692 => x"0201360c",
			1693 => x"03002e04",
			1694 => x"ffe21a95",
			1695 => x"0d001a04",
			1696 => x"01031a95",
			1697 => x"ffed1a95",
			1698 => x"0a003604",
			1699 => x"00421a95",
			1700 => x"ffa21a95",
			1701 => x"07002304",
			1702 => x"feed1b41",
			1703 => x"03002108",
			1704 => x"0000e904",
			1705 => x"ff681b41",
			1706 => x"014a1b41",
			1707 => x"0b00171c",
			1708 => x"05002f10",
			1709 => x"07002804",
			1710 => x"00d81b41",
			1711 => x"0a002704",
			1712 => x"fe9e1b41",
			1713 => x"01000904",
			1714 => x"ff5f1b41",
			1715 => x"006a1b41",
			1716 => x"03003304",
			1717 => x"fea41b41",
			1718 => x"01000a04",
			1719 => x"ff721b41",
			1720 => x"00ce1b41",
			1721 => x"0a003418",
			1722 => x"07002f08",
			1723 => x"06005d04",
			1724 => x"ffe11b41",
			1725 => x"013c1b41",
			1726 => x"00013b08",
			1727 => x"05002804",
			1728 => x"00941b41",
			1729 => x"febb1b41",
			1730 => x"05002f04",
			1731 => x"ffc81b41",
			1732 => x"01421b41",
			1733 => x"0c001d0c",
			1734 => x"08001908",
			1735 => x"01000804",
			1736 => x"ffca1b41",
			1737 => x"00d21b41",
			1738 => x"feb21b41",
			1739 => x"00014304",
			1740 => x"ff981b41",
			1741 => x"01001804",
			1742 => x"00f21b41",
			1743 => x"ffee1b41",
			1744 => x"04002e68",
			1745 => x"05002420",
			1746 => x"0500231c",
			1747 => x"06009510",
			1748 => x"0b00130c",
			1749 => x"0b001104",
			1750 => x"fed01c17",
			1751 => x"01000904",
			1752 => x"ffb51c17",
			1753 => x"01241c17",
			1754 => x"fe9d1c17",
			1755 => x"0e008a08",
			1756 => x"01000704",
			1757 => x"00d61c17",
			1758 => x"01721c17",
			1759 => x"fef81c17",
			1760 => x"fe441c17",
			1761 => x"03002418",
			1762 => x"04001704",
			1763 => x"fe871c17",
			1764 => x"04001e0c",
			1765 => x"04001c08",
			1766 => x"03002204",
			1767 => x"006c1c17",
			1768 => x"015b1c17",
			1769 => x"01e01c17",
			1770 => x"08001d04",
			1771 => x"008b1c17",
			1772 => x"feab1c17",
			1773 => x"08001f1c",
			1774 => x"0b001710",
			1775 => x"01000908",
			1776 => x"07002504",
			1777 => x"01581c17",
			1778 => x"fe621c17",
			1779 => x"07002e04",
			1780 => x"00c41c17",
			1781 => x"ff7f1c17",
			1782 => x"05002e04",
			1783 => x"00071c17",
			1784 => x"0a003404",
			1785 => x"01961c17",
			1786 => x"000e1c17",
			1787 => x"04002608",
			1788 => x"0e005604",
			1789 => x"00f01c17",
			1790 => x"fe6e1c17",
			1791 => x"09002408",
			1792 => x"0c001a04",
			1793 => x"ff521c17",
			1794 => x"01411c17",
			1795 => x"ff2d1c17",
			1796 => x"fea31c17",
			1797 => x"0200f218",
			1798 => x"0c001508",
			1799 => x"0f009804",
			1800 => x"fe6f1c81",
			1801 => x"02541c81",
			1802 => x"07002708",
			1803 => x"0f006704",
			1804 => x"fe671c81",
			1805 => x"02991c81",
			1806 => x"0f00a004",
			1807 => x"fe641c81",
			1808 => x"fe021c81",
			1809 => x"0100121c",
			1810 => x"04002a18",
			1811 => x"0c001a14",
			1812 => x"0600b810",
			1813 => x"04002208",
			1814 => x"04002004",
			1815 => x"01011c81",
			1816 => x"03291c81",
			1817 => x"08001c04",
			1818 => x"01421c81",
			1819 => x"fe431c81",
			1820 => x"fe5f1c81",
			1821 => x"02891c81",
			1822 => x"fe661c81",
			1823 => x"fe661c81",
			1824 => x"0f007d0c",
			1825 => x"0f006904",
			1826 => x"fe6a1cf5",
			1827 => x"0200a204",
			1828 => x"02051cf5",
			1829 => x"fe741cf5",
			1830 => x"01001024",
			1831 => x"03001f08",
			1832 => x"0000e904",
			1833 => x"ff051cf5",
			1834 => x"01ab1cf5",
			1835 => x"0e006704",
			1836 => x"03d81cf5",
			1837 => x"0001180c",
			1838 => x"0e007908",
			1839 => x"09001d04",
			1840 => x"01171cf5",
			1841 => x"fe651cf5",
			1842 => x"fe1e1cf5",
			1843 => x"0e007b04",
			1844 => x"fe391cf5",
			1845 => x"02011904",
			1846 => x"02171cf5",
			1847 => x"00961cf5",
			1848 => x"0f00e208",
			1849 => x"04001e04",
			1850 => x"ffea1cf5",
			1851 => x"fe5a1cf5",
			1852 => x"01171cf5",
			1853 => x"0f009d10",
			1854 => x"09001e0c",
			1855 => x"06006104",
			1856 => x"fe611d79",
			1857 => x"07002704",
			1858 => x"05ef1d79",
			1859 => x"fe6a1d79",
			1860 => x"fe5f1d79",
			1861 => x"0100102c",
			1862 => x"0b001720",
			1863 => x"0a00280c",
			1864 => x"0e007604",
			1865 => x"011e1d79",
			1866 => x"0d001204",
			1867 => x"02991d79",
			1868 => x"03d61d79",
			1869 => x"0e007f08",
			1870 => x"02011904",
			1871 => x"04bf1d79",
			1872 => x"fe601d79",
			1873 => x"01000d08",
			1874 => x"0b001604",
			1875 => x"fe5c1d79",
			1876 => x"00481d79",
			1877 => x"020e1d79",
			1878 => x"02012d08",
			1879 => x"0e008204",
			1880 => x"04801d79",
			1881 => x"fe331d79",
			1882 => x"05a91d79",
			1883 => x"04001e04",
			1884 => x"ffc01d79",
			1885 => x"fe5d1d79",
			1886 => x"0a002828",
			1887 => x"04001a18",
			1888 => x"0c00150c",
			1889 => x"07002504",
			1890 => x"ffe01e3d",
			1891 => x"0000e904",
			1892 => x"fff71e3d",
			1893 => x"004a1e3d",
			1894 => x"03002108",
			1895 => x"05001e04",
			1896 => x"fff51e3d",
			1897 => x"00181e3d",
			1898 => x"ffa21e3d",
			1899 => x"04001e08",
			1900 => x"07002304",
			1901 => x"fff61e3d",
			1902 => x"007f1e3d",
			1903 => x"03002104",
			1904 => x"00091e3d",
			1905 => x"ffd51e3d",
			1906 => x"0b001714",
			1907 => x"02011910",
			1908 => x"00011b0c",
			1909 => x"05002d04",
			1910 => x"ffac1e3d",
			1911 => x"05002f04",
			1912 => x"00381e3d",
			1913 => x"ffd11e3d",
			1914 => x"002d1e3d",
			1915 => x"ff691e3d",
			1916 => x"0a003414",
			1917 => x"05002e0c",
			1918 => x"0e008308",
			1919 => x"0a002c04",
			1920 => x"00301e3d",
			1921 => x"fff51e3d",
			1922 => x"ffc71e3d",
			1923 => x"01000f04",
			1924 => x"00671e3d",
			1925 => x"ffed1e3d",
			1926 => x"0c001d0c",
			1927 => x"08001908",
			1928 => x"01000804",
			1929 => x"fffa1e3d",
			1930 => x"00131e3d",
			1931 => x"ffa51e3d",
			1932 => x"09002504",
			1933 => x"002d1e3d",
			1934 => x"fff31e3d",
			1935 => x"0f009214",
			1936 => x"09001e10",
			1937 => x"08001d04",
			1938 => x"fe731ec1",
			1939 => x"01000e08",
			1940 => x"05001b04",
			1941 => x"fee41ec1",
			1942 => x"02021ec1",
			1943 => x"fe981ec1",
			1944 => x"fe6b1ec1",
			1945 => x"01001024",
			1946 => x"06008904",
			1947 => x"02881ec1",
			1948 => x"0d001714",
			1949 => x"03001f04",
			1950 => x"01651ec1",
			1951 => x"05002a08",
			1952 => x"0c001504",
			1953 => x"00361ec1",
			1954 => x"fed91ec1",
			1955 => x"07002c04",
			1956 => x"fe6b1ec1",
			1957 => x"01071ec1",
			1958 => x"00013708",
			1959 => x"0e008104",
			1960 => x"013c1ec1",
			1961 => x"fe651ec1",
			1962 => x"02291ec1",
			1963 => x"0d001908",
			1964 => x"0b001904",
			1965 => x"fe641ec1",
			1966 => x"01c91ec1",
			1967 => x"fe681ec1",
			1968 => x"0d001420",
			1969 => x"00011918",
			1970 => x"08001b0c",
			1971 => x"0f009204",
			1972 => x"ffdc1f6d",
			1973 => x"07002d04",
			1974 => x"007e1f6d",
			1975 => x"ffec1f6d",
			1976 => x"07002404",
			1977 => x"00161f6d",
			1978 => x"0a002104",
			1979 => x"000a1f6d",
			1980 => x"ffba1f6d",
			1981 => x"07003004",
			1982 => x"ff511f6d",
			1983 => x"00131f6d",
			1984 => x"02012020",
			1985 => x"09001b08",
			1986 => x"04001a04",
			1987 => x"ffee1f6d",
			1988 => x"00421f6d",
			1989 => x"03002904",
			1990 => x"ff771f6d",
			1991 => x"04002108",
			1992 => x"00010704",
			1993 => x"ffe61f6d",
			1994 => x"00511f6d",
			1995 => x"00012404",
			1996 => x"ffb31f6d",
			1997 => x"00012704",
			1998 => x"00131f6d",
			1999 => x"fff71f6d",
			2000 => x"01000c04",
			2001 => x"00751f6d",
			2002 => x"04002608",
			2003 => x"05002c04",
			2004 => x"00131f6d",
			2005 => x"ff991f6d",
			2006 => x"00014304",
			2007 => x"ffe21f6d",
			2008 => x"07003f04",
			2009 => x"004c1f6d",
			2010 => x"fff61f6d",
			2011 => x"01000f2c",
			2012 => x"07002304",
			2013 => x"fe931fe9",
			2014 => x"0a002308",
			2015 => x"0000e904",
			2016 => x"fefd1fe9",
			2017 => x"018f1fe9",
			2018 => x"0a002404",
			2019 => x"fe971fe9",
			2020 => x"02010f10",
			2021 => x"07002508",
			2022 => x"00009b04",
			2023 => x"ffb21fe9",
			2024 => x"01c41fe9",
			2025 => x"0e007d04",
			2026 => x"ffd11fe9",
			2027 => x"fe591fe9",
			2028 => x"09001904",
			2029 => x"fe941fe9",
			2030 => x"02013104",
			2031 => x"00e71fe9",
			2032 => x"00191fe9",
			2033 => x"0500260c",
			2034 => x"07003204",
			2035 => x"ff401fe9",
			2036 => x"0c002504",
			2037 => x"00f61fe9",
			2038 => x"ffb71fe9",
			2039 => x"0f00e204",
			2040 => x"fe7d1fe9",
			2041 => x"00961fe9",
			2042 => x"0000e50c",
			2043 => x"03002f04",
			2044 => x"fe872075",
			2045 => x"04002604",
			2046 => x"01032075",
			2047 => x"fec92075",
			2048 => x"0400170c",
			2049 => x"0e008504",
			2050 => x"004c2075",
			2051 => x"05002204",
			2052 => x"ffc82075",
			2053 => x"fe102075",
			2054 => x"0300240c",
			2055 => x"0d001204",
			2056 => x"ffba2075",
			2057 => x"00012e04",
			2058 => x"00d62075",
			2059 => x"01a92075",
			2060 => x"08001f18",
			2061 => x"04001d08",
			2062 => x"0f00d004",
			2063 => x"fe632075",
			2064 => x"005c2075",
			2065 => x"0d001308",
			2066 => x"0b001304",
			2067 => x"015e2075",
			2068 => x"fe812075",
			2069 => x"0d001504",
			2070 => x"01402075",
			2071 => x"00102075",
			2072 => x"04002604",
			2073 => x"fe662075",
			2074 => x"09002404",
			2075 => x"00ff2075",
			2076 => x"fed32075",
			2077 => x"0c00183c",
			2078 => x"0a002814",
			2079 => x"03002410",
			2080 => x"07002304",
			2081 => x"ffd02129",
			2082 => x"0000f408",
			2083 => x"0e006b04",
			2084 => x"000e2129",
			2085 => x"ffd62129",
			2086 => x"008d2129",
			2087 => x"ffd62129",
			2088 => x"01000d1c",
			2089 => x"0200fd0c",
			2090 => x"0e006f04",
			2091 => x"ffdb2129",
			2092 => x"0e008204",
			2093 => x"002f2129",
			2094 => x"fff92129",
			2095 => x"01000504",
			2096 => x"000a2129",
			2097 => x"05002508",
			2098 => x"05002304",
			2099 => x"ffe32129",
			2100 => x"00052129",
			2101 => x"ff702129",
			2102 => x"01001008",
			2103 => x"0e008f04",
			2104 => x"003e2129",
			2105 => x"ffe52129",
			2106 => x"ffd72129",
			2107 => x"0500290c",
			2108 => x"05002608",
			2109 => x"05002104",
			2110 => x"fff82129",
			2111 => x"001a2129",
			2112 => x"ffc12129",
			2113 => x"05003f10",
			2114 => x"0100110c",
			2115 => x"0a003108",
			2116 => x"0b001904",
			2117 => x"ffeb2129",
			2118 => x"003d2129",
			2119 => x"00832129",
			2120 => x"ffe02129",
			2121 => x"ffd72129",
			2122 => x"0f00ca48",
			2123 => x"03002420",
			2124 => x"05002410",
			2125 => x"0a002108",
			2126 => x"0f009804",
			2127 => x"ffe721f5",
			2128 => x"002f21f5",
			2129 => x"03001e04",
			2130 => x"000721f5",
			2131 => x"ff9c21f5",
			2132 => x"01000a08",
			2133 => x"0000f404",
			2134 => x"fff721f5",
			2135 => x"008321f5",
			2136 => x"04001d04",
			2137 => x"ffd121f5",
			2138 => x"001d21f5",
			2139 => x"00013a20",
			2140 => x"01000b0c",
			2141 => x"0000f208",
			2142 => x"0f009204",
			2143 => x"ffda21f5",
			2144 => x"003221f5",
			2145 => x"ff4a21f5",
			2146 => x"07002f10",
			2147 => x"01000e08",
			2148 => x"08002004",
			2149 => x"006821f5",
			2150 => x"fffb21f5",
			2151 => x"05002e04",
			2152 => x"ffda21f5",
			2153 => x"000b21f5",
			2154 => x"ffb021f5",
			2155 => x"02012f04",
			2156 => x"004221f5",
			2157 => x"ffeb21f5",
			2158 => x"0f00d614",
			2159 => x"0e00960c",
			2160 => x"08002408",
			2161 => x"0600af04",
			2162 => x"fff321f5",
			2163 => x"008621f5",
			2164 => x"ffea21f5",
			2165 => x"03002c04",
			2166 => x"000621f5",
			2167 => x"ffd821f5",
			2168 => x"07003404",
			2169 => x"ffab21f5",
			2170 => x"00015304",
			2171 => x"ffef21f5",
			2172 => x"004a21f5",
			2173 => x"0f009810",
			2174 => x"09001e0c",
			2175 => x"08001d04",
			2176 => x"fe632279",
			2177 => x"0c001604",
			2178 => x"fe772279",
			2179 => x"02bf2279",
			2180 => x"fe612279",
			2181 => x"01001230",
			2182 => x"0a002c14",
			2183 => x"0000e904",
			2184 => x"fe582279",
			2185 => x"0e00910c",
			2186 => x"0d001104",
			2187 => x"00eb2279",
			2188 => x"00012d04",
			2189 => x"024f2279",
			2190 => x"04042279",
			2191 => x"fe5f2279",
			2192 => x"0b00160c",
			2193 => x"01000b04",
			2194 => x"fe5b2279",
			2195 => x"08001c04",
			2196 => x"05892279",
			2197 => x"fe552279",
			2198 => x"07002f04",
			2199 => x"045e2279",
			2200 => x"02012d04",
			2201 => x"fe5c2279",
			2202 => x"0c001a04",
			2203 => x"00a12279",
			2204 => x"03e62279",
			2205 => x"fe602279",
			2206 => x"0f009810",
			2207 => x"09001e0c",
			2208 => x"08001d04",
			2209 => x"fe6c22ed",
			2210 => x"05002804",
			2211 => x"fe8f22ed",
			2212 => x"01cc22ed",
			2213 => x"fe6822ed",
			2214 => x"01001228",
			2215 => x"0a002304",
			2216 => x"01ca22ed",
			2217 => x"09001908",
			2218 => x"05002104",
			2219 => x"ff9b22ed",
			2220 => x"fe3e22ed",
			2221 => x"0001180c",
			2222 => x"07002d04",
			2223 => x"013222ed",
			2224 => x"03002604",
			2225 => x"fdbb22ed",
			2226 => x"fe6022ed",
			2227 => x"03002708",
			2228 => x"04001804",
			2229 => x"005f22ed",
			2230 => x"022822ed",
			2231 => x"02011c04",
			2232 => x"026722ed",
			2233 => x"001c22ed",
			2234 => x"fe6b22ed",
			2235 => x"0000e50c",
			2236 => x"03002f04",
			2237 => x"fe822391",
			2238 => x"04002604",
			2239 => x"01072391",
			2240 => x"fec02391",
			2241 => x"05002718",
			2242 => x"0500230c",
			2243 => x"0e008a08",
			2244 => x"06009f04",
			2245 => x"004e2391",
			2246 => x"01b42391",
			2247 => x"fed22391",
			2248 => x"07003008",
			2249 => x"0c001504",
			2250 => x"00092391",
			2251 => x"fe3c2391",
			2252 => x"01272391",
			2253 => x"08001d1c",
			2254 => x"09001f14",
			2255 => x"0f00c20c",
			2256 => x"05003808",
			2257 => x"02012204",
			2258 => x"01542391",
			2259 => x"000b2391",
			2260 => x"fec12391",
			2261 => x"0600b404",
			2262 => x"fe732391",
			2263 => x"00712391",
			2264 => x"0f009c04",
			2265 => x"ff6b2391",
			2266 => x"01fc2391",
			2267 => x"07002f04",
			2268 => x"00ed2391",
			2269 => x"0f00e20c",
			2270 => x"0c001d04",
			2271 => x"fe5b2391",
			2272 => x"0d001a04",
			2273 => x"01632391",
			2274 => x"fed32391",
			2275 => x"013f2391",
			2276 => x"0f00be40",
			2277 => x"07002a1c",
			2278 => x"00011114",
			2279 => x"0f009210",
			2280 => x"08001d04",
			2281 => x"ff9b2465",
			2282 => x"08002008",
			2283 => x"01000b04",
			2284 => x"ffe82465",
			2285 => x"005d2465",
			2286 => x"ffd12465",
			2287 => x"00a52465",
			2288 => x"0e007904",
			2289 => x"ff5f2465",
			2290 => x"001e2465",
			2291 => x"0400200c",
			2292 => x"03001e08",
			2293 => x"03001c04",
			2294 => x"fffc2465",
			2295 => x"000f2465",
			2296 => x"feff2465",
			2297 => x"02010b0c",
			2298 => x"07002b08",
			2299 => x"01000804",
			2300 => x"fff82465",
			2301 => x"00142465",
			2302 => x"ff892465",
			2303 => x"02011304",
			2304 => x"00942465",
			2305 => x"04002804",
			2306 => x"ff872465",
			2307 => x"00152465",
			2308 => x"0f00c30c",
			2309 => x"04002108",
			2310 => x"09001a04",
			2311 => x"ffe12465",
			2312 => x"00c42465",
			2313 => x"ff9e2465",
			2314 => x"09001f10",
			2315 => x"0300270c",
			2316 => x"0600ac04",
			2317 => x"ff752465",
			2318 => x"0f00da04",
			2319 => x"00772465",
			2320 => x"ffc22465",
			2321 => x"ff202465",
			2322 => x"01001004",
			2323 => x"00a12465",
			2324 => x"00013204",
			2325 => x"001a2465",
			2326 => x"02014804",
			2327 => x"ff922465",
			2328 => x"00102465",
			2329 => x"0f00980c",
			2330 => x"07002708",
			2331 => x"06006104",
			2332 => x"fe7424e1",
			2333 => x"012a24e1",
			2334 => x"fe6c24e1",
			2335 => x"08002430",
			2336 => x"0d00120c",
			2337 => x"0a002304",
			2338 => x"010424e1",
			2339 => x"04001504",
			2340 => x"ffd024e1",
			2341 => x"fe3824e1",
			2342 => x"0e008310",
			2343 => x"0f00c00c",
			2344 => x"07002f08",
			2345 => x"05002a04",
			2346 => x"003f24e1",
			2347 => x"019624e1",
			2348 => x"fe6c24e1",
			2349 => x"027324e1",
			2350 => x"0c001c10",
			2351 => x"08001f08",
			2352 => x"04001704",
			2353 => x"fe8624e1",
			2354 => x"00c924e1",
			2355 => x"05002904",
			2356 => x"00ec24e1",
			2357 => x"fe4b24e1",
			2358 => x"022b24e1",
			2359 => x"fe7024e1",
			2360 => x"04001a24",
			2361 => x"03002118",
			2362 => x"07002504",
			2363 => x"ff3d25ad",
			2364 => x"08001c08",
			2365 => x"0000e904",
			2366 => x"ffe125ad",
			2367 => x"012625ad",
			2368 => x"03001c08",
			2369 => x"03001a04",
			2370 => x"ffee25ad",
			2371 => x"003d25ad",
			2372 => x"ffbd25ad",
			2373 => x"0c001508",
			2374 => x"09001904",
			2375 => x"ff1025ad",
			2376 => x"009625ad",
			2377 => x"fe9425ad",
			2378 => x"0a002814",
			2379 => x"0e007610",
			2380 => x"07002708",
			2381 => x"0d001204",
			2382 => x"00ff25ad",
			2383 => x"ffbc25ad",
			2384 => x"05001d04",
			2385 => x"001c25ad",
			2386 => x"ff1325ad",
			2387 => x"013125ad",
			2388 => x"05002a0c",
			2389 => x"0600af08",
			2390 => x"0a002a04",
			2391 => x"ff9f25ad",
			2392 => x"feb325ad",
			2393 => x"003825ad",
			2394 => x"0a003614",
			2395 => x"0d001408",
			2396 => x"01000a04",
			2397 => x"fecb25ad",
			2398 => x"00a125ad",
			2399 => x"01000a04",
			2400 => x"013125ad",
			2401 => x"07002f04",
			2402 => x"009025ad",
			2403 => x"ff6b25ad",
			2404 => x"08001908",
			2405 => x"01000804",
			2406 => x"ffbb25ad",
			2407 => x"009925ad",
			2408 => x"0f00e104",
			2409 => x"fed025ad",
			2410 => x"003525ad",
			2411 => x"05002a3c",
			2412 => x"0a002828",
			2413 => x"0f00b520",
			2414 => x"0c00150c",
			2415 => x"07002404",
			2416 => x"ffc02691",
			2417 => x"07002804",
			2418 => x"00822691",
			2419 => x"ffe42691",
			2420 => x"07002408",
			2421 => x"00009b04",
			2422 => x"fff82691",
			2423 => x"00292691",
			2424 => x"0a001c08",
			2425 => x"03001a04",
			2426 => x"fff82691",
			2427 => x"000a2691",
			2428 => x"ff642691",
			2429 => x"04001704",
			2430 => x"000c2691",
			2431 => x"00952691",
			2432 => x"01000d0c",
			2433 => x"05002208",
			2434 => x"0b001504",
			2435 => x"000c2691",
			2436 => x"ffea2691",
			2437 => x"ff1a2691",
			2438 => x"01001004",
			2439 => x"001c2691",
			2440 => x"ffc32691",
			2441 => x"0a003424",
			2442 => x"0b001610",
			2443 => x"01000b08",
			2444 => x"0000f304",
			2445 => x"00172691",
			2446 => x"ff702691",
			2447 => x"0a002d04",
			2448 => x"ffbf2691",
			2449 => x"00812691",
			2450 => x"01000a04",
			2451 => x"00eb2691",
			2452 => x"0b001704",
			2453 => x"ffae2691",
			2454 => x"07002f04",
			2455 => x"00712691",
			2456 => x"0e009104",
			2457 => x"ff9a2691",
			2458 => x"00442691",
			2459 => x"0c001d0c",
			2460 => x"04002d04",
			2461 => x"ff5d2691",
			2462 => x"04003104",
			2463 => x"001c2691",
			2464 => x"ffd32691",
			2465 => x"09002504",
			2466 => x"00612691",
			2467 => x"ffea2691",
			2468 => x"0f00b630",
			2469 => x"0e007c20",
			2470 => x"0001101c",
			2471 => x"0e007514",
			2472 => x"0c001508",
			2473 => x"0000d104",
			2474 => x"ffa12765",
			2475 => x"00f92765",
			2476 => x"0000f208",
			2477 => x"0000ed04",
			2478 => x"ff8e2765",
			2479 => x"00962765",
			2480 => x"ff092765",
			2481 => x"0200f704",
			2482 => x"ffc92765",
			2483 => x"01252765",
			2484 => x"ff402765",
			2485 => x"01000d08",
			2486 => x"04001804",
			2487 => x"00082765",
			2488 => x"feba2765",
			2489 => x"02010f04",
			2490 => x"ffd42765",
			2491 => x"00942765",
			2492 => x"0d001418",
			2493 => x"0001270c",
			2494 => x"0f00bb04",
			2495 => x"ffc52765",
			2496 => x"07002e04",
			2497 => x"012a2765",
			2498 => x"ffa92765",
			2499 => x"0f00cc04",
			2500 => x"feb82765",
			2501 => x"0f00db04",
			2502 => x"00b72765",
			2503 => x"ff1a2765",
			2504 => x"01000c0c",
			2505 => x"04001d04",
			2506 => x"003f2765",
			2507 => x"01000a04",
			2508 => x"01592765",
			2509 => x"001a2765",
			2510 => x"03002604",
			2511 => x"00992765",
			2512 => x"07003704",
			2513 => x"fed92765",
			2514 => x"04002608",
			2515 => x"07003a04",
			2516 => x"ff692765",
			2517 => x"00042765",
			2518 => x"0b001b04",
			2519 => x"00e52765",
			2520 => x"ffb92765",
			2521 => x"0e007518",
			2522 => x"01000904",
			2523 => x"ffb12809",
			2524 => x"0e006a0c",
			2525 => x"0e005908",
			2526 => x"0000a804",
			2527 => x"ffe72809",
			2528 => x"002c2809",
			2529 => x"ffc32809",
			2530 => x"0e007004",
			2531 => x"003b2809",
			2532 => x"fff52809",
			2533 => x"0600b730",
			2534 => x"05002308",
			2535 => x"00010804",
			2536 => x"fff72809",
			2537 => x"006e2809",
			2538 => x"04001808",
			2539 => x"0600a504",
			2540 => x"000b2809",
			2541 => x"ffb12809",
			2542 => x"01000c10",
			2543 => x"01000708",
			2544 => x"05003404",
			2545 => x"ffb12809",
			2546 => x"002b2809",
			2547 => x"06009f04",
			2548 => x"00012809",
			2549 => x"00802809",
			2550 => x"02012608",
			2551 => x"0b001604",
			2552 => x"ffe22809",
			2553 => x"00402809",
			2554 => x"0c001e04",
			2555 => x"ff8b2809",
			2556 => x"001c2809",
			2557 => x"07003404",
			2558 => x"ff952809",
			2559 => x"00015304",
			2560 => x"ffe12809",
			2561 => x"00502809",
			2562 => x"08001b28",
			2563 => x"0600940c",
			2564 => x"0c001508",
			2565 => x"05002404",
			2566 => x"ffd428ed",
			2567 => x"002528ed",
			2568 => x"ffb028ed",
			2569 => x"0e008a14",
			2570 => x"02012e10",
			2571 => x"08001604",
			2572 => x"ffe728ed",
			2573 => x"0a002c04",
			2574 => x"009a28ed",
			2575 => x"09001a04",
			2576 => x"ffea28ed",
			2577 => x"001b28ed",
			2578 => x"ffdf28ed",
			2579 => x"0e009304",
			2580 => x"ffa128ed",
			2581 => x"003728ed",
			2582 => x"05002e2c",
			2583 => x"0d00181c",
			2584 => x"03002210",
			2585 => x"0500250c",
			2586 => x"0a002308",
			2587 => x"05001c04",
			2588 => x"fffa28ed",
			2589 => x"001628ed",
			2590 => x"ffb428ed",
			2591 => x"003f28ed",
			2592 => x"0e007008",
			2593 => x"07002404",
			2594 => x"001c28ed",
			2595 => x"fff628ed",
			2596 => x"ff5528ed",
			2597 => x"07002e08",
			2598 => x"07002c04",
			2599 => x"fffa28ed",
			2600 => x"004c28ed",
			2601 => x"05002704",
			2602 => x"000f28ed",
			2603 => x"ffbd28ed",
			2604 => x"0d00150c",
			2605 => x"07002c04",
			2606 => x"ffe328ed",
			2607 => x"0a003704",
			2608 => x"007528ed",
			2609 => x"fff128ed",
			2610 => x"0b001a0c",
			2611 => x"07002e08",
			2612 => x"0f006904",
			2613 => x"fff328ed",
			2614 => x"002528ed",
			2615 => x"ff7528ed",
			2616 => x"09002404",
			2617 => x"006528ed",
			2618 => x"ffe128ed",
			2619 => x"0a002828",
			2620 => x"0f00b520",
			2621 => x"07002814",
			2622 => x"07002304",
			2623 => x"ffaa29c9",
			2624 => x"0c001504",
			2625 => x"00b029c9",
			2626 => x"01000b04",
			2627 => x"ffc329c9",
			2628 => x"08001f04",
			2629 => x"003929c9",
			2630 => x"ffec29c9",
			2631 => x"03001e08",
			2632 => x"05001c04",
			2633 => x"fffa29c9",
			2634 => x"002229c9",
			2635 => x"ff6129c9",
			2636 => x"04001804",
			2637 => x"001629c9",
			2638 => x"00a529c9",
			2639 => x"0b001720",
			2640 => x"01000d18",
			2641 => x"05002508",
			2642 => x"0d001204",
			2643 => x"003229c9",
			2644 => x"ffb129c9",
			2645 => x"03003308",
			2646 => x"01000404",
			2647 => x"fff629c9",
			2648 => x"fef829c9",
			2649 => x"0a003704",
			2650 => x"003329c9",
			2651 => x"ffdf29c9",
			2652 => x"09001c04",
			2653 => x"008129c9",
			2654 => x"ff9a29c9",
			2655 => x"00013b18",
			2656 => x"07002f0c",
			2657 => x"05003508",
			2658 => x"09002004",
			2659 => x"008c29c9",
			2660 => x"fff629c9",
			2661 => x"ffd729c9",
			2662 => x"05003e04",
			2663 => x"ff5429c9",
			2664 => x"04002c04",
			2665 => x"003429c9",
			2666 => x"fff329c9",
			2667 => x"08002004",
			2668 => x"009329c9",
			2669 => x"02013608",
			2670 => x"02013204",
			2671 => x"fff529c9",
			2672 => x"004029c9",
			2673 => x"ff9629c9",
			2674 => x"09001918",
			2675 => x"00011914",
			2676 => x"0c00140c",
			2677 => x"0d001208",
			2678 => x"0000d104",
			2679 => x"ffb92a75",
			2680 => x"010c2a75",
			2681 => x"ff822a75",
			2682 => x"03001d04",
			2683 => x"002a2a75",
			2684 => x"ff1f2a75",
			2685 => x"fed02a75",
			2686 => x"00010714",
			2687 => x"09001b08",
			2688 => x"0000e204",
			2689 => x"ffad2a75",
			2690 => x"01052a75",
			2691 => x"0e005908",
			2692 => x"06006004",
			2693 => x"ff502a75",
			2694 => x"00c02a75",
			2695 => x"feac2a75",
			2696 => x"00010c04",
			2697 => x"01332a75",
			2698 => x"01000a14",
			2699 => x"04001804",
			2700 => x"ff742a75",
			2701 => x"01000708",
			2702 => x"05003304",
			2703 => x"ff7d2a75",
			2704 => x"00eb2a75",
			2705 => x"06009f04",
			2706 => x"00022a75",
			2707 => x"01452a75",
			2708 => x"00011804",
			2709 => x"feca2a75",
			2710 => x"02011c08",
			2711 => x"0b001804",
			2712 => x"00db2a75",
			2713 => x"ff772a75",
			2714 => x"05002c04",
			2715 => x"00a22a75",
			2716 => x"ff472a75",
			2717 => x"04002e2c",
			2718 => x"0000a804",
			2719 => x"fe7c2ad1",
			2720 => x"01001124",
			2721 => x"0b001918",
			2722 => x"0600890c",
			2723 => x"07002a08",
			2724 => x"0d001104",
			2725 => x"02ea2ad1",
			2726 => x"014f2ad1",
			2727 => x"fe962ad1",
			2728 => x"0e007504",
			2729 => x"fec62ad1",
			2730 => x"05003504",
			2731 => x"00122ad1",
			2732 => x"01ab2ad1",
			2733 => x"0a003608",
			2734 => x"0f00bf04",
			2735 => x"ff3a2ad1",
			2736 => x"02282ad1",
			2737 => x"ff8d2ad1",
			2738 => x"fe802ad1",
			2739 => x"fe6f2ad1",
			2740 => x"0f00be3c",
			2741 => x"02011830",
			2742 => x"05002c18",
			2743 => x"08001b10",
			2744 => x"0a00280c",
			2745 => x"0e006604",
			2746 => x"ff212bad",
			2747 => x"0e007604",
			2748 => x"008c2bad",
			2749 => x"01602bad",
			2750 => x"feca2bad",
			2751 => x"0d001204",
			2752 => x"00af2bad",
			2753 => x"fe6b2bad",
			2754 => x"01000b08",
			2755 => x"05002f04",
			2756 => x"00d52bad",
			2757 => x"fe8a2bad",
			2758 => x"07002f0c",
			2759 => x"0a002f04",
			2760 => x"ff242bad",
			2761 => x"09002004",
			2762 => x"01ac2bad",
			2763 => x"ffb02bad",
			2764 => x"feec2bad",
			2765 => x"01000d04",
			2766 => x"fe7a2bad",
			2767 => x"02011c04",
			2768 => x"00c22bad",
			2769 => x"ffb72bad",
			2770 => x"0f00c30c",
			2771 => x"05002f08",
			2772 => x"0c001504",
			2773 => x"ff532bad",
			2774 => x"01af2bad",
			2775 => x"febc2bad",
			2776 => x"0c001a1c",
			2777 => x"0800190c",
			2778 => x"02013108",
			2779 => x"0600a904",
			2780 => x"00362bad",
			2781 => x"01502bad",
			2782 => x"fed22bad",
			2783 => x"0f00ce04",
			2784 => x"fe842bad",
			2785 => x"0f00da08",
			2786 => x"01000c04",
			2787 => x"015c2bad",
			2788 => x"ff9a2bad",
			2789 => x"fea62bad",
			2790 => x"08002408",
			2791 => x"02013904",
			2792 => x"01952bad",
			2793 => x"006c2bad",
			2794 => x"ff022bad",
			2795 => x"0600af48",
			2796 => x"02012638",
			2797 => x"0f00b520",
			2798 => x"0e007c1c",
			2799 => x"0e007510",
			2800 => x"0000f208",
			2801 => x"0f009004",
			2802 => x"ff992c81",
			2803 => x"00aa2c81",
			2804 => x"01000b04",
			2805 => x"ff022c81",
			2806 => x"ffef2c81",
			2807 => x"01000c08",
			2808 => x"03002f04",
			2809 => x"00d92c81",
			2810 => x"ffcb2c81",
			2811 => x"ff922c81",
			2812 => x"fef92c81",
			2813 => x"0e008108",
			2814 => x"0600a004",
			2815 => x"002e2c81",
			2816 => x"011d2c81",
			2817 => x"07002d04",
			2818 => x"ff5a2c81",
			2819 => x"0f00bf04",
			2820 => x"ff8f2c81",
			2821 => x"0600ac04",
			2822 => x"00d52c81",
			2823 => x"fff72c81",
			2824 => x"0800190c",
			2825 => x"03002704",
			2826 => x"ff4d2c81",
			2827 => x"09001a04",
			2828 => x"fff42c81",
			2829 => x"00b72c81",
			2830 => x"fed72c81",
			2831 => x"0f00d614",
			2832 => x"0e00960c",
			2833 => x"01001008",
			2834 => x"01000a04",
			2835 => x"00582c81",
			2836 => x"00f32c81",
			2837 => x"ffa72c81",
			2838 => x"0f00d304",
			2839 => x"ff732c81",
			2840 => x"00192c81",
			2841 => x"07003404",
			2842 => x"ff102c81",
			2843 => x"00015304",
			2844 => x"ffc32c81",
			2845 => x"08002904",
			2846 => x"00d62c81",
			2847 => x"fff72c81",
			2848 => x"0f00be34",
			2849 => x"02011828",
			2850 => x"02010f20",
			2851 => x"07002d1c",
			2852 => x"04002110",
			2853 => x"04001d08",
			2854 => x"08001b04",
			2855 => x"00552d4d",
			2856 => x"fec22d4d",
			2857 => x"0000be04",
			2858 => x"ff812d4d",
			2859 => x"01222d4d",
			2860 => x"0c001a04",
			2861 => x"fe9b2d4d",
			2862 => x"01000c04",
			2863 => x"ffb32d4d",
			2864 => x"00d92d4d",
			2865 => x"fe812d4d",
			2866 => x"0b001604",
			2867 => x"ff852d4d",
			2868 => x"014b2d4d",
			2869 => x"01000d04",
			2870 => x"fe822d4d",
			2871 => x"02011c04",
			2872 => x"00b22d4d",
			2873 => x"ffbb2d4d",
			2874 => x"0f00c30c",
			2875 => x"05002f08",
			2876 => x"0c001504",
			2877 => x"ff612d4d",
			2878 => x"01982d4d",
			2879 => x"fec32d4d",
			2880 => x"0c001a1c",
			2881 => x"0800190c",
			2882 => x"02013108",
			2883 => x"0600a904",
			2884 => x"00392d4d",
			2885 => x"01362d4d",
			2886 => x"feda2d4d",
			2887 => x"0f00ce04",
			2888 => x"fe902d4d",
			2889 => x"0f00da08",
			2890 => x"01000c04",
			2891 => x"014f2d4d",
			2892 => x"ff9e2d4d",
			2893 => x"feb02d4d",
			2894 => x"08002408",
			2895 => x"05003604",
			2896 => x"018c2d4d",
			2897 => x"00662d4d",
			2898 => x"ff0a2d4d",
			2899 => x"0f009814",
			2900 => x"09001e10",
			2901 => x"0c001a0c",
			2902 => x"0000be04",
			2903 => x"fe682dd9",
			2904 => x"07002404",
			2905 => x"02492dd9",
			2906 => x"fe6e2dd9",
			2907 => x"02742dd9",
			2908 => x"fe652dd9",
			2909 => x"01001230",
			2910 => x"03001f04",
			2911 => x"021c2dd9",
			2912 => x"0d001318",
			2913 => x"0c00150c",
			2914 => x"09001908",
			2915 => x"00012704",
			2916 => x"00b62dd9",
			2917 => x"fe522dd9",
			2918 => x"02292dd9",
			2919 => x"0f00ca08",
			2920 => x"03002604",
			2921 => x"fdd42dd9",
			2922 => x"fe6a2dd9",
			2923 => x"ffbb2dd9",
			2924 => x"00010708",
			2925 => x"09001b04",
			2926 => x"006d2dd9",
			2927 => x"fe252dd9",
			2928 => x"0a002a04",
			2929 => x"02922dd9",
			2930 => x"04001e04",
			2931 => x"ff352dd9",
			2932 => x"01882dd9",
			2933 => x"fe672dd9",
			2934 => x"01000a2c",
			2935 => x"09001c24",
			2936 => x"0c001510",
			2937 => x"07002404",
			2938 => x"ffc92ea5",
			2939 => x"0a002c08",
			2940 => x"0000e504",
			2941 => x"fff42ea5",
			2942 => x"008d2ea5",
			2943 => x"ffd62ea5",
			2944 => x"04001d0c",
			2945 => x"03002108",
			2946 => x"0a002104",
			2947 => x"fffd2ea5",
			2948 => x"00142ea5",
			2949 => x"ff442ea5",
			2950 => x"04001f04",
			2951 => x"00552ea5",
			2952 => x"ffb32ea5",
			2953 => x"0f00ac04",
			2954 => x"ffc52ea5",
			2955 => x"00842ea5",
			2956 => x"0500230c",
			2957 => x"0e008a08",
			2958 => x"0e006a04",
			2959 => x"ffec2ea5",
			2960 => x"00532ea5",
			2961 => x"ffe32ea5",
			2962 => x"0c001d28",
			2963 => x"02012620",
			2964 => x"04002010",
			2965 => x"0f00c008",
			2966 => x"07002404",
			2967 => x"001f2ea5",
			2968 => x"ff4d2ea5",
			2969 => x"00012404",
			2970 => x"ffe72ea5",
			2971 => x"004e2ea5",
			2972 => x"0d001508",
			2973 => x"07002c04",
			2974 => x"ffee2ea5",
			2975 => x"007e2ea5",
			2976 => x"07002b04",
			2977 => x"00132ea5",
			2978 => x"ffc32ea5",
			2979 => x"07003a04",
			2980 => x"ff402ea5",
			2981 => x"ffff2ea5",
			2982 => x"09002404",
			2983 => x"00512ea5",
			2984 => x"ffdb2ea5",
			2985 => x"00010f28",
			2986 => x"07002b24",
			2987 => x"0c001408",
			2988 => x"0000b804",
			2989 => x"ff6e2f71",
			2990 => x"013f2f71",
			2991 => x"0d001510",
			2992 => x"08001d08",
			2993 => x"0c001504",
			2994 => x"00062f71",
			2995 => x"fe9f2f71",
			2996 => x"01000b04",
			2997 => x"ff912f71",
			2998 => x"00b82f71",
			2999 => x"05002d04",
			3000 => x"ff212f71",
			3001 => x"04002304",
			3002 => x"01482f71",
			3003 => x"ff9a2f71",
			3004 => x"fe762f71",
			3005 => x"0300271c",
			3006 => x"0d001718",
			3007 => x"02011908",
			3008 => x"0d001204",
			3009 => x"ffe52f71",
			3010 => x"01002f71",
			3011 => x"0c001508",
			3012 => x"09001804",
			3013 => x"ff122f71",
			3014 => x"01252f71",
			3015 => x"07002d04",
			3016 => x"feaa2f71",
			3017 => x"ffcc2f71",
			3018 => x"01732f71",
			3019 => x"03002904",
			3020 => x"fe7e2f71",
			3021 => x"01000e10",
			3022 => x"07002d04",
			3023 => x"fec32f71",
			3024 => x"05002c04",
			3025 => x"fee52f71",
			3026 => x"08001d04",
			3027 => x"013d2f71",
			3028 => x"00302f71",
			3029 => x"04002604",
			3030 => x"fe8c2f71",
			3031 => x"0f00cb04",
			3032 => x"ff602f71",
			3033 => x"07003f04",
			3034 => x"013b2f71",
			3035 => x"ffb82f71",
			3036 => x"0b001630",
			3037 => x"04001e24",
			3038 => x"0a002c20",
			3039 => x"04001d1c",
			3040 => x"01000910",
			3041 => x"0c001508",
			3042 => x"00011104",
			3043 => x"00943035",
			3044 => x"ffaa3035",
			3045 => x"03001e04",
			3046 => x"000e3035",
			3047 => x"ff153035",
			3048 => x"0f00b408",
			3049 => x"08001b04",
			3050 => x"00833035",
			3051 => x"ff463035",
			3052 => x"00ba3035",
			3053 => x"00e43035",
			3054 => x"ff143035",
			3055 => x"0a002d04",
			3056 => x"fef83035",
			3057 => x"01000b04",
			3058 => x"ff303035",
			3059 => x"00713035",
			3060 => x"0e008218",
			3061 => x"05003814",
			3062 => x"0c001704",
			3063 => x"ffb23035",
			3064 => x"07002f08",
			3065 => x"0f006904",
			3066 => x"ffe13035",
			3067 => x"01213035",
			3068 => x"03002404",
			3069 => x"00193035",
			3070 => x"ffaa3035",
			3071 => x"ff8f3035",
			3072 => x"0600a904",
			3073 => x"ff133035",
			3074 => x"01000c04",
			3075 => x"008c3035",
			3076 => x"04002608",
			3077 => x"00013204",
			3078 => x"00253035",
			3079 => x"ff203035",
			3080 => x"00014304",
			3081 => x"ffa73035",
			3082 => x"03003304",
			3083 => x"00a73035",
			3084 => x"ffdf3035",
			3085 => x"0e007524",
			3086 => x"07002718",
			3087 => x"04001810",
			3088 => x"01000904",
			3089 => x"feff30f9",
			3090 => x"03001c08",
			3091 => x"03001704",
			3092 => x"ffd030f9",
			3093 => x"005630f9",
			3094 => x"ffc530f9",
			3095 => x"06006104",
			3096 => x"ff3f30f9",
			3097 => x"010830f9",
			3098 => x"0a002008",
			3099 => x"0a001c04",
			3100 => x"ffc930f9",
			3101 => x"007430f9",
			3102 => x"fe8d30f9",
			3103 => x"08001808",
			3104 => x"00011d04",
			3105 => x"006c30f9",
			3106 => x"fecd30f9",
			3107 => x"00010704",
			3108 => x"fec530f9",
			3109 => x"0e008314",
			3110 => x"07002f0c",
			3111 => x"04002208",
			3112 => x"0d001404",
			3113 => x"004730f9",
			3114 => x"013730f9",
			3115 => x"ffd730f9",
			3116 => x"0d001a04",
			3117 => x"fed430f9",
			3118 => x"002b30f9",
			3119 => x"09001f10",
			3120 => x"01000d08",
			3121 => x"0d001304",
			3122 => x"007730f9",
			3123 => x"fec730f9",
			3124 => x"09001c04",
			3125 => x"013730f9",
			3126 => x"fedd30f9",
			3127 => x"0a003408",
			3128 => x"09002104",
			3129 => x"017630f9",
			3130 => x"ff7630f9",
			3131 => x"04002604",
			3132 => x"febc30f9",
			3133 => x"009a30f9",
			3134 => x"0f00b538",
			3135 => x"07002d34",
			3136 => x"07002c28",
			3137 => x"0300291c",
			3138 => x"05002710",
			3139 => x"07002808",
			3140 => x"0c001504",
			3141 => x"00d931cd",
			3142 => x"fed731cd",
			3143 => x"03001d04",
			3144 => x"003b31cd",
			3145 => x"fe8f31cd",
			3146 => x"09001d08",
			3147 => x"0000be04",
			3148 => x"ff8f31cd",
			3149 => x"014a31cd",
			3150 => x"feeb31cd",
			3151 => x"01000c04",
			3152 => x"fe8331cd",
			3153 => x"0000a804",
			3154 => x"ffc531cd",
			3155 => x"010331cd",
			3156 => x"01000b04",
			3157 => x"ffa831cd",
			3158 => x"08002204",
			3159 => x"018a31cd",
			3160 => x"ffee31cd",
			3161 => x"fe6331cd",
			3162 => x"0400170c",
			3163 => x"05002208",
			3164 => x"0e009104",
			3165 => x"014d31cd",
			3166 => x"fefd31cd",
			3167 => x"fe6431cd",
			3168 => x"0300260c",
			3169 => x"0f00c604",
			3170 => x"01a331cd",
			3171 => x"0600b104",
			3172 => x"ff5431cd",
			3173 => x"015031cd",
			3174 => x"01000e14",
			3175 => x"09001e10",
			3176 => x"08001c08",
			3177 => x"0e008704",
			3178 => x"ff8331cd",
			3179 => x"011931cd",
			3180 => x"00012a04",
			3181 => x"ffc831cd",
			3182 => x"fe8131cd",
			3183 => x"011d31cd",
			3184 => x"02014804",
			3185 => x"fe7e31cd",
			3186 => x"00f431cd",
			3187 => x"06009f34",
			3188 => x"0700281c",
			3189 => x"07002304",
			3190 => x"ffc732c1",
			3191 => x"0a002810",
			3192 => x"0c001504",
			3193 => x"005e32c1",
			3194 => x"01000b04",
			3195 => x"ffda32c1",
			3196 => x"08001f04",
			3197 => x"002632c1",
			3198 => x"fff532c1",
			3199 => x"0c001a04",
			3200 => x"ffc732c1",
			3201 => x"001532c1",
			3202 => x"0300230c",
			3203 => x"01000504",
			3204 => x"002132c1",
			3205 => x"03001e04",
			3206 => x"001932c1",
			3207 => x"ffdb32c1",
			3208 => x"0b001704",
			3209 => x"ff5b32c1",
			3210 => x"0b001804",
			3211 => x"001432c1",
			3212 => x"ffe532c1",
			3213 => x"0f00da40",
			3214 => x"05002d18",
			3215 => x"09001908",
			3216 => x"00012a04",
			3217 => x"000232c1",
			3218 => x"ffd932c1",
			3219 => x"01000704",
			3220 => x"000832c1",
			3221 => x"04001704",
			3222 => x"fff932c1",
			3223 => x"00011b04",
			3224 => x"fffc32c1",
			3225 => x"009c32c1",
			3226 => x"0c001910",
			3227 => x"0d00180c",
			3228 => x"0c001608",
			3229 => x"0f00c204",
			3230 => x"001632c1",
			3231 => x"fff832c1",
			3232 => x"ff8132c1",
			3233 => x"001432c1",
			3234 => x"0a00360c",
			3235 => x"00013b04",
			3236 => x"ffe132c1",
			3237 => x"0b001c04",
			3238 => x"008932c1",
			3239 => x"fffa32c1",
			3240 => x"0b001d04",
			3241 => x"ffc132c1",
			3242 => x"04002904",
			3243 => x"001732c1",
			3244 => x"fffb32c1",
			3245 => x"04002604",
			3246 => x"ffa532c1",
			3247 => x"001532c1",
			3248 => x"04002e34",
			3249 => x"07002304",
			3250 => x"fe85332d",
			3251 => x"0100112c",
			3252 => x"0b001714",
			3253 => x"0a002308",
			3254 => x"0000e904",
			3255 => x"ff17332d",
			3256 => x"0197332d",
			3257 => x"07002504",
			3258 => x"01a7332d",
			3259 => x"01000904",
			3260 => x"ff44332d",
			3261 => x"004b332d",
			3262 => x"07002f0c",
			3263 => x"09001f08",
			3264 => x"06005d04",
			3265 => x"ffcc332d",
			3266 => x"01b5332d",
			3267 => x"fefa332d",
			3268 => x"0f00c508",
			3269 => x"05002704",
			3270 => x"006c332d",
			3271 => x"fe88332d",
			3272 => x"00d2332d",
			3273 => x"fea3332d",
			3274 => x"fe8d332d",
			3275 => x"0a003460",
			3276 => x"05002410",
			3277 => x"0500230c",
			3278 => x"06009504",
			3279 => x"fee93411",
			3280 => x"0e008f04",
			3281 => x"01063411",
			3282 => x"ff4a3411",
			3283 => x"feba3411",
			3284 => x"01000a24",
			3285 => x"0a00280c",
			3286 => x"04001a04",
			3287 => x"001e3411",
			3288 => x"0000c204",
			3289 => x"ffe33411",
			3290 => x"01513411",
			3291 => x"0b001610",
			3292 => x"0c001408",
			3293 => x"0600a504",
			3294 => x"ff8a3411",
			3295 => x"00fb3411",
			3296 => x"0000f204",
			3297 => x"00af3411",
			3298 => x"fecd3411",
			3299 => x"05002b04",
			3300 => x"00423411",
			3301 => x"01453411",
			3302 => x"04002014",
			3303 => x"0f00c008",
			3304 => x"07002504",
			3305 => x"006b3411",
			3306 => x"fe993411",
			3307 => x"03002704",
			3308 => x"00793411",
			3309 => x"09001f04",
			3310 => x"fedd3411",
			3311 => x"007c3411",
			3312 => x"02011c0c",
			3313 => x"0a002f04",
			3314 => x"ff2b3411",
			3315 => x"07002f04",
			3316 => x"01673411",
			3317 => x"ff8e3411",
			3318 => x"0600b604",
			3319 => x"fee13411",
			3320 => x"01001604",
			3321 => x"00e63411",
			3322 => x"ffec3411",
			3323 => x"0c001d0c",
			3324 => x"03003504",
			3325 => x"feb13411",
			3326 => x"0d001804",
			3327 => x"ff853411",
			3328 => x"009e3411",
			3329 => x"09002504",
			3330 => x"00f53411",
			3331 => x"ffa63411",
			3332 => x"09001918",
			3333 => x"00011914",
			3334 => x"0c00140c",
			3335 => x"0a002708",
			3336 => x"0000aa04",
			3337 => x"ffe234f5",
			3338 => x"00ef34f5",
			3339 => x"ff8c34f5",
			3340 => x"03001d04",
			3341 => x"001134f5",
			3342 => x"ff7a34f5",
			3343 => x"ff0f34f5",
			3344 => x"0400212c",
			3345 => x"0f00da28",
			3346 => x"0d001108",
			3347 => x"0a002304",
			3348 => x"001034f5",
			3349 => x"ff5234f5",
			3350 => x"01000c10",
			3351 => x"04001708",
			3352 => x"05002204",
			3353 => x"008534f5",
			3354 => x"ff3834f5",
			3355 => x"02010304",
			3356 => x"001d34f5",
			3357 => x"00c134f5",
			3358 => x"04001808",
			3359 => x"03002404",
			3360 => x"ffda34f5",
			3361 => x"00c334f5",
			3362 => x"0b001704",
			3363 => x"ff2a34f5",
			3364 => x"002e34f5",
			3365 => x"ff4b34f5",
			3366 => x"0500340c",
			3367 => x"0b001904",
			3368 => x"fee834f5",
			3369 => x"0b001c04",
			3370 => x"006b34f5",
			3371 => x"fff234f5",
			3372 => x"01000b0c",
			3373 => x"08001908",
			3374 => x"01000804",
			3375 => x"ffe234f5",
			3376 => x"006234f5",
			3377 => x"ff5034f5",
			3378 => x"0800200c",
			3379 => x"0d001808",
			3380 => x"04003104",
			3381 => x"00db34f5",
			3382 => x"fff934f5",
			3383 => x"ffe834f5",
			3384 => x"0a003608",
			3385 => x"03003104",
			3386 => x"ffe134f5",
			3387 => x"007f34f5",
			3388 => x"ff7534f5",
			3389 => x"0a002308",
			3390 => x"0e006a04",
			3391 => x"ffc535c1",
			3392 => x"007c35c1",
			3393 => x"05002a24",
			3394 => x"0e006c08",
			3395 => x"0d001404",
			3396 => x"004135c1",
			3397 => x"ffe835c1",
			3398 => x"0d001718",
			3399 => x"0c00150c",
			3400 => x"09001904",
			3401 => x"ff9635c1",
			3402 => x"0a002c04",
			3403 => x"005435c1",
			3404 => x"ffdb35c1",
			3405 => x"03002104",
			3406 => x"001735c1",
			3407 => x"09001c04",
			3408 => x"ff5935c1",
			3409 => x"fff235c1",
			3410 => x"001235c1",
			3411 => x"01000a18",
			3412 => x"0d001408",
			3413 => x"00014404",
			3414 => x"ff9035c1",
			3415 => x"000535c1",
			3416 => x"0600980c",
			3417 => x"0000f208",
			3418 => x"0000dd04",
			3419 => x"fff635c1",
			3420 => x"002735c1",
			3421 => x"ffc635c1",
			3422 => x"00be35c1",
			3423 => x"07002f10",
			3424 => x"01000b04",
			3425 => x"ffc435c1",
			3426 => x"00010708",
			3427 => x"05003404",
			3428 => x"ffe135c1",
			3429 => x"001435c1",
			3430 => x"007a35c1",
			3431 => x"0c001d0c",
			3432 => x"0c001704",
			3433 => x"fff335c1",
			3434 => x"07003a04",
			3435 => x"ff4035c1",
			3436 => x"ffff35c1",
			3437 => x"09002504",
			3438 => x"005035c1",
			3439 => x"ffdf35c1",
			3440 => x"04002e3c",
			3441 => x"07002304",
			3442 => x"fe7e363f",
			3443 => x"09002434",
			3444 => x"0b001718",
			3445 => x"0a002308",
			3446 => x"0000e904",
			3447 => x"ff0c363f",
			3448 => x"019d363f",
			3449 => x"01000908",
			3450 => x"00012e04",
			3451 => x"001b363f",
			3452 => x"fe55363f",
			3453 => x"00011d04",
			3454 => x"ffaf363f",
			3455 => x"00d1363f",
			3456 => x"07002f0c",
			3457 => x"09001f08",
			3458 => x"06005d04",
			3459 => x"ffc8363f",
			3460 => x"01d7363f",
			3461 => x"ff0a363f",
			3462 => x"0600a908",
			3463 => x"08002004",
			3464 => x"fe8a363f",
			3465 => x"ff78363f",
			3466 => x"04002304",
			3467 => x"003e363f",
			3468 => x"014e363f",
			3469 => x"fe9d363f",
			3470 => x"fe88363f",
			3471 => x"0f009810",
			3472 => x"09001e0c",
			3473 => x"08001d04",
			3474 => x"fe6f36a1",
			3475 => x"0c001604",
			3476 => x"fe8636a1",
			3477 => x"01a236a1",
			3478 => x"fe6936a1",
			3479 => x"01001220",
			3480 => x"0a002304",
			3481 => x"01b136a1",
			3482 => x"09001908",
			3483 => x"05002104",
			3484 => x"ff9d36a1",
			3485 => x"fe4536a1",
			3486 => x"00011808",
			3487 => x"07002d04",
			3488 => x"010b36a1",
			3489 => x"fe1836a1",
			3490 => x"0b001908",
			3491 => x"08001d04",
			3492 => x"012636a1",
			3493 => x"ff8236a1",
			3494 => x"01ec36a1",
			3495 => x"fe6d36a1",
			3496 => x"0d001428",
			3497 => x"00012720",
			3498 => x"05002714",
			3499 => x"0300210c",
			3500 => x"0e006a04",
			3501 => x"ff8c373d",
			3502 => x"0000e904",
			3503 => x"ffec373d",
			3504 => x"0106373d",
			3505 => x"07002804",
			3506 => x"fff5373d",
			3507 => x"fed8373d",
			3508 => x"03002a08",
			3509 => x"06006c04",
			3510 => x"ffec373d",
			3511 => x"0102373d",
			3512 => x"ff69373d",
			3513 => x"03002304",
			3514 => x"ffea373d",
			3515 => x"fea4373d",
			3516 => x"02010f0c",
			3517 => x"07002d08",
			3518 => x"0e006e04",
			3519 => x"ff13373d",
			3520 => x"00b5373d",
			3521 => x"fec8373d",
			3522 => x"05002c08",
			3523 => x"03002604",
			3524 => x"0115373d",
			3525 => x"fff8373d",
			3526 => x"03002904",
			3527 => x"fee2373d",
			3528 => x"01000c04",
			3529 => x"010c373d",
			3530 => x"0f00b604",
			3531 => x"0104373d",
			3532 => x"07003704",
			3533 => x"fefb373d",
			3534 => x"0058373d",
			3535 => x"06009e20",
			3536 => x"02010c18",
			3537 => x"07002d14",
			3538 => x"0f00920c",
			3539 => x"0c001a04",
			3540 => x"ffa837e1",
			3541 => x"0b001804",
			3542 => x"001f37e1",
			3543 => x"fff437e1",
			3544 => x"03002c04",
			3545 => x"008237e1",
			3546 => x"ffc537e1",
			3547 => x"ff9237e1",
			3548 => x"04002704",
			3549 => x"ff5737e1",
			3550 => x"003b37e1",
			3551 => x"0d001414",
			3552 => x"02011b08",
			3553 => x"00011304",
			3554 => x"ffd937e1",
			3555 => x"007637e1",
			3556 => x"0600af04",
			3557 => x"ff4537e1",
			3558 => x"03002704",
			3559 => x"006a37e1",
			3560 => x"ffbc37e1",
			3561 => x"01000c08",
			3562 => x"0e009204",
			3563 => x"00c137e1",
			3564 => x"000c37e1",
			3565 => x"01000d04",
			3566 => x"ff8e37e1",
			3567 => x"0201370c",
			3568 => x"0600b508",
			3569 => x"0a003604",
			3570 => x"008037e1",
			3571 => x"ffe437e1",
			3572 => x"ffcd37e1",
			3573 => x"0f00e204",
			3574 => x"ff9f37e1",
			3575 => x"002637e1",
			3576 => x"0a002828",
			3577 => x"04001a18",
			3578 => x"0c00150c",
			3579 => x"07002504",
			3580 => x"ffe038a5",
			3581 => x"0000e904",
			3582 => x"fff738a5",
			3583 => x"004838a5",
			3584 => x"03002108",
			3585 => x"05001e04",
			3586 => x"fff538a5",
			3587 => x"001838a5",
			3588 => x"ffa538a5",
			3589 => x"04001e08",
			3590 => x"07002304",
			3591 => x"fff638a5",
			3592 => x"007b38a5",
			3593 => x"03002104",
			3594 => x"000938a5",
			3595 => x"ffd638a5",
			3596 => x"0b001714",
			3597 => x"02011910",
			3598 => x"00011b0c",
			3599 => x"05002d04",
			3600 => x"ffae38a5",
			3601 => x"05002f04",
			3602 => x"003638a5",
			3603 => x"ffd238a5",
			3604 => x"002d38a5",
			3605 => x"ff6f38a5",
			3606 => x"0a003414",
			3607 => x"05002e0c",
			3608 => x"0e008308",
			3609 => x"0a002c04",
			3610 => x"003038a5",
			3611 => x"fff538a5",
			3612 => x"ffc938a5",
			3613 => x"01000f04",
			3614 => x"006438a5",
			3615 => x"ffed38a5",
			3616 => x"0c001d0c",
			3617 => x"08001908",
			3618 => x"01000804",
			3619 => x"fffa38a5",
			3620 => x"001238a5",
			3621 => x"ffa738a5",
			3622 => x"09002504",
			3623 => x"002b38a5",
			3624 => x"fff438a5",
			3625 => x"0b001934",
			3626 => x"0700322c",
			3627 => x"02013724",
			3628 => x"0e008718",
			3629 => x"0e008210",
			3630 => x"0b001608",
			3631 => x"04001e04",
			3632 => x"00303931",
			3633 => x"ff393931",
			3634 => x"05003804",
			3635 => x"00b63931",
			3636 => x"ff8f3931",
			3637 => x"09001a04",
			3638 => x"fffd3931",
			3639 => x"ff083931",
			3640 => x"02012808",
			3641 => x"0600ad04",
			3642 => x"001f3931",
			3643 => x"ffa53931",
			3644 => x"00ef3931",
			3645 => x"0c001504",
			3646 => x"ffd13931",
			3647 => x"ff0a3931",
			3648 => x"00014a04",
			3649 => x"fed63931",
			3650 => x"00593931",
			3651 => x"0d001a0c",
			3652 => x"0a003908",
			3653 => x"0f00c004",
			3654 => x"ffe03931",
			3655 => x"01023931",
			3656 => x"ffaa3931",
			3657 => x"01000c04",
			3658 => x"001c3931",
			3659 => x"ff613931",
			3660 => x"05002a30",
			3661 => x"0c001514",
			3662 => x"00011108",
			3663 => x"0000e504",
			3664 => x"ffc039f5",
			3665 => x"00e739f5",
			3666 => x"0600a504",
			3667 => x"ff4e39f5",
			3668 => x"0e009104",
			3669 => x"00c639f5",
			3670 => x"ff8d39f5",
			3671 => x"03002108",
			3672 => x"0200c504",
			3673 => x"ffc339f5",
			3674 => x"009839f5",
			3675 => x"0f00d510",
			3676 => x"0b001908",
			3677 => x"03002204",
			3678 => x"ff9f39f5",
			3679 => x"fed939f5",
			3680 => x"09002104",
			3681 => x"003a39f5",
			3682 => x"ffe939f5",
			3683 => x"004339f5",
			3684 => x"0b001614",
			3685 => x"05002f10",
			3686 => x"0a002d08",
			3687 => x"07002a04",
			3688 => x"003339f5",
			3689 => x"ff5839f5",
			3690 => x"01000a04",
			3691 => x"ffd039f5",
			3692 => x"00b239f5",
			3693 => x"ff4d39f5",
			3694 => x"01000a08",
			3695 => x"0f00ba04",
			3696 => x"ffac39f5",
			3697 => x"010339f5",
			3698 => x"07002f0c",
			3699 => x"01000b04",
			3700 => x"ffce39f5",
			3701 => x"09001f04",
			3702 => x"00af39f5",
			3703 => x"ffee39f5",
			3704 => x"07003704",
			3705 => x"ff0539f5",
			3706 => x"0d001a04",
			3707 => x"00b339f5",
			3708 => x"ffad39f5",
			3709 => x"0f009214",
			3710 => x"09001e10",
			3711 => x"0c001a0c",
			3712 => x"0000be04",
			3713 => x"fe643a79",
			3714 => x"0a002d04",
			3715 => x"01463a79",
			3716 => x"fe903a79",
			3717 => x"02d83a79",
			3718 => x"fe623a79",
			3719 => x"0100122c",
			3720 => x"03002d20",
			3721 => x"0900190c",
			3722 => x"00012708",
			3723 => x"01000804",
			3724 => x"02543a79",
			3725 => x"ff153a79",
			3726 => x"fe2c3a79",
			3727 => x"0000e904",
			3728 => x"fe6f3a79",
			3729 => x"01000708",
			3730 => x"03002704",
			3731 => x"00f53a79",
			3732 => x"fe623a79",
			3733 => x"07002f04",
			3734 => x"03233a79",
			3735 => x"01563a79",
			3736 => x"00013a04",
			3737 => x"fe583a79",
			3738 => x"0b001704",
			3739 => x"fe5f3a79",
			3740 => x"025d3a79",
			3741 => x"fe623a79",
			3742 => x"0f009210",
			3743 => x"09001e0c",
			3744 => x"08001d04",
			3745 => x"fe693b15",
			3746 => x"0c001604",
			3747 => x"fe7c3b15",
			3748 => x"021b3b15",
			3749 => x"fe663b15",
			3750 => x"0300271c",
			3751 => x"0d001714",
			3752 => x"0f009d04",
			3753 => x"054b3b15",
			3754 => x"08001d0c",
			3755 => x"03002608",
			3756 => x"00012704",
			3757 => x"018a3b15",
			3758 => x"00053b15",
			3759 => x"030a3b15",
			3760 => x"fe5d3b15",
			3761 => x"0d001b04",
			3762 => x"037e3b15",
			3763 => x"fead3b15",
			3764 => x"0800201c",
			3765 => x"0b001710",
			3766 => x"0001270c",
			3767 => x"0a003108",
			3768 => x"05002904",
			3769 => x"fe6d3b15",
			3770 => x"02783b15",
			3771 => x"fe663b15",
			3772 => x"fe473b15",
			3773 => x"0a003d08",
			3774 => x"01000c04",
			3775 => x"02573b15",
			3776 => x"00f83b15",
			3777 => x"fe7e3b15",
			3778 => x"01001004",
			3779 => x"ff983b15",
			3780 => x"fe673b15",
			3781 => x"0e008234",
			3782 => x"0e007514",
			3783 => x"0c001408",
			3784 => x"07002204",
			3785 => x"ffe43bd9",
			3786 => x"00283bd9",
			3787 => x"07002408",
			3788 => x"07002304",
			3789 => x"fff43bd9",
			3790 => x"00103bd9",
			3791 => x"ffa73bd9",
			3792 => x"04002214",
			3793 => x"0c001408",
			3794 => x"00011e04",
			3795 => x"00133bd9",
			3796 => x"ffd03bd9",
			3797 => x"0d001204",
			3798 => x"ffe93bd9",
			3799 => x"07002f04",
			3800 => x"00823bd9",
			3801 => x"ffee3bd9",
			3802 => x"04002d04",
			3803 => x"ffc93bd9",
			3804 => x"0d001804",
			3805 => x"00173bd9",
			3806 => x"fff63bd9",
			3807 => x"09001f14",
			3808 => x"00015810",
			3809 => x"0c001508",
			3810 => x"03002704",
			3811 => x"00363bd9",
			3812 => x"ffe03bd9",
			3813 => x"05002304",
			3814 => x"00193bd9",
			3815 => x"ff5a3bd9",
			3816 => x"001b3bd9",
			3817 => x"01000c04",
			3818 => x"005b3bd9",
			3819 => x"0f00e214",
			3820 => x"0c001e0c",
			3821 => x"02012508",
			3822 => x"02011d04",
			3823 => x"fffb3bd9",
			3824 => x"000b3bd9",
			3825 => x"ffa83bd9",
			3826 => x"09002704",
			3827 => x"00203bd9",
			3828 => x"fff83bd9",
			3829 => x"00223bd9",
			3830 => x"0f00b528",
			3831 => x"05002d18",
			3832 => x"0c00150c",
			3833 => x"07002808",
			3834 => x"07002404",
			3835 => x"ffad3c9d",
			3836 => x"00923c9d",
			3837 => x"ffb53c9d",
			3838 => x"03001e08",
			3839 => x"03001d04",
			3840 => x"ffe33c9d",
			3841 => x"00133c9d",
			3842 => x"ff193c9d",
			3843 => x"01000b08",
			3844 => x"09001b04",
			3845 => x"00333c9d",
			3846 => x"ff623c9d",
			3847 => x"09001e04",
			3848 => x"00aa3c9d",
			3849 => x"ffdc3c9d",
			3850 => x"0e008314",
			3851 => x"05002d0c",
			3852 => x"0d001208",
			3853 => x"0d001004",
			3854 => x"001f3c9d",
			3855 => x"ffb33c9d",
			3856 => x"00e93c9d",
			3857 => x"05003204",
			3858 => x"ff6d3c9d",
			3859 => x"003d3c9d",
			3860 => x"0e008704",
			3861 => x"ff603c9d",
			3862 => x"0001350c",
			3863 => x"0600a708",
			3864 => x"0600a504",
			3865 => x"fff23c9d",
			3866 => x"00463c9d",
			3867 => x"ff6d3c9d",
			3868 => x"0001450c",
			3869 => x"07003204",
			3870 => x"00c53c9d",
			3871 => x"0c001b04",
			3872 => x"ff793c9d",
			3873 => x"00853c9d",
			3874 => x"07003204",
			3875 => x"ff533c9d",
			3876 => x"08002004",
			3877 => x"00763c9d",
			3878 => x"ffba3c9d",
			3879 => x"0f009810",
			3880 => x"09001e0c",
			3881 => x"08001d04",
			3882 => x"fe623d11",
			3883 => x"05002804",
			3884 => x"fe783d11",
			3885 => x"038c3d11",
			3886 => x"fe603d11",
			3887 => x"01001228",
			3888 => x"03001f04",
			3889 => x"03023d11",
			3890 => x"00011808",
			3891 => x"07002b04",
			3892 => x"02773d11",
			3893 => x"fe303d11",
			3894 => x"0d001410",
			3895 => x"00012708",
			3896 => x"06009f04",
			3897 => x"011b3d11",
			3898 => x"04a13d11",
			3899 => x"0600af04",
			3900 => x"fe423d11",
			3901 => x"00c23d11",
			3902 => x"0e008204",
			3903 => x"065e3d11",
			3904 => x"0f00c404",
			3905 => x"fe353d11",
			3906 => x"02f43d11",
			3907 => x"fe5e3d11",
			3908 => x"0f00ca48",
			3909 => x"03002420",
			3910 => x"05002410",
			3911 => x"0a002108",
			3912 => x"0f009804",
			3913 => x"ffe73ddd",
			3914 => x"002e3ddd",
			3915 => x"03001e04",
			3916 => x"00063ddd",
			3917 => x"ff9f3ddd",
			3918 => x"01000a08",
			3919 => x"0000f404",
			3920 => x"fff73ddd",
			3921 => x"007f3ddd",
			3922 => x"04001d04",
			3923 => x"ffd33ddd",
			3924 => x"001d3ddd",
			3925 => x"00013a20",
			3926 => x"01000b0c",
			3927 => x"0000f208",
			3928 => x"0f009204",
			3929 => x"ffdb3ddd",
			3930 => x"00313ddd",
			3931 => x"ff513ddd",
			3932 => x"07002f10",
			3933 => x"01000e08",
			3934 => x"08002004",
			3935 => x"00633ddd",
			3936 => x"fffb3ddd",
			3937 => x"05002e04",
			3938 => x"ffdc3ddd",
			3939 => x"000b3ddd",
			3940 => x"ffb23ddd",
			3941 => x"02012f04",
			3942 => x"00413ddd",
			3943 => x"ffeb3ddd",
			3944 => x"0d001308",
			3945 => x"03002704",
			3946 => x"00683ddd",
			3947 => x"fff73ddd",
			3948 => x"0b001910",
			3949 => x"09001c08",
			3950 => x"01000b04",
			3951 => x"ffe13ddd",
			3952 => x"00403ddd",
			3953 => x"0a003204",
			3954 => x"ff983ddd",
			3955 => x"00033ddd",
			3956 => x"09002404",
			3957 => x"00523ddd",
			3958 => x"ffe43ddd",
			3959 => x"0f00b53c",
			3960 => x"05002820",
			3961 => x"07002814",
			3962 => x"0500240c",
			3963 => x"04001308",
			3964 => x"05001c04",
			3965 => x"ffe23ec1",
			3966 => x"00333ec1",
			3967 => x"ff7f3ec1",
			3968 => x"0c001504",
			3969 => x"006d3ec1",
			3970 => x"ffe13ec1",
			3971 => x"0a002108",
			3972 => x"04001304",
			3973 => x"fff93ec1",
			3974 => x"00143ec1",
			3975 => x"ff1c3ec1",
			3976 => x"04002110",
			3977 => x"0b001404",
			3978 => x"ffc93ec1",
			3979 => x"0f009d08",
			3980 => x"05002a04",
			3981 => x"00313ec1",
			3982 => x"ffbb3ec1",
			3983 => x"00bd3ec1",
			3984 => x"0e005608",
			3985 => x"0200a104",
			3986 => x"ffe43ec1",
			3987 => x"00373ec1",
			3988 => x"ff603ec1",
			3989 => x"0d001724",
			3990 => x"02011c08",
			3991 => x"07002f04",
			3992 => x"00ca3ec1",
			3993 => x"ff803ec1",
			3994 => x"0600a90c",
			3995 => x"07002d08",
			3996 => x"01000504",
			3997 => x"00263ec1",
			3998 => x"ff0d3ec1",
			3999 => x"00163ec1",
			4000 => x"02013308",
			4001 => x"0e008e04",
			4002 => x"00b03ec1",
			4003 => x"ffea3ec1",
			4004 => x"07003004",
			4005 => x"ff4f3ec1",
			4006 => x"004c3ec1",
			4007 => x"04001e04",
			4008 => x"00e03ec1",
			4009 => x"04002608",
			4010 => x"00014b04",
			4011 => x"ff4d3ec1",
			4012 => x"00233ec1",
			4013 => x"09002404",
			4014 => x"00a53ec1",
			4015 => x"ffd73ec1",
			4016 => x"0f009810",
			4017 => x"09001e0c",
			4018 => x"08001d04",
			4019 => x"fe743f45",
			4020 => x"0c001604",
			4021 => x"fe933f45",
			4022 => x"01603f45",
			4023 => x"fe6c3f45",
			4024 => x"08002430",
			4025 => x"0d00120c",
			4026 => x"0a002304",
			4027 => x"011c3f45",
			4028 => x"0f00d004",
			4029 => x"fe2e3f45",
			4030 => x"ffbd3f45",
			4031 => x"0e008310",
			4032 => x"0f00c00c",
			4033 => x"07002f08",
			4034 => x"05003804",
			4035 => x"01283f45",
			4036 => x"fe7e3f45",
			4037 => x"fe673f45",
			4038 => x"02df3f45",
			4039 => x"0c001c10",
			4040 => x"08001f08",
			4041 => x"04001e04",
			4042 => x"ffa23f45",
			4043 => x"01763f45",
			4044 => x"05002904",
			4045 => x"00f93f45",
			4046 => x"fe433f45",
			4047 => x"024a3f45",
			4048 => x"fe6c3f45",
			4049 => x"0e007518",
			4050 => x"01000904",
			4051 => x"ffac3fe9",
			4052 => x"0e006a0c",
			4053 => x"0e005908",
			4054 => x"0000a804",
			4055 => x"ffe73fe9",
			4056 => x"002e3fe9",
			4057 => x"ffc13fe9",
			4058 => x"0e007004",
			4059 => x"003c3fe9",
			4060 => x"fff53fe9",
			4061 => x"0600b730",
			4062 => x"05002308",
			4063 => x"00010804",
			4064 => x"fff63fe9",
			4065 => x"00713fe9",
			4066 => x"0100070c",
			4067 => x"05003408",
			4068 => x"0e007f04",
			4069 => x"000e3fe9",
			4070 => x"ff8e3fe9",
			4071 => x"002c3fe9",
			4072 => x"01000a0c",
			4073 => x"04001a04",
			4074 => x"ffcf3fe9",
			4075 => x"06009f04",
			4076 => x"ffdb3fe9",
			4077 => x"00a13fe9",
			4078 => x"02012608",
			4079 => x"09001b04",
			4080 => x"ffb33fe9",
			4081 => x"00533fe9",
			4082 => x"0e009004",
			4083 => x"ff6d3fe9",
			4084 => x"003b3fe9",
			4085 => x"07003404",
			4086 => x"ff913fe9",
			4087 => x"00015304",
			4088 => x"ffe03fe9",
			4089 => x"00533fe9",
			4090 => x"01000f4c",
			4091 => x"04001720",
			4092 => x"0b001614",
			4093 => x"0e008510",
			4094 => x"0600960c",
			4095 => x"03001c08",
			4096 => x"05001904",
			4097 => x"ff7b40a5",
			4098 => x"009440a5",
			4099 => x"fe9f40a5",
			4100 => x"016140a5",
			4101 => x"fea740a5",
			4102 => x"03002108",
			4103 => x"05001e04",
			4104 => x"ff4940a5",
			4105 => x"00a940a5",
			4106 => x"fe0e40a5",
			4107 => x"0e008718",
			4108 => x"0f00c514",
			4109 => x"0600a510",
			4110 => x"0e008108",
			4111 => x"01000e04",
			4112 => x"006940a5",
			4113 => x"fe8d40a5",
			4114 => x"07002f04",
			4115 => x"fe7040a5",
			4116 => x"ffae40a5",
			4117 => x"01cc40a5",
			4118 => x"fe7c40a5",
			4119 => x"0e008b08",
			4120 => x"01000a04",
			4121 => x"023c40a5",
			4122 => x"006340a5",
			4123 => x"00013c04",
			4124 => x"fe7f40a5",
			4125 => x"0f00d604",
			4126 => x"00f640a5",
			4127 => x"ffda40a5",
			4128 => x"0500260c",
			4129 => x"07003204",
			4130 => x"ff4940a5",
			4131 => x"0c002504",
			4132 => x"00e940a5",
			4133 => x"ffbd40a5",
			4134 => x"0f00e204",
			4135 => x"fe8240a5",
			4136 => x"008d40a5",
			4137 => x"08002044",
			4138 => x"0600af30",
			4139 => x"00013028",
			4140 => x"0f00b518",
			4141 => x"02010210",
			4142 => x"04002108",
			4143 => x"05002504",
			4144 => x"ffac4151",
			4145 => x"00bf4151",
			4146 => x"08001f04",
			4147 => x"ff2d4151",
			4148 => x"00614151",
			4149 => x"04002004",
			4150 => x"ff0c4151",
			4151 => x"000e4151",
			4152 => x"07002f0c",
			4153 => x"0e008308",
			4154 => x"08001804",
			4155 => x"ffdd4151",
			4156 => x"012f4151",
			4157 => x"ffc64151",
			4158 => x"ff444151",
			4159 => x"0b001604",
			4160 => x"fec34151",
			4161 => x"001f4151",
			4162 => x"04001708",
			4163 => x"00013904",
			4164 => x"fff84151",
			4165 => x"ff4e4151",
			4166 => x"00013504",
			4167 => x"ff704151",
			4168 => x"0a002f04",
			4169 => x"01024151",
			4170 => x"00404151",
			4171 => x"0a002c10",
			4172 => x"0100110c",
			4173 => x"0b001904",
			4174 => x"ffc64151",
			4175 => x"00008f04",
			4176 => x"fff94151",
			4177 => x"00c74151",
			4178 => x"ff8f4151",
			4179 => x"feef4151",
			4180 => x"0f006904",
			4181 => x"fe7341cd",
			4182 => x"01000e20",
			4183 => x"04002e1c",
			4184 => x"0d001718",
			4185 => x"0001270c",
			4186 => x"07002f08",
			4187 => x"01000b04",
			4188 => x"00ca41cd",
			4189 => x"022c41cd",
			4190 => x"fe7341cd",
			4191 => x"0e008004",
			4192 => x"fe4841cd",
			4193 => x"0a003404",
			4194 => x"008e41cd",
			4195 => x"fe6b41cd",
			4196 => x"01ba41cd",
			4197 => x"fe7a41cd",
			4198 => x"03002910",
			4199 => x"0c001604",
			4200 => x"fe5b41cd",
			4201 => x"00010a04",
			4202 => x"fe9941cd",
			4203 => x"04002104",
			4204 => x"018441cd",
			4205 => x"fec841cd",
			4206 => x"0c001d04",
			4207 => x"fe4e41cd",
			4208 => x"0d001b04",
			4209 => x"01f841cd",
			4210 => x"fe8d41cd",
			4211 => x"0c00183c",
			4212 => x"0a002814",
			4213 => x"03002410",
			4214 => x"07002304",
			4215 => x"ffd14291",
			4216 => x"0000f408",
			4217 => x"0e006b04",
			4218 => x"000e4291",
			4219 => x"ffd74291",
			4220 => x"00864291",
			4221 => x"ffda4291",
			4222 => x"01000d1c",
			4223 => x"0200fd0c",
			4224 => x"0e006f04",
			4225 => x"ffdc4291",
			4226 => x"0e008204",
			4227 => x"002d4291",
			4228 => x"fff94291",
			4229 => x"01000504",
			4230 => x"00094291",
			4231 => x"05002508",
			4232 => x"05002304",
			4233 => x"ffe44291",
			4234 => x"00044291",
			4235 => x"ff764291",
			4236 => x"01001008",
			4237 => x"0e008f04",
			4238 => x"003a4291",
			4239 => x"ffe54291",
			4240 => x"ffd84291",
			4241 => x"0500290c",
			4242 => x"05002608",
			4243 => x"05002104",
			4244 => x"fff84291",
			4245 => x"00194291",
			4246 => x"ffc34291",
			4247 => x"05003f18",
			4248 => x"01001114",
			4249 => x"00011b0c",
			4250 => x"0000a904",
			4251 => x"00144291",
			4252 => x"0d001704",
			4253 => x"ffe54291",
			4254 => x"000a4291",
			4255 => x"0a003104",
			4256 => x"001a4291",
			4257 => x"00814291",
			4258 => x"ffe14291",
			4259 => x"ffd84291",
			4260 => x"00010f28",
			4261 => x"07002b24",
			4262 => x"0c001408",
			4263 => x"0000b804",
			4264 => x"ff74434d",
			4265 => x"0136434d",
			4266 => x"0d001510",
			4267 => x"08001d08",
			4268 => x"0c001504",
			4269 => x"000a434d",
			4270 => x"fea9434d",
			4271 => x"01000b04",
			4272 => x"ff97434d",
			4273 => x"00b2434d",
			4274 => x"05002d04",
			4275 => x"ff28434d",
			4276 => x"04002304",
			4277 => x"013d434d",
			4278 => x"ff9e434d",
			4279 => x"fe7d434d",
			4280 => x"02012b24",
			4281 => x"07002f1c",
			4282 => x"0e007b08",
			4283 => x"00011e04",
			4284 => x"006a434d",
			4285 => x"fea8434d",
			4286 => x"0e008108",
			4287 => x"06009f04",
			4288 => x"00a7434d",
			4289 => x"0173434d",
			4290 => x"0600a504",
			4291 => x"fed7434d",
			4292 => x"01000804",
			4293 => x"0011434d",
			4294 => x"00c7434d",
			4295 => x"05002704",
			4296 => x"0049434d",
			4297 => x"fe9a434d",
			4298 => x"07003004",
			4299 => x"fe8a434d",
			4300 => x"09001f04",
			4301 => x"ffbe434d",
			4302 => x"01001004",
			4303 => x"00e9434d",
			4304 => x"02014804",
			4305 => x"feff434d",
			4306 => x"004c434d",
			4307 => x"0a002828",
			4308 => x"0f00b520",
			4309 => x"07002814",
			4310 => x"07002304",
			4311 => x"ffae4429",
			4312 => x"0c001504",
			4313 => x"00ab4429",
			4314 => x"01000b04",
			4315 => x"ffc44429",
			4316 => x"08001f04",
			4317 => x"00364429",
			4318 => x"ffed4429",
			4319 => x"03001e08",
			4320 => x"05001c04",
			4321 => x"fffa4429",
			4322 => x"00204429",
			4323 => x"ff674429",
			4324 => x"0e008504",
			4325 => x"009d4429",
			4326 => x"00154429",
			4327 => x"0b001720",
			4328 => x"01000d18",
			4329 => x"05002508",
			4330 => x"03002604",
			4331 => x"ffb54429",
			4332 => x"002e4429",
			4333 => x"03003308",
			4334 => x"01000404",
			4335 => x"fff64429",
			4336 => x"ff074429",
			4337 => x"0a003704",
			4338 => x"00304429",
			4339 => x"ffdf4429",
			4340 => x"09001c04",
			4341 => x"00784429",
			4342 => x"ff9e4429",
			4343 => x"00013b18",
			4344 => x"07002f0c",
			4345 => x"05003508",
			4346 => x"09002004",
			4347 => x"00864429",
			4348 => x"fff74429",
			4349 => x"ffd84429",
			4350 => x"05003e04",
			4351 => x"ff5d4429",
			4352 => x"04002c04",
			4353 => x"00324429",
			4354 => x"fff44429",
			4355 => x"08002004",
			4356 => x"008b4429",
			4357 => x"02013608",
			4358 => x"02013204",
			4359 => x"fff54429",
			4360 => x"003e4429",
			4361 => x"ff994429",
			4362 => x"01000e4c",
			4363 => x"04001818",
			4364 => x"0a002308",
			4365 => x"06008e04",
			4366 => x"ffc544ed",
			4367 => x"007944ed",
			4368 => x"01000c0c",
			4369 => x"0b001304",
			4370 => x"fffe44ed",
			4371 => x"04001304",
			4372 => x"001744ed",
			4373 => x"ff2544ed",
			4374 => x"002f44ed",
			4375 => x"01000714",
			4376 => x"0a002a08",
			4377 => x"01000404",
			4378 => x"005544ed",
			4379 => x"ffc844ed",
			4380 => x"0d001308",
			4381 => x"0b001704",
			4382 => x"ffaa44ed",
			4383 => x"004c44ed",
			4384 => x"ff6544ed",
			4385 => x"0f00d71c",
			4386 => x"0e00800c",
			4387 => x"00011e08",
			4388 => x"0d001604",
			4389 => x"008244ed",
			4390 => x"ff9744ed",
			4391 => x"ff8b44ed",
			4392 => x"0d001408",
			4393 => x"0c001404",
			4394 => x"005144ed",
			4395 => x"ffc544ed",
			4396 => x"01000c04",
			4397 => x"00e944ed",
			4398 => x"ffea44ed",
			4399 => x"ffb544ed",
			4400 => x"03002608",
			4401 => x"00012304",
			4402 => x"ffa344ed",
			4403 => x"005544ed",
			4404 => x"0201480c",
			4405 => x"07002b08",
			4406 => x"00009404",
			4407 => x"fffa44ed",
			4408 => x"000644ed",
			4409 => x"ff3e44ed",
			4410 => x"002b44ed",
			4411 => x"0d001430",
			4412 => x"0a002710",
			4413 => x"07002304",
			4414 => x"ffba45b9",
			4415 => x"0000be04",
			4416 => x"ffe345b9",
			4417 => x"0a002304",
			4418 => x"009c45b9",
			4419 => x"002945b9",
			4420 => x"01000d1c",
			4421 => x"09001c14",
			4422 => x"0b001410",
			4423 => x"0600af08",
			4424 => x"0e006e04",
			4425 => x"001b45b9",
			4426 => x"ff9045b9",
			4427 => x"00013904",
			4428 => x"005545b9",
			4429 => x"ffc645b9",
			4430 => x"ff1b45b9",
			4431 => x"03002704",
			4432 => x"006345b9",
			4433 => x"ffb945b9",
			4434 => x"003b45b9",
			4435 => x"02010f18",
			4436 => x"05002a04",
			4437 => x"ff7b45b9",
			4438 => x"05002f08",
			4439 => x"0000d504",
			4440 => x"ffea45b9",
			4441 => x"007345b9",
			4442 => x"07002708",
			4443 => x"00009504",
			4444 => x"fff345b9",
			4445 => x"002245b9",
			4446 => x"ff9a45b9",
			4447 => x"01000c08",
			4448 => x"0b001704",
			4449 => x"00a145b9",
			4450 => x"002e45b9",
			4451 => x"05002c04",
			4452 => x"004445b9",
			4453 => x"04002608",
			4454 => x"0f00bc04",
			4455 => x"000345b9",
			4456 => x"ff5a45b9",
			4457 => x"05003504",
			4458 => x"ffcc45b9",
			4459 => x"0d001a04",
			4460 => x"007545b9",
			4461 => x"ffe845b9",
			4462 => x"0e007524",
			4463 => x"07002718",
			4464 => x"04001810",
			4465 => x"01000904",
			4466 => x"ff084675",
			4467 => x"03001c08",
			4468 => x"03001704",
			4469 => x"ffd24675",
			4470 => x"00524675",
			4471 => x"ffc64675",
			4472 => x"06006104",
			4473 => x"ff484675",
			4474 => x"00fc4675",
			4475 => x"0a002008",
			4476 => x"0a001c04",
			4477 => x"ffcc4675",
			4478 => x"00764675",
			4479 => x"fe934675",
			4480 => x"0800180c",
			4481 => x"00011d04",
			4482 => x"00694675",
			4483 => x"02011d04",
			4484 => x"ffa24675",
			4485 => x"fec34675",
			4486 => x"00010704",
			4487 => x"fed14675",
			4488 => x"0e008210",
			4489 => x"07002f0c",
			4490 => x"02010f04",
			4491 => x"00234675",
			4492 => x"0d001404",
			4493 => x"000b4675",
			4494 => x"014f4675",
			4495 => x"ff024675",
			4496 => x"09001f0c",
			4497 => x"0a002a04",
			4498 => x"00824675",
			4499 => x"0a002d04",
			4500 => x"fe854675",
			4501 => x"ffde4675",
			4502 => x"0a003408",
			4503 => x"09002104",
			4504 => x"016c4675",
			4505 => x"ff774675",
			4506 => x"04002604",
			4507 => x"fec74675",
			4508 => x"008a4675",
			4509 => x"0a002824",
			4510 => x"05002410",
			4511 => x"0300210c",
			4512 => x"07002504",
			4513 => x"ff864761",
			4514 => x"0000e904",
			4515 => x"ffcd4761",
			4516 => x"00e54761",
			4517 => x"ff1d4761",
			4518 => x"03002610",
			4519 => x"01000c0c",
			4520 => x"04001e08",
			4521 => x"06006c04",
			4522 => x"fff34761",
			4523 => x"00f64761",
			4524 => x"ffec4761",
			4525 => x"ffce4761",
			4526 => x"ffa24761",
			4527 => x"0b001728",
			4528 => x"01000b14",
			4529 => x"0000f208",
			4530 => x"0f009d04",
			4531 => x"ffc64761",
			4532 => x"004f4761",
			4533 => x"0b001608",
			4534 => x"01000504",
			4535 => x"ffe24761",
			4536 => x"fed04761",
			4537 => x"ffe04761",
			4538 => x"0b001404",
			4539 => x"ff704761",
			4540 => x"0d001508",
			4541 => x"07002f04",
			4542 => x"00f14761",
			4543 => x"ffcb4761",
			4544 => x"04001b04",
			4545 => x"00524761",
			4546 => x"ff604761",
			4547 => x"0a003418",
			4548 => x"05002904",
			4549 => x"ff814761",
			4550 => x"0d001908",
			4551 => x"06006104",
			4552 => x"fff84761",
			4553 => x"00be4761",
			4554 => x"0f00d404",
			4555 => x"ffb24761",
			4556 => x"0e00a204",
			4557 => x"001d4761",
			4558 => x"fffc4761",
			4559 => x"0c001d0c",
			4560 => x"08001908",
			4561 => x"01000804",
			4562 => x"fff04761",
			4563 => x"00464761",
			4564 => x"ff3a4761",
			4565 => x"0b001b04",
			4566 => x"00764761",
			4567 => x"ffd94761",
			4568 => x"01000e50",
			4569 => x"04001820",
			4570 => x"0a002308",
			4571 => x"06008e04",
			4572 => x"ffc3482d",
			4573 => x"007d482d",
			4574 => x"01000c14",
			4575 => x"0500220c",
			4576 => x"0e008c08",
			4577 => x"0b001504",
			4578 => x"0034482d",
			4579 => x"fff9482d",
			4580 => x"ffd0482d",
			4581 => x"0f00a804",
			4582 => x"001e482d",
			4583 => x"ff1d482d",
			4584 => x"002d482d",
			4585 => x"01000714",
			4586 => x"0a002a08",
			4587 => x"01000404",
			4588 => x"005a482d",
			4589 => x"ffc6482d",
			4590 => x"0d001308",
			4591 => x"0b001704",
			4592 => x"ffa8482d",
			4593 => x"004f482d",
			4594 => x"ff5e482d",
			4595 => x"0f00d718",
			4596 => x"0e00800c",
			4597 => x"00011e08",
			4598 => x"0d001604",
			4599 => x"008b482d",
			4600 => x"ff93482d",
			4601 => x"ff87482d",
			4602 => x"0a002d04",
			4603 => x"00da482d",
			4604 => x"05002e04",
			4605 => x"ffba482d",
			4606 => x"0052482d",
			4607 => x"ffb1482d",
			4608 => x"04001808",
			4609 => x"04001604",
			4610 => x"fff4482d",
			4611 => x"004a482d",
			4612 => x"0201480c",
			4613 => x"03002408",
			4614 => x"03002204",
			4615 => x"ffe1482d",
			4616 => x"0021482d",
			4617 => x"ff47482d",
			4618 => x"002c482d",
			4619 => x"0e006610",
			4620 => x"08001f04",
			4621 => x"fe6848e9",
			4622 => x"08002008",
			4623 => x"0000a804",
			4624 => x"ff3648e9",
			4625 => x"017c48e9",
			4626 => x"fe9f48e9",
			4627 => x"0300272c",
			4628 => x"0c001514",
			4629 => x"0a002c10",
			4630 => x"0f00c30c",
			4631 => x"00011108",
			4632 => x"0000d304",
			4633 => x"ff1448e9",
			4634 => x"020d48e9",
			4635 => x"ff2f48e9",
			4636 => x"029748e9",
			4637 => x"fea048e9",
			4638 => x"00011108",
			4639 => x"04001504",
			4640 => x"002748e9",
			4641 => x"fe2a48e9",
			4642 => x"0d00170c",
			4643 => x"02011904",
			4644 => x"010448e9",
			4645 => x"07002d04",
			4646 => x"fe4048e9",
			4647 => x"004b48e9",
			4648 => x"021848e9",
			4649 => x"0b001608",
			4650 => x"0000f304",
			4651 => x"014748e9",
			4652 => x"fe5748e9",
			4653 => x"07002f08",
			4654 => x"05003904",
			4655 => x"018d48e9",
			4656 => x"fe9d48e9",
			4657 => x"08001c04",
			4658 => x"012148e9",
			4659 => x"0b001a08",
			4660 => x"09002204",
			4661 => x"fe5048e9",
			4662 => x"ff2b48e9",
			4663 => x"09002404",
			4664 => x"019b48e9",
			4665 => x"fe9048e9",
			4666 => x"0f007d04",
			4667 => x"fe7e495d",
			4668 => x"0100102c",
			4669 => x"0a003928",
			4670 => x"05003520",
			4671 => x"03002710",
			4672 => x"0c001508",
			4673 => x"0a002c04",
			4674 => x"013c495d",
			4675 => x"feb1495d",
			4676 => x"00011104",
			4677 => x"fee3495d",
			4678 => x"0064495d",
			4679 => x"0c001808",
			4680 => x"00010804",
			4681 => x"ffd7495d",
			4682 => x"fe68495d",
			4683 => x"01000c04",
			4684 => x"0096495d",
			4685 => x"ffc6495d",
			4686 => x"0c001804",
			4687 => x"fed7495d",
			4688 => x"01a1495d",
			4689 => x"fe86495d",
			4690 => x"0c001b04",
			4691 => x"fe73495d",
			4692 => x"09002404",
			4693 => x"00e8495d",
			4694 => x"fea5495d",
			4695 => x"0d00174c",
			4696 => x"0a00230c",
			4697 => x"07002504",
			4698 => x"ffc94a29",
			4699 => x"0000e904",
			4700 => x"fff44a29",
			4701 => x"008c4a29",
			4702 => x"0c001934",
			4703 => x"08001b1c",
			4704 => x"03002710",
			4705 => x"09001908",
			4706 => x"0000ed04",
			4707 => x"00234a29",
			4708 => x"ff984a29",
			4709 => x"0d001104",
			4710 => x"ffe54a29",
			4711 => x"006e4a29",
			4712 => x"0b001704",
			4713 => x"ff864a29",
			4714 => x"07002a04",
			4715 => x"fffa4a29",
			4716 => x"00254a29",
			4717 => x"0001290c",
			4718 => x"05002704",
			4719 => x"ff7e4a29",
			4720 => x"07002f04",
			4721 => x"006b4a29",
			4722 => x"ffc34a29",
			4723 => x"0f00d204",
			4724 => x"ff314a29",
			4725 => x"0600c104",
			4726 => x"00144a29",
			4727 => x"ffd34a29",
			4728 => x"05002f04",
			4729 => x"ffcc4a29",
			4730 => x"04002704",
			4731 => x"007f4a29",
			4732 => x"ffe84a29",
			4733 => x"01000f10",
			4734 => x"0001240c",
			4735 => x"07002b08",
			4736 => x"07002a04",
			4737 => x"fffb4a29",
			4738 => x"00104a29",
			4739 => x"ffc84a29",
			4740 => x"00a44a29",
			4741 => x"03002408",
			4742 => x"09002204",
			4743 => x"003a4a29",
			4744 => x"ffe84a29",
			4745 => x"ff9b4a29",
			4746 => x"04002e30",
			4747 => x"0000a804",
			4748 => x"fe804a8d",
			4749 => x"01001128",
			4750 => x"0b00191c",
			4751 => x"0600890c",
			4752 => x"07002a08",
			4753 => x"04001d04",
			4754 => x"00b84a8d",
			4755 => x"02084a8d",
			4756 => x"fe9b4a8d",
			4757 => x"03002108",
			4758 => x"00012004",
			4759 => x"01864a8d",
			4760 => x"007b4a8d",
			4761 => x"09001904",
			4762 => x"fe574a8d",
			4763 => x"001b4a8d",
			4764 => x"0a003608",
			4765 => x"0f00bf04",
			4766 => x"ff484a8d",
			4767 => x"02054a8d",
			4768 => x"ff9f4a8d",
			4769 => x"fe854a8d",
			4770 => x"fe724a8d",
			4771 => x"0400215c",
			4772 => x"04001d38",
			4773 => x"0d001728",
			4774 => x"0c001514",
			4775 => x"01000c10",
			4776 => x"09001908",
			4777 => x"00011904",
			4778 => x"00924b69",
			4779 => x"fec24b69",
			4780 => x"08001c04",
			4781 => x"01c14b69",
			4782 => x"ff5a4b69",
			4783 => x"fe9c4b69",
			4784 => x"07003410",
			4785 => x"03002108",
			4786 => x"0e007504",
			4787 => x"ff184b69",
			4788 => x"014e4b69",
			4789 => x"01000c04",
			4790 => x"feab4b69",
			4791 => x"00a64b69",
			4792 => x"00fb4b69",
			4793 => x"0d001808",
			4794 => x"08001d04",
			4795 => x"ffcc4b69",
			4796 => x"01d94b69",
			4797 => x"0c001b04",
			4798 => x"00044b69",
			4799 => x"ff404b69",
			4800 => x"0201311c",
			4801 => x"0b001710",
			4802 => x"09001d0c",
			4803 => x"0a002804",
			4804 => x"01ae4b69",
			4805 => x"08001804",
			4806 => x"feb14b69",
			4807 => x"00cb4b69",
			4808 => x"fe824b69",
			4809 => x"07003208",
			4810 => x"09002004",
			4811 => x"01a44b69",
			4812 => x"ffc64b69",
			4813 => x"ffcf4b69",
			4814 => x"0b001b04",
			4815 => x"fe914b69",
			4816 => x"002f4b69",
			4817 => x"09001e04",
			4818 => x"fe684b69",
			4819 => x"08001d08",
			4820 => x"0e007604",
			4821 => x"fed64b69",
			4822 => x"01734b69",
			4823 => x"00015304",
			4824 => x"fe764b69",
			4825 => x"01214b69",
			4826 => x"01000e60",
			4827 => x"0d001438",
			4828 => x"0100091c",
			4829 => x"0a00230c",
			4830 => x"0e007508",
			4831 => x"04001804",
			4832 => x"ffde4c55",
			4833 => x"00054c55",
			4834 => x"002a4c55",
			4835 => x"0b00170c",
			4836 => x"0200db08",
			4837 => x"0000d204",
			4838 => x"fff44c55",
			4839 => x"001b4c55",
			4840 => x"ff744c55",
			4841 => x"000d4c55",
			4842 => x"0e008f18",
			4843 => x"0500290c",
			4844 => x"0b001608",
			4845 => x"09001904",
			4846 => x"ffed4c55",
			4847 => x"008f4c55",
			4848 => x"ffe14c55",
			4849 => x"00012708",
			4850 => x"0b001604",
			4851 => x"000f4c55",
			4852 => x"fffc4c55",
			4853 => x"ffd24c55",
			4854 => x"ffc94c55",
			4855 => x"01000a10",
			4856 => x"06009c0c",
			4857 => x"0000f208",
			4858 => x"0000dd04",
			4859 => x"fff24c55",
			4860 => x"001e4c55",
			4861 => x"ffc54c55",
			4862 => x"00a24c55",
			4863 => x"04002008",
			4864 => x"08001c04",
			4865 => x"00244c55",
			4866 => x"ff924c55",
			4867 => x"01000b04",
			4868 => x"ffcf4c55",
			4869 => x"0e008108",
			4870 => x"07002f04",
			4871 => x"00664c55",
			4872 => x"ffee4c55",
			4873 => x"fff64c55",
			4874 => x"02014814",
			4875 => x"04001808",
			4876 => x"04001604",
			4877 => x"fff84c55",
			4878 => x"001b4c55",
			4879 => x"03002408",
			4880 => x"03002304",
			4881 => x"fff24c55",
			4882 => x"00104c55",
			4883 => x"ff7a4c55",
			4884 => x"00224c55",
			4885 => x"0f009214",
			4886 => x"09001e10",
			4887 => x"0c001a0c",
			4888 => x"0d001208",
			4889 => x"01000b04",
			4890 => x"fe9d4d19",
			4891 => x"019b4d19",
			4892 => x"fe784d19",
			4893 => x"01b54d19",
			4894 => x"fe714d19",
			4895 => x"03002728",
			4896 => x"0b001924",
			4897 => x"0c001510",
			4898 => x"0c001204",
			4899 => x"ff314d19",
			4900 => x"0a002c08",
			4901 => x"04001804",
			4902 => x"015f4d19",
			4903 => x"02fd4d19",
			4904 => x"fe9b4d19",
			4905 => x"00011108",
			4906 => x"04001704",
			4907 => x"000d4d19",
			4908 => x"fe114d19",
			4909 => x"08001804",
			4910 => x"ff464d19",
			4911 => x"0f00c304",
			4912 => x"01824d19",
			4913 => x"00414d19",
			4914 => x"02804d19",
			4915 => x"05002b04",
			4916 => x"fe4a4d19",
			4917 => x"08001f18",
			4918 => x"0400210c",
			4919 => x"08001804",
			4920 => x"fe954d19",
			4921 => x"0f00c504",
			4922 => x"02114d19",
			4923 => x"013f4d19",
			4924 => x"09001e04",
			4925 => x"fe524d19",
			4926 => x"07003304",
			4927 => x"01844d19",
			4928 => x"ff2b4d19",
			4929 => x"0c001d04",
			4930 => x"fe4d4d19",
			4931 => x"08002404",
			4932 => x"01f74d19",
			4933 => x"fe904d19",
			4934 => x"04001e48",
			4935 => x"0d00173c",
			4936 => x"0d001324",
			4937 => x"05002414",
			4938 => x"0300210c",
			4939 => x"07002504",
			4940 => x"ff1b4dfd",
			4941 => x"0000fc04",
			4942 => x"ffa94dfd",
			4943 => x"01304dfd",
			4944 => x"05002004",
			4945 => x"fffa4dfd",
			4946 => x"fec64dfd",
			4947 => x"0300270c",
			4948 => x"04001804",
			4949 => x"ffee4dfd",
			4950 => x"0c001504",
			4951 => x"01594dfd",
			4952 => x"00b84dfd",
			4953 => x"ff354dfd",
			4954 => x"07002b0c",
			4955 => x"01000c08",
			4956 => x"0c001604",
			4957 => x"01004dfd",
			4958 => x"ff6e4dfd",
			4959 => x"fef34dfd",
			4960 => x"0a003108",
			4961 => x"0a002804",
			4962 => x"fffc4dfd",
			4963 => x"fe814dfd",
			4964 => x"005a4dfd",
			4965 => x"05002c08",
			4966 => x"0000e704",
			4967 => x"ffb04dfd",
			4968 => x"01814dfd",
			4969 => x"ff264dfd",
			4970 => x"05002a04",
			4971 => x"fe854dfd",
			4972 => x"05002f10",
			4973 => x"0400210c",
			4974 => x"0f00c308",
			4975 => x"04002004",
			4976 => x"ff8a4dfd",
			4977 => x"01874dfd",
			4978 => x"ff9d4dfd",
			4979 => x"ff024dfd",
			4980 => x"03002a04",
			4981 => x"feaf4dfd",
			4982 => x"09001d04",
			4983 => x"fecf4dfd",
			4984 => x"0d001508",
			4985 => x"05003a04",
			4986 => x"014e4dfd",
			4987 => x"ff474dfd",
			4988 => x"0c001d04",
			4989 => x"ff874dfd",
			4990 => x"00c14dfd",
			4991 => x"0f00b538",
			4992 => x"07002d34",
			4993 => x"07002c28",
			4994 => x"0300291c",
			4995 => x"05002710",
			4996 => x"07002808",
			4997 => x"0c001504",
			4998 => x"00c44ed1",
			4999 => x"fede4ed1",
			5000 => x"03001d04",
			5001 => x"003c4ed1",
			5002 => x"fe974ed1",
			5003 => x"09001d08",
			5004 => x"0000be04",
			5005 => x"ff954ed1",
			5006 => x"01384ed1",
			5007 => x"fef94ed1",
			5008 => x"01000c04",
			5009 => x"fe894ed1",
			5010 => x"0000a804",
			5011 => x"ffc94ed1",
			5012 => x"00f64ed1",
			5013 => x"01000b04",
			5014 => x"ffad4ed1",
			5015 => x"08002204",
			5016 => x"017f4ed1",
			5017 => x"fff04ed1",
			5018 => x"fe6a4ed1",
			5019 => x"0d001928",
			5020 => x"0d001720",
			5021 => x"0500351c",
			5022 => x"0800190c",
			5023 => x"02013108",
			5024 => x"05002c04",
			5025 => x"01284ed1",
			5026 => x"fed24ed1",
			5027 => x"fec54ed1",
			5028 => x"04001708",
			5029 => x"05002204",
			5030 => x"ffac4ed1",
			5031 => x"fe754ed1",
			5032 => x"00012904",
			5033 => x"00a24ed1",
			5034 => x"ff864ed1",
			5035 => x"013b4ed1",
			5036 => x"05002f04",
			5037 => x"019f4ed1",
			5038 => x"000c4ed1",
			5039 => x"0f00db04",
			5040 => x"febd4ed1",
			5041 => x"0600c704",
			5042 => x"00244ed1",
			5043 => x"ffc74ed1",
			5044 => x"0d001430",
			5045 => x"0a002710",
			5046 => x"07002304",
			5047 => x"ffb94fbd",
			5048 => x"0000be04",
			5049 => x"ffe24fbd",
			5050 => x"0a002304",
			5051 => x"00a24fbd",
			5052 => x"002d4fbd",
			5053 => x"01000d1c",
			5054 => x"09001c14",
			5055 => x"0b001410",
			5056 => x"0600af08",
			5057 => x"0e006e04",
			5058 => x"001b4fbd",
			5059 => x"ff8b4fbd",
			5060 => x"00013904",
			5061 => x"005a4fbd",
			5062 => x"ffc64fbd",
			5063 => x"ff134fbd",
			5064 => x"03002704",
			5065 => x"00654fbd",
			5066 => x"ffb64fbd",
			5067 => x"003e4fbd",
			5068 => x"09001b08",
			5069 => x"0a002c04",
			5070 => x"00ba4fbd",
			5071 => x"ffd44fbd",
			5072 => x"0b001610",
			5073 => x"05002704",
			5074 => x"00254fbd",
			5075 => x"0d001508",
			5076 => x"0a002f04",
			5077 => x"ffd44fbd",
			5078 => x"002f4fbd",
			5079 => x"ff4f4fbd",
			5080 => x"0e008214",
			5081 => x"07002f0c",
			5082 => x"05003808",
			5083 => x"0f006904",
			5084 => x"ffe94fbd",
			5085 => x"00cd4fbd",
			5086 => x"ffd34fbd",
			5087 => x"03002404",
			5088 => x"000e4fbd",
			5089 => x"ffc34fbd",
			5090 => x"05003510",
			5091 => x"0b001908",
			5092 => x"0b001704",
			5093 => x"00164fbd",
			5094 => x"ff354fbd",
			5095 => x"02013704",
			5096 => x"ffcb4fbd",
			5097 => x"00694fbd",
			5098 => x"02012d04",
			5099 => x"ffcc4fbd",
			5100 => x"02013604",
			5101 => x"00a94fbd",
			5102 => x"fff34fbd",
			5103 => x"07002304",
			5104 => x"fee35059",
			5105 => x"03002108",
			5106 => x"0000e904",
			5107 => x"ff5f5059",
			5108 => x"01505059",
			5109 => x"0b00161c",
			5110 => x"04002118",
			5111 => x"0f00a908",
			5112 => x"04001d04",
			5113 => x"ffe15059",
			5114 => x"00ea5059",
			5115 => x"0f00bf08",
			5116 => x"0f00b104",
			5117 => x"00045059",
			5118 => x"fe865059",
			5119 => x"00012f04",
			5120 => x"01215059",
			5121 => x"ffa35059",
			5122 => x"fea95059",
			5123 => x"01000a0c",
			5124 => x"05002a04",
			5125 => x"ff055059",
			5126 => x"00011b04",
			5127 => x"ff205059",
			5128 => x"01385059",
			5129 => x"07002f0c",
			5130 => x"0d001404",
			5131 => x"ff005059",
			5132 => x"01000b04",
			5133 => x"ff7b5059",
			5134 => x"01155059",
			5135 => x"0e009008",
			5136 => x"05002904",
			5137 => x"00985059",
			5138 => x"fe945059",
			5139 => x"0e009204",
			5140 => x"01195059",
			5141 => x"ff7b5059",
			5142 => x"07002304",
			5143 => x"ff015127",
			5144 => x"0a002820",
			5145 => x"04001e1c",
			5146 => x"04001d18",
			5147 => x"0c00160c",
			5148 => x"0f00b408",
			5149 => x"09001904",
			5150 => x"ff765127",
			5151 => x"006b5127",
			5152 => x"01545127",
			5153 => x"03002108",
			5154 => x"05001e04",
			5155 => x"ffc35127",
			5156 => x"00b75127",
			5157 => x"feb85127",
			5158 => x"01695127",
			5159 => x"ff0d5127",
			5160 => x"05002a14",
			5161 => x"0f00c004",
			5162 => x"fe9e5127",
			5163 => x"01000908",
			5164 => x"0b001304",
			5165 => x"00275127",
			5166 => x"fec05127",
			5167 => x"0600b704",
			5168 => x"00eb5127",
			5169 => x"ff1a5127",
			5170 => x"0a00341c",
			5171 => x"05003310",
			5172 => x"04002108",
			5173 => x"0f00c304",
			5174 => x"00f15127",
			5175 => x"ff905127",
			5176 => x"0b001904",
			5177 => x"feb85127",
			5178 => x"00bf5127",
			5179 => x"0d001808",
			5180 => x"0c001804",
			5181 => x"ffa65127",
			5182 => x"014e5127",
			5183 => x"ff7e5127",
			5184 => x"0c001d0c",
			5185 => x"07003208",
			5186 => x"07002e04",
			5187 => x"ff175127",
			5188 => x"00b05127",
			5189 => x"feb75127",
			5190 => x"09002504",
			5191 => x"01025127",
			5192 => x"ff9b5127",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1797, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3471, initial_addr_3'length));
	end generate gen_rom_4;

	gen_rom_5: if SELECT_ROM = 5 generate
		bank <= (
			0 => x"06009510",
			1 => x"0f008004",
			2 => x"fe630085",
			3 => x"0000d708",
			4 => x"05002704",
			5 => x"fe690085",
			6 => x"02e60085",
			7 => x"fe5f0085",
			8 => x"01000c10",
			9 => x"0e009308",
			10 => x"07002904",
			11 => x"00680085",
			12 => x"fe550085",
			13 => x"00013a04",
			14 => x"fe910085",
			15 => x"00be0085",
			16 => x"05003918",
			17 => x"07004414",
			18 => x"0001460c",
			19 => x"0f00b104",
			20 => x"02db0085",
			21 => x"08001f04",
			22 => x"fefc0085",
			23 => x"013c0085",
			24 => x"08002404",
			25 => x"01c30085",
			26 => x"02b20085",
			27 => x"fe700085",
			28 => x"0a004308",
			29 => x"07003704",
			30 => x"00a70085",
			31 => x"fe590085",
			32 => x"02950085",
			33 => x"00011f18",
			34 => x"0f008004",
			35 => x"fe600101",
			36 => x"07002f08",
			37 => x"08001d04",
			38 => x"fe560101",
			39 => x"04c40101",
			40 => x"01001604",
			41 => x"fe510101",
			42 => x"00011404",
			43 => x"00300101",
			44 => x"fe720101",
			45 => x"08001c04",
			46 => x"fe600101",
			47 => x"0d00211c",
			48 => x"0a004218",
			49 => x"05003910",
			50 => x"0600a608",
			51 => x"0600a204",
			52 => x"01a00101",
			53 => x"fe380101",
			54 => x"0f00c404",
			55 => x"045a0101",
			56 => x"02360101",
			57 => x"07003904",
			58 => x"012d0101",
			59 => x"fe500101",
			60 => x"04af0101",
			61 => x"01001804",
			62 => x"00bb0101",
			63 => x"fe500101",
			64 => x"0f00a90c",
			65 => x"0f008004",
			66 => x"fe5e0175",
			67 => x"0e006804",
			68 => x"007d0175",
			69 => x"fe600175",
			70 => x"01000a04",
			71 => x"fe5c0175",
			72 => x"07004024",
			73 => x"02012e14",
			74 => x"01000e08",
			75 => x"0000fa04",
			76 => x"00d50175",
			77 => x"fe570175",
			78 => x"07003104",
			79 => x"03f10175",
			80 => x"03003804",
			81 => x"005c0175",
			82 => x"03ce0175",
			83 => x"0f00c904",
			84 => x"03a90175",
			85 => x"0e008f04",
			86 => x"008e0175",
			87 => x"07003c04",
			88 => x"02cc0175",
			89 => x"01310175",
			90 => x"05003504",
			91 => x"00010175",
			92 => x"fe610175",
			93 => x"02012634",
			94 => x"0c001a20",
			95 => x"04002210",
			96 => x"0700300c",
			97 => x"01000c04",
			98 => x"ff820241",
			99 => x"0000c704",
			100 => x"ffa70241",
			101 => x"00a60241",
			102 => x"ff3a0241",
			103 => x"06007404",
			104 => x"ff9e0241",
			105 => x"03003308",
			106 => x"08001c04",
			107 => x"fff30241",
			108 => x"00df0241",
			109 => x"ffda0241",
			110 => x"01001a0c",
			111 => x"03004404",
			112 => x"feda0241",
			113 => x"0b001b04",
			114 => x"00380241",
			115 => x"ffe70241",
			116 => x"0e009104",
			117 => x"ffe00241",
			118 => x"00950241",
			119 => x"01001928",
			120 => x"01001010",
			121 => x"0b00170c",
			122 => x"01000a04",
			123 => x"ff7e0241",
			124 => x"08001c04",
			125 => x"ff9f0241",
			126 => x"00a40241",
			127 => x"ff3d0241",
			128 => x"07004010",
			129 => x"03002c04",
			130 => x"00d30241",
			131 => x"05003604",
			132 => x"ffa30241",
			133 => x"05003904",
			134 => x"00f80241",
			135 => x"002d0241",
			136 => x"04002b04",
			137 => x"ff780241",
			138 => x"00370241",
			139 => x"01001a04",
			140 => x"ff3a0241",
			141 => x"0f00d904",
			142 => x"ffc70241",
			143 => x"00430241",
			144 => x"0f00ae14",
			145 => x"0f008004",
			146 => x"fe5902e5",
			147 => x"0e006804",
			148 => x"028c02e5",
			149 => x"0200cb08",
			150 => x"0000c304",
			151 => x"fe6a02e5",
			152 => x"014402e5",
			153 => x"fe5402e5",
			154 => x"0d001f34",
			155 => x"01000c10",
			156 => x"00014508",
			157 => x"07003404",
			158 => x"fe5802e5",
			159 => x"005602e5",
			160 => x"0b001404",
			161 => x"031102e5",
			162 => x"ff3e02e5",
			163 => x"00014618",
			164 => x"0e009110",
			165 => x"01001008",
			166 => x"0e008a04",
			167 => x"ff9102e5",
			168 => x"047502e5",
			169 => x"0b001b04",
			170 => x"067f02e5",
			171 => x"00fc02e5",
			172 => x"00013b04",
			173 => x"fe6202e5",
			174 => x"022a02e5",
			175 => x"05003908",
			176 => x"0f00db04",
			177 => x"05e002e5",
			178 => x"047602e5",
			179 => x"012802e5",
			180 => x"01001708",
			181 => x"0d002004",
			182 => x"fe5902e5",
			183 => x"031f02e5",
			184 => x"fe4f02e5",
			185 => x"0f008c0c",
			186 => x"0b001308",
			187 => x"04001d04",
			188 => x"fe930369",
			189 => x"03cc0369",
			190 => x"fe610369",
			191 => x"01000a04",
			192 => x"fe650369",
			193 => x"0b001718",
			194 => x"05002408",
			195 => x"0a002a04",
			196 => x"ffb50369",
			197 => x"fe450369",
			198 => x"06009a04",
			199 => x"02ac0369",
			200 => x"02010f04",
			201 => x"fe7c0369",
			202 => x"08001c04",
			203 => x"fe870369",
			204 => x"01af0369",
			205 => x"0d00180c",
			206 => x"0a003d08",
			207 => x"04002504",
			208 => x"fdff0369",
			209 => x"fec30369",
			210 => x"010d0369",
			211 => x"0f00af04",
			212 => x"fe5b0369",
			213 => x"0d002208",
			214 => x"01001a04",
			215 => x"00ca0369",
			216 => x"02f00369",
			217 => x"fe610369",
			218 => x"02012e34",
			219 => x"0f00a914",
			220 => x"0f008004",
			221 => x"fe57041d",
			222 => x"0e006804",
			223 => x"0390041d",
			224 => x"0a002a08",
			225 => x"0000c604",
			226 => x"fe67041d",
			227 => x"010b041d",
			228 => x"fe5a041d",
			229 => x"01000c04",
			230 => x"fe5b041d",
			231 => x"08002610",
			232 => x"0600a104",
			233 => x"0a2a041d",
			234 => x"00012404",
			235 => x"fe60041d",
			236 => x"02012004",
			237 => x"0875041d",
			238 => x"01cb041d",
			239 => x"05003504",
			240 => x"0247041d",
			241 => x"05004904",
			242 => x"fe56041d",
			243 => x"0049041d",
			244 => x"07004020",
			245 => x"01000c08",
			246 => x"01000a04",
			247 => x"fe56041d",
			248 => x"0210041d",
			249 => x"07003c10",
			250 => x"08001f04",
			251 => x"04c4041d",
			252 => x"03002f08",
			253 => x"03002c04",
			254 => x"07ff041d",
			255 => x"064e041d",
			256 => x"0a2e041d",
			257 => x"05003804",
			258 => x"0574041d",
			259 => x"ff54041d",
			260 => x"03002e04",
			261 => x"018f041d",
			262 => x"fe5d041d",
			263 => x"0d002130",
			264 => x"08001b04",
			265 => x"fe8d0481",
			266 => x"0d00201c",
			267 => x"0d001e18",
			268 => x"07003e10",
			269 => x"0d001a08",
			270 => x"0b001804",
			271 => x"006a0481",
			272 => x"ff420481",
			273 => x"02013304",
			274 => x"00570481",
			275 => x"01c00481",
			276 => x"01001404",
			277 => x"00120481",
			278 => x"fe890481",
			279 => x"fe700481",
			280 => x"03003108",
			281 => x"05001f04",
			282 => x"ffe10481",
			283 => x"01e90481",
			284 => x"0a004a04",
			285 => x"fea70481",
			286 => x"01580481",
			287 => x"fe840481",
			288 => x"02012638",
			289 => x"0c001a24",
			290 => x"04002210",
			291 => x"0700300c",
			292 => x"01000c04",
			293 => x"ff87055d",
			294 => x"0000c704",
			295 => x"ffab055d",
			296 => x"009c055d",
			297 => x"ff44055d",
			298 => x"09001f0c",
			299 => x"0000c008",
			300 => x"0000ab04",
			301 => x"fff6055d",
			302 => x"0058055d",
			303 => x"ff77055d",
			304 => x"06007c04",
			305 => x"ffd8055d",
			306 => x"00cc055d",
			307 => x"01001a0c",
			308 => x"03004404",
			309 => x"fee6055d",
			310 => x"0b001b04",
			311 => x"0037055d",
			312 => x"ffe8055d",
			313 => x"0e009104",
			314 => x"ffe0055d",
			315 => x"008f055d",
			316 => x"0100192c",
			317 => x"08002014",
			318 => x"03002708",
			319 => x"08001b04",
			320 => x"ffcc055d",
			321 => x"0089055d",
			322 => x"05003608",
			323 => x"0e009b04",
			324 => x"ff0f055d",
			325 => x"000c055d",
			326 => x"003b055d",
			327 => x"04002104",
			328 => x"00d8055d",
			329 => x"08002a10",
			330 => x"0b001b08",
			331 => x"08002304",
			332 => x"00a2055d",
			333 => x"ffe6055d",
			334 => x"02013004",
			335 => x"ff2d055d",
			336 => x"000a055d",
			337 => x"00a7055d",
			338 => x"01001a04",
			339 => x"ff44055d",
			340 => x"0f00d904",
			341 => x"ffc8055d",
			342 => x"0041055d",
			343 => x"0f008c0c",
			344 => x"0c001608",
			345 => x"01001004",
			346 => x"fe7005d1",
			347 => x"024d05d1",
			348 => x"fe6505d1",
			349 => x"01000a04",
			350 => x"fe6b05d1",
			351 => x"07002a04",
			352 => x"022105d1",
			353 => x"0e008e14",
			354 => x"09002610",
			355 => x"01001008",
			356 => x"06009604",
			357 => x"019d05d1",
			358 => x"feb005d1",
			359 => x"04001e04",
			360 => x"ff9405d1",
			361 => x"012f05d1",
			362 => x"fe5405d1",
			363 => x"0e00a30c",
			364 => x"00012204",
			365 => x"fe7805d1",
			366 => x"00012804",
			367 => x"035605d1",
			368 => x"010505d1",
			369 => x"03002e04",
			370 => x"00c805d1",
			371 => x"fe5005d1",
			372 => x"0d002134",
			373 => x"0e00a42c",
			374 => x"0f00d620",
			375 => x"04001804",
			376 => x"fed1063d",
			377 => x"01001210",
			378 => x"05003408",
			379 => x"08002204",
			380 => x"ffeb063d",
			381 => x"00fa063d",
			382 => x"02013404",
			383 => x"fed2063d",
			384 => x"002a063d",
			385 => x"04001b04",
			386 => x"fec5063d",
			387 => x"0d001b04",
			388 => x"00d9063d",
			389 => x"0021063d",
			390 => x"0c001404",
			391 => x"ff77063d",
			392 => x"0e009a04",
			393 => x"0134063d",
			394 => x"0095063d",
			395 => x"0f00e504",
			396 => x"febc063d",
			397 => x"003c063d",
			398 => x"feab063d",
			399 => x"0f008c0c",
			400 => x"0c001608",
			401 => x"01001004",
			402 => x"fe6c06c1",
			403 => x"020306c1",
			404 => x"fe6106c1",
			405 => x"01000a04",
			406 => x"fe6206c1",
			407 => x"0b00161c",
			408 => x"05002408",
			409 => x"0c001404",
			410 => x"fe2606c1",
			411 => x"003906c1",
			412 => x"08001c08",
			413 => x"0f00bf04",
			414 => x"017506c1",
			415 => x"fe7f06c1",
			416 => x"0f00c904",
			417 => x"02d306c1",
			418 => x"00014704",
			419 => x"ff7206c1",
			420 => x"021f06c1",
			421 => x"01000e04",
			422 => x"fe0f06c1",
			423 => x"03004110",
			424 => x"05003508",
			425 => x"0600b704",
			426 => x"007b06c1",
			427 => x"022006c1",
			428 => x"07003f04",
			429 => x"002906c1",
			430 => x"fe5e06c1",
			431 => x"02f906c1",
			432 => x"06007404",
			433 => x"fe74071d",
			434 => x"09002b28",
			435 => x"01001a20",
			436 => x"0b00201c",
			437 => x"08002610",
			438 => x"04002308",
			439 => x"01000c04",
			440 => x"fecf071d",
			441 => x"002b071d",
			442 => x"07003404",
			443 => x"014f071d",
			444 => x"0027071d",
			445 => x"03002a04",
			446 => x"0083071d",
			447 => x"0a003704",
			448 => x"fe52071d",
			449 => x"ff8d071d",
			450 => x"0201071d",
			451 => x"03003304",
			452 => x"0285071d",
			453 => x"ff16071d",
			454 => x"fe77071d",
			455 => x"0f008004",
			456 => x"fe700771",
			457 => x"08001b04",
			458 => x"fe7b0771",
			459 => x"07002a04",
			460 => x"01dd0771",
			461 => x"0a002804",
			462 => x"fec30771",
			463 => x"0300290c",
			464 => x"01001608",
			465 => x"0c001804",
			466 => x"011d0771",
			467 => x"ff140771",
			468 => x"028f0771",
			469 => x"05003308",
			470 => x"0b001a04",
			471 => x"00550771",
			472 => x"fe7e0771",
			473 => x"01001204",
			474 => x"ffce0771",
			475 => x"00e40771",
			476 => x"05002718",
			477 => x"07002908",
			478 => x"03002404",
			479 => x"fff20835",
			480 => x"00170835",
			481 => x"03002108",
			482 => x"03001f04",
			483 => x"fff40835",
			484 => x"00160835",
			485 => x"0e00a104",
			486 => x"ff7b0835",
			487 => x"00040835",
			488 => x"02011a24",
			489 => x"0f00b31c",
			490 => x"05003518",
			491 => x"0a002d0c",
			492 => x"05002904",
			493 => x"001d0835",
			494 => x"05002d04",
			495 => x"ffc90835",
			496 => x"00090835",
			497 => x"0b001a08",
			498 => x"08001c04",
			499 => x"fff90835",
			500 => x"007b0835",
			501 => x"fff30835",
			502 => x"ffc20835",
			503 => x"07003104",
			504 => x"fffc0835",
			505 => x"ff760835",
			506 => x"0c001808",
			507 => x"01000a04",
			508 => x"ffd60835",
			509 => x"00880835",
			510 => x"09002108",
			511 => x"09001e04",
			512 => x"fffc0835",
			513 => x"ff870835",
			514 => x"05003308",
			515 => x"00014604",
			516 => x"ff9d0835",
			517 => x"00340835",
			518 => x"05003808",
			519 => x"09002b04",
			520 => x"00980835",
			521 => x"ffcf0835",
			522 => x"0a004304",
			523 => x"ffb80835",
			524 => x"00540835",
			525 => x"0201264c",
			526 => x"0c001c38",
			527 => x"0600951c",
			528 => x"01000b10",
			529 => x"0b00150c",
			530 => x"03002404",
			531 => x"fff50939",
			532 => x"0000d704",
			533 => x"00430939",
			534 => x"fffa0939",
			535 => x"ffd90939",
			536 => x"03002108",
			537 => x"03001d04",
			538 => x"fff00939",
			539 => x"00280939",
			540 => x"ff520939",
			541 => x"06009d0c",
			542 => x"0f00b308",
			543 => x"01000a04",
			544 => x"fffb0939",
			545 => x"00b60939",
			546 => x"ffe10939",
			547 => x"00012704",
			548 => x"ff620939",
			549 => x"0600a204",
			550 => x"ffbf0939",
			551 => x"0f00c804",
			552 => x"00880939",
			553 => x"ffed0939",
			554 => x"01001a0c",
			555 => x"0a005404",
			556 => x"ff470939",
			557 => x"05007604",
			558 => x"000c0939",
			559 => x"fffb0939",
			560 => x"0e009104",
			561 => x"fff00939",
			562 => x"00460939",
			563 => x"0600ad14",
			564 => x"0600a708",
			565 => x"00013c04",
			566 => x"ff9a0939",
			567 => x"003b0939",
			568 => x"0f00c908",
			569 => x"01000e04",
			570 => x"00130939",
			571 => x"00f00939",
			572 => x"ffef0939",
			573 => x"00014810",
			574 => x"0d001c08",
			575 => x"03002f04",
			576 => x"ff2d0939",
			577 => x"00280939",
			578 => x"05003804",
			579 => x"00520939",
			580 => x"ff950939",
			581 => x"0100180c",
			582 => x"02014408",
			583 => x"08002204",
			584 => x"ffcc0939",
			585 => x"00530939",
			586 => x"00af0939",
			587 => x"01001a04",
			588 => x"ff9c0939",
			589 => x"001e0939",
			590 => x"09002540",
			591 => x"0c001b2c",
			592 => x"0d001a28",
			593 => x"0b00181c",
			594 => x"01000e0c",
			595 => x"0b001508",
			596 => x"08001c04",
			597 => x"fe940a15",
			598 => x"00a00a15",
			599 => x"fe6f0a15",
			600 => x"0e008808",
			601 => x"0000c704",
			602 => x"fed20a15",
			603 => x"01510a15",
			604 => x"03002d04",
			605 => x"fed60a15",
			606 => x"00c40a15",
			607 => x"0a003704",
			608 => x"fe6f0a15",
			609 => x"09002104",
			610 => x"ff3e0a15",
			611 => x"00d30a15",
			612 => x"01390a15",
			613 => x"0a003b08",
			614 => x"02013504",
			615 => x"fe260a15",
			616 => x"00030a15",
			617 => x"0c001c08",
			618 => x"09002204",
			619 => x"ff550a15",
			620 => x"01b80a15",
			621 => x"ff390a15",
			622 => x"05003820",
			623 => x"0300270c",
			624 => x"0d001b08",
			625 => x"0d001a04",
			626 => x"ffec0a15",
			627 => x"00230a15",
			628 => x"fe900a15",
			629 => x"09002b10",
			630 => x"0e008604",
			631 => x"fecf0a15",
			632 => x"05003304",
			633 => x"00c60a15",
			634 => x"01001704",
			635 => x"02110a15",
			636 => x"008f0a15",
			637 => x"fec00a15",
			638 => x"03004608",
			639 => x"08002404",
			640 => x"007c0a15",
			641 => x"fe790a15",
			642 => x"04004a04",
			643 => x"017d0a15",
			644 => x"ff350a15",
			645 => x"0b001838",
			646 => x"02011b20",
			647 => x"0e00841c",
			648 => x"0e007910",
			649 => x"0f008108",
			650 => x"06007104",
			651 => x"ffd90b01",
			652 => x"00310b01",
			653 => x"04002604",
			654 => x"ffaf0b01",
			655 => x"00070b01",
			656 => x"02011508",
			657 => x"01000b04",
			658 => x"fff90b01",
			659 => x"00740b01",
			660 => x"ffec0b01",
			661 => x"ff960b01",
			662 => x"01000a04",
			663 => x"ffc90b01",
			664 => x"0e008e0c",
			665 => x"0600a404",
			666 => x"00230b01",
			667 => x"0f00c704",
			668 => x"ffca0b01",
			669 => x"00110b01",
			670 => x"0c001404",
			671 => x"00010b01",
			672 => x"00ab0b01",
			673 => x"0d001a10",
			674 => x"00012e0c",
			675 => x"03002d04",
			676 => x"ffd00b01",
			677 => x"00010604",
			678 => x"fff00b01",
			679 => x"00470b01",
			680 => x"ff690b01",
			681 => x"02012614",
			682 => x"0200fd08",
			683 => x"0000ff04",
			684 => x"ffed0b01",
			685 => x"003f0b01",
			686 => x"03003804",
			687 => x"ff6f0b01",
			688 => x"03003b04",
			689 => x"00230b01",
			690 => x"fff20b01",
			691 => x"0d001f0c",
			692 => x"04002708",
			693 => x"05003304",
			694 => x"00100b01",
			695 => x"008a0b01",
			696 => x"ffed0b01",
			697 => x"04002b04",
			698 => x"ff880b01",
			699 => x"08002a04",
			700 => x"ffe90b01",
			701 => x"07004404",
			702 => x"005e0b01",
			703 => x"fff20b01",
			704 => x"0d002134",
			705 => x"0e00a52c",
			706 => x"02013f24",
			707 => x"01001a20",
			708 => x"0600aa10",
			709 => x"01001208",
			710 => x"07003304",
			711 => x"00350b6d",
			712 => x"fea70b6d",
			713 => x"01001704",
			714 => x"00a20b6d",
			715 => x"ff240b6d",
			716 => x"0e008e08",
			717 => x"0e008804",
			718 => x"007b0b6d",
			719 => x"fea10b6d",
			720 => x"07003f04",
			721 => x"001b0b6d",
			722 => x"fed90b6d",
			723 => x"00f40b6d",
			724 => x"04001d04",
			725 => x"00000b6d",
			726 => x"01370b6d",
			727 => x"03002e04",
			728 => x"ffd20b6d",
			729 => x"fedb0b6d",
			730 => x"feb80b6d",
			731 => x"0a004350",
			732 => x"05003934",
			733 => x"0b001f28",
			734 => x"08002010",
			735 => x"0c00190c",
			736 => x"09001f08",
			737 => x"0b001304",
			738 => x"00500c19",
			739 => x"ff830c19",
			740 => x"00b00c19",
			741 => x"ff280c19",
			742 => x"00014610",
			743 => x"0f00c608",
			744 => x"0600a804",
			745 => x"001d0c19",
			746 => x"00c00c19",
			747 => x"03002d04",
			748 => x"003a0c19",
			749 => x"ff5f0c19",
			750 => x"0d001c04",
			751 => x"01030c19",
			752 => x"00510c19",
			753 => x"01001708",
			754 => x"09002a04",
			755 => x"ff8d0c19",
			756 => x"00bb0c19",
			757 => x"ff060c19",
			758 => x"08002414",
			759 => x"0c001b0c",
			760 => x"0f00b908",
			761 => x"0000f204",
			762 => x"ffe10c19",
			763 => x"00460c19",
			764 => x"ff470c19",
			765 => x"0a003d04",
			766 => x"00990c19",
			767 => x"ffd60c19",
			768 => x"02013a04",
			769 => x"feea0c19",
			770 => x"fff40c19",
			771 => x"00012804",
			772 => x"ffd80c19",
			773 => x"00ce0c19",
			774 => x"0700404c",
			775 => x"0f00a918",
			776 => x"01000b0c",
			777 => x"0b001508",
			778 => x"03002404",
			779 => x"fff70cb5",
			780 => x"00330cb5",
			781 => x"ffe00cb5",
			782 => x"03002108",
			783 => x"03001d04",
			784 => x"fff10cb5",
			785 => x"00200cb5",
			786 => x"ff6f0cb5",
			787 => x"0f00cd20",
			788 => x"00013c14",
			789 => x"00013710",
			790 => x"0c001c08",
			791 => x"01000c04",
			792 => x"ffc70cb5",
			793 => x"00620cb5",
			794 => x"0e009104",
			795 => x"ffa70cb5",
			796 => x"004c0cb5",
			797 => x"ff9e0cb5",
			798 => x"01001008",
			799 => x"0e008704",
			800 => x"002e0cb5",
			801 => x"ffc30cb5",
			802 => x"00a70cb5",
			803 => x"00015710",
			804 => x"0500330c",
			805 => x"00014604",
			806 => x"ff5f0cb5",
			807 => x"0600b704",
			808 => x"ffdb0cb5",
			809 => x"00310cb5",
			810 => x"fff30cb5",
			811 => x"00610cb5",
			812 => x"ff730cb5",
			813 => x"07004058",
			814 => x"00011f28",
			815 => x"0f00b31c",
			816 => x"0f00ae18",
			817 => x"06007f0c",
			818 => x"0f008004",
			819 => x"ff590d81",
			820 => x"0d001504",
			821 => x"ff980d81",
			822 => x"00a10d81",
			823 => x"03002408",
			824 => x"09001a04",
			825 => x"ffcf0d81",
			826 => x"00280d81",
			827 => x"ff020d81",
			828 => x"00c30d81",
			829 => x"04001a08",
			830 => x"07003204",
			831 => x"00250d81",
			832 => x"ffef0d81",
			833 => x"fee90d81",
			834 => x"0d001d20",
			835 => x"07003714",
			836 => x"01001210",
			837 => x"0600a908",
			838 => x"00013e04",
			839 => x"ff000d81",
			840 => x"00700d81",
			841 => x"0f00cd04",
			842 => x"00a80d81",
			843 => x"ffda0d81",
			844 => x"00da0d81",
			845 => x"0600b708",
			846 => x"01001604",
			847 => x"ff9c0d81",
			848 => x"fee60d81",
			849 => x"00600d81",
			850 => x"03003308",
			851 => x"09002804",
			852 => x"01060d81",
			853 => x"00610d81",
			854 => x"04003104",
			855 => x"ff4d0d81",
			856 => x"008f0d81",
			857 => x"0c002104",
			858 => x"ff020d81",
			859 => x"00014904",
			860 => x"ff830d81",
			861 => x"02014204",
			862 => x"008d0d81",
			863 => x"ffbb0d81",
			864 => x"0f008004",
			865 => x"fe7e0dfd",
			866 => x"0e00a534",
			867 => x"02013f28",
			868 => x"01001a20",
			869 => x"0f00cd10",
			870 => x"0c001c08",
			871 => x"08001f04",
			872 => x"ffd50dfd",
			873 => x"00c80dfd",
			874 => x"0d002004",
			875 => x"ff470dfd",
			876 => x"01700dfd",
			877 => x"0600b808",
			878 => x"02013704",
			879 => x"fe1e0dfd",
			880 => x"ffbb0dfd",
			881 => x"07003f04",
			882 => x"01340dfd",
			883 => x"fe8a0dfd",
			884 => x"08002a04",
			885 => x"02a70dfd",
			886 => x"feb30dfd",
			887 => x"04002208",
			888 => x"02014b04",
			889 => x"00710dfd",
			890 => x"00fb0dfd",
			891 => x"01bc0dfd",
			892 => x"03002e04",
			893 => x"ffe40dfd",
			894 => x"fe670dfd",
			895 => x"06007404",
			896 => x"fe710e61",
			897 => x"09002b2c",
			898 => x"01001a24",
			899 => x"0b002020",
			900 => x"0b001910",
			901 => x"01000e08",
			902 => x"0b001504",
			903 => x"00700e61",
			904 => x"fe560e61",
			905 => x"0f00ce04",
			906 => x"013d0e61",
			907 => x"00250e61",
			908 => x"02011a08",
			909 => x"0a003604",
			910 => x"fe220e61",
			911 => x"ffe40e61",
			912 => x"05003304",
			913 => x"ff430e61",
			914 => x"005f0e61",
			915 => x"02570e61",
			916 => x"03003304",
			917 => x"02e80e61",
			918 => x"ff060e61",
			919 => x"fe710e61",
			920 => x"08002764",
			921 => x"07003648",
			922 => x"0c001828",
			923 => x"0500240c",
			924 => x"03002108",
			925 => x"03001f04",
			926 => x"ffe00f45",
			927 => x"001a0f45",
			928 => x"ff730f45",
			929 => x"05002e10",
			930 => x"0f008c08",
			931 => x"03002104",
			932 => x"00390f45",
			933 => x"ffa40f45",
			934 => x"08001b04",
			935 => x"ffda0f45",
			936 => x"00b20f45",
			937 => x"04002004",
			938 => x"ff810f45",
			939 => x"0e008604",
			940 => x"ffda0f45",
			941 => x"006c0f45",
			942 => x"08002310",
			943 => x"05003808",
			944 => x"04002604",
			945 => x"ff010f45",
			946 => x"00060f45",
			947 => x"04002a04",
			948 => x"004b0f45",
			949 => x"ffd10f45",
			950 => x"0c001c08",
			951 => x"00011f04",
			952 => x"00080f45",
			953 => x"005e0f45",
			954 => x"05003e04",
			955 => x"ff910f45",
			956 => x"000e0f45",
			957 => x"0a00360c",
			958 => x"0e008f04",
			959 => x"fff00f45",
			960 => x"08002004",
			961 => x"00140f45",
			962 => x"00d40f45",
			963 => x"03003508",
			964 => x"08002404",
			965 => x"00140f45",
			966 => x"ff5a0f45",
			967 => x"0c001f04",
			968 => x"008e0f45",
			969 => x"ffe60f45",
			970 => x"02013708",
			971 => x"0b001d04",
			972 => x"00020f45",
			973 => x"ff1c0f45",
			974 => x"03002e04",
			975 => x"004e0f45",
			976 => x"ff8b0f45",
			977 => x"08002030",
			978 => x"02013f2c",
			979 => x"06009e20",
			980 => x"0e006f0c",
			981 => x"0b001308",
			982 => x"0b001204",
			983 => x"fff01039",
			984 => x"001e1039",
			985 => x"ffab1039",
			986 => x"06009a0c",
			987 => x"0a002a04",
			988 => x"004c1039",
			989 => x"0b001704",
			990 => x"fff41039",
			991 => x"00041039",
			992 => x"0f00b704",
			993 => x"ffdc1039",
			994 => x"00151039",
			995 => x"04002608",
			996 => x"07002a04",
			997 => x"00061039",
			998 => x"ff3b1039",
			999 => x"000b1039",
			1000 => x"001a1039",
			1001 => x"0b001b1c",
			1002 => x"02011c10",
			1003 => x"0600a00c",
			1004 => x"04002508",
			1005 => x"05002704",
			1006 => x"ffed1039",
			1007 => x"006b1039",
			1008 => x"ffba1039",
			1009 => x"ff791039",
			1010 => x"05003908",
			1011 => x"0d001904",
			1012 => x"000c1039",
			1013 => x"00a51039",
			1014 => x"00041039",
			1015 => x"0e009110",
			1016 => x"03002a08",
			1017 => x"08002704",
			1018 => x"ffe91039",
			1019 => x"00311039",
			1020 => x"0a005b04",
			1021 => x"ff4f1039",
			1022 => x"00091039",
			1023 => x"0e009508",
			1024 => x"0a003804",
			1025 => x"00811039",
			1026 => x"fffa1039",
			1027 => x"0100170c",
			1028 => x"0c001e04",
			1029 => x"ffbe1039",
			1030 => x"01001604",
			1031 => x"ffe81039",
			1032 => x"006f1039",
			1033 => x"01001a04",
			1034 => x"ff751039",
			1035 => x"09002b04",
			1036 => x"00211039",
			1037 => x"ffe11039",
			1038 => x"0200b704",
			1039 => x"fec310d5",
			1040 => x"0500392c",
			1041 => x"04002824",
			1042 => x"0d001f1c",
			1043 => x"0d001a10",
			1044 => x"0c001808",
			1045 => x"0d001204",
			1046 => x"ff0210d5",
			1047 => x"006510d5",
			1048 => x"06009f04",
			1049 => x"004310d5",
			1050 => x"fef210d5",
			1051 => x"03002f08",
			1052 => x"03002d04",
			1053 => x"00a110d5",
			1054 => x"ff1710d5",
			1055 => x"013410d5",
			1056 => x"08002d04",
			1057 => x"fe9a10d5",
			1058 => x"005c10d5",
			1059 => x"0600af04",
			1060 => x"000810d5",
			1061 => x"013510d5",
			1062 => x"0a004318",
			1063 => x"0c001908",
			1064 => x"00012404",
			1065 => x"ff8b10d5",
			1066 => x"00a010d5",
			1067 => x"0a003404",
			1068 => x"005e10d5",
			1069 => x"08002308",
			1070 => x"04003304",
			1071 => x"000b10d5",
			1072 => x"ff4710d5",
			1073 => x"fe8710d5",
			1074 => x"00012b04",
			1075 => x"ff7510d5",
			1076 => x"011410d5",
			1077 => x"02012640",
			1078 => x"03003234",
			1079 => x"0a002d1c",
			1080 => x"08002614",
			1081 => x"09001c10",
			1082 => x"0b001508",
			1083 => x"0f00ae04",
			1084 => x"ffd011c1",
			1085 => x"000111c1",
			1086 => x"04001804",
			1087 => x"fff611c1",
			1088 => x"003211c1",
			1089 => x"ff8011c1",
			1090 => x"08002704",
			1091 => x"002f11c1",
			1092 => x"fff811c1",
			1093 => x"08002610",
			1094 => x"0e00930c",
			1095 => x"00012a08",
			1096 => x"06007404",
			1097 => x"ffe911c1",
			1098 => x"009011c1",
			1099 => x"fff211c1",
			1100 => x"ffd111c1",
			1101 => x"0a003704",
			1102 => x"ff9c11c1",
			1103 => x"001b11c1",
			1104 => x"03004404",
			1105 => x"ff6a11c1",
			1106 => x"05005004",
			1107 => x"001011c1",
			1108 => x"fff311c1",
			1109 => x"0600ac14",
			1110 => x"07003210",
			1111 => x"0c001504",
			1112 => x"003e11c1",
			1113 => x"0600a404",
			1114 => x"fffe11c1",
			1115 => x"05002d04",
			1116 => x"fffe11c1",
			1117 => x"ffb511c1",
			1118 => x"00b211c1",
			1119 => x"02013008",
			1120 => x"0c001804",
			1121 => x"fffe11c1",
			1122 => x"ff8611c1",
			1123 => x"0a002c04",
			1124 => x"ffa911c1",
			1125 => x"03002e08",
			1126 => x"0f00d204",
			1127 => x"ffdd11c1",
			1128 => x"009511c1",
			1129 => x"0a003708",
			1130 => x"0c001b04",
			1131 => x"000111c1",
			1132 => x"ff8611c1",
			1133 => x"0600b904",
			1134 => x"006211c1",
			1135 => x"ffe411c1",
			1136 => x"01000e34",
			1137 => x"0b001530",
			1138 => x"05002710",
			1139 => x"03002108",
			1140 => x"0e007e04",
			1141 => x"fff712c5",
			1142 => x"002212c5",
			1143 => x"0e009e04",
			1144 => x"ff7912c5",
			1145 => x"000112c5",
			1146 => x"0a002f10",
			1147 => x"0a002c08",
			1148 => x"0e006f04",
			1149 => x"ffd912c5",
			1150 => x"000e12c5",
			1151 => x"08001b04",
			1152 => x"fffa12c5",
			1153 => x"009312c5",
			1154 => x"03002d08",
			1155 => x"05002e04",
			1156 => x"000812c5",
			1157 => x"ffb112c5",
			1158 => x"02012904",
			1159 => x"ffee12c5",
			1160 => x"003612c5",
			1161 => x"ff5a12c5",
			1162 => x"0b001b28",
			1163 => x"0d001a20",
			1164 => x"0b001814",
			1165 => x"05002404",
			1166 => x"ffc912c5",
			1167 => x"03002708",
			1168 => x"06006704",
			1169 => x"fffc12c5",
			1170 => x"00a412c5",
			1171 => x"03002d04",
			1172 => x"ffd112c5",
			1173 => x"004f12c5",
			1174 => x"0e008508",
			1175 => x"09002204",
			1176 => x"ffc812c5",
			1177 => x"006612c5",
			1178 => x"ff7b12c5",
			1179 => x"00013204",
			1180 => x"001812c5",
			1181 => x"00c812c5",
			1182 => x"0d001d10",
			1183 => x"0001460c",
			1184 => x"08002308",
			1185 => x"08002204",
			1186 => x"ffd912c5",
			1187 => x"002c12c5",
			1188 => x"ff4612c5",
			1189 => x"003212c5",
			1190 => x"0600b610",
			1191 => x"0f00c308",
			1192 => x"05006304",
			1193 => x"ff8f12c5",
			1194 => x"001f12c5",
			1195 => x"0e009704",
			1196 => x"009912c5",
			1197 => x"fff412c5",
			1198 => x"09002904",
			1199 => x"000812c5",
			1200 => x"ff6712c5",
			1201 => x"08001c04",
			1202 => x"fe661349",
			1203 => x"0f008004",
			1204 => x"fe6f1349",
			1205 => x"0b001718",
			1206 => x"04001808",
			1207 => x"0d001404",
			1208 => x"00a91349",
			1209 => x"fedb1349",
			1210 => x"05002e08",
			1211 => x"07003104",
			1212 => x"020c1349",
			1213 => x"00d41349",
			1214 => x"0a003404",
			1215 => x"ff5f1349",
			1216 => x"01a31349",
			1217 => x"08002210",
			1218 => x"0a004f0c",
			1219 => x"06009a08",
			1220 => x"0e007a04",
			1221 => x"feaf1349",
			1222 => x"00701349",
			1223 => x"fe281349",
			1224 => x"012a1349",
			1225 => x"0d002210",
			1226 => x"00013508",
			1227 => x"00012c04",
			1228 => x"009b1349",
			1229 => x"fe301349",
			1230 => x"01001904",
			1231 => x"01341349",
			1232 => x"fe6e1349",
			1233 => x"fe5f1349",
			1234 => x"01000e34",
			1235 => x"0b001530",
			1236 => x"05002710",
			1237 => x"03002108",
			1238 => x"0e007e04",
			1239 => x"fff7145d",
			1240 => x"0020145d",
			1241 => x"0e009e04",
			1242 => x"ff7f145d",
			1243 => x"0002145d",
			1244 => x"0a002f10",
			1245 => x"0a002c08",
			1246 => x"0e006f04",
			1247 => x"ffdb145d",
			1248 => x"000e145d",
			1249 => x"08001b04",
			1250 => x"fffa145d",
			1251 => x"008e145d",
			1252 => x"03002d08",
			1253 => x"05002e04",
			1254 => x"0008145d",
			1255 => x"ffb4145d",
			1256 => x"02012904",
			1257 => x"ffee145d",
			1258 => x"0034145d",
			1259 => x"ff5f145d",
			1260 => x"0b001b28",
			1261 => x"0400251c",
			1262 => x"04001e10",
			1263 => x"0c001708",
			1264 => x"05002404",
			1265 => x"ffdc145d",
			1266 => x"0083145d",
			1267 => x"04001704",
			1268 => x"000e145d",
			1269 => x"ff8d145d",
			1270 => x"0f00ab04",
			1271 => x"ffbd145d",
			1272 => x"0d001804",
			1273 => x"0014145d",
			1274 => x"00d6145d",
			1275 => x"03003808",
			1276 => x"0e008504",
			1277 => x"0039145d",
			1278 => x"ff99145d",
			1279 => x"0059145d",
			1280 => x"03002a10",
			1281 => x"0d001f0c",
			1282 => x"0d001c08",
			1283 => x"0d001b04",
			1284 => x"000e145d",
			1285 => x"ffd7145d",
			1286 => x"009b145d",
			1287 => x"ffa1145d",
			1288 => x"0d002010",
			1289 => x"0001480c",
			1290 => x"08002308",
			1291 => x"08002204",
			1292 => x"ffda145d",
			1293 => x"002b145d",
			1294 => x"ff3a145d",
			1295 => x"000e145d",
			1296 => x"0100190c",
			1297 => x"0e009708",
			1298 => x"02011a04",
			1299 => x"fff5145d",
			1300 => x"008c145d",
			1301 => x"ffde145d",
			1302 => x"ffae145d",
			1303 => x"08001c08",
			1304 => x"01000e04",
			1305 => x"fe711529",
			1306 => x"00d71529",
			1307 => x"0c001820",
			1308 => x"04002014",
			1309 => x"01001010",
			1310 => x"0b00150c",
			1311 => x"00012708",
			1312 => x"04001b04",
			1313 => x"fe7d1529",
			1314 => x"00761529",
			1315 => x"01151529",
			1316 => x"fe841529",
			1317 => x"01631529",
			1318 => x"0d001404",
			1319 => x"ffbb1529",
			1320 => x"06007404",
			1321 => x"ff241529",
			1322 => x"019a1529",
			1323 => x"01001224",
			1324 => x"05003414",
			1325 => x"0d001a0c",
			1326 => x"0b001808",
			1327 => x"09001f04",
			1328 => x"ff0c1529",
			1329 => x"007a1529",
			1330 => x"fe541529",
			1331 => x"03002904",
			1332 => x"ff071529",
			1333 => x"02601529",
			1334 => x"09001f04",
			1335 => x"ff981529",
			1336 => x"0d001b04",
			1337 => x"fe401529",
			1338 => x"0d001c04",
			1339 => x"002e1529",
			1340 => x"fef11529",
			1341 => x"04001d0c",
			1342 => x"04001608",
			1343 => x"04001504",
			1344 => x"ffb01529",
			1345 => x"00721529",
			1346 => x"fe031529",
			1347 => x"0f00b004",
			1348 => x"fe7f1529",
			1349 => x"03002904",
			1350 => x"01781529",
			1351 => x"05003304",
			1352 => x"feb61529",
			1353 => x"00b61529",
			1354 => x"02013f64",
			1355 => x"0f00cd4c",
			1356 => x"0e008e30",
			1357 => x"0c001c1c",
			1358 => x"01001010",
			1359 => x"0b001308",
			1360 => x"0d001304",
			1361 => x"ff3c1605",
			1362 => x"01501605",
			1363 => x"05003404",
			1364 => x"ff9c1605",
			1365 => x"fe821605",
			1366 => x"0f00bc08",
			1367 => x"0f00aa04",
			1368 => x"ffe81605",
			1369 => x"01821605",
			1370 => x"ffbb1605",
			1371 => x"0300460c",
			1372 => x"08002308",
			1373 => x"07003304",
			1374 => x"ff281605",
			1375 => x"00df1605",
			1376 => x"fe631605",
			1377 => x"04004504",
			1378 => x"01171605",
			1379 => x"ff891605",
			1380 => x"05002e08",
			1381 => x"0200ee04",
			1382 => x"ff811605",
			1383 => x"01c71605",
			1384 => x"03002f04",
			1385 => x"ff171605",
			1386 => x"03003308",
			1387 => x"01001704",
			1388 => x"01771605",
			1389 => x"ff1d1605",
			1390 => x"0600ac04",
			1391 => x"00841605",
			1392 => x"ff0c1605",
			1393 => x"0800220c",
			1394 => x"07002e04",
			1395 => x"000d1605",
			1396 => x"03002d04",
			1397 => x"fe621605",
			1398 => x"ff711605",
			1399 => x"0d001f08",
			1400 => x"05003404",
			1401 => x"ffbe1605",
			1402 => x"00f21605",
			1403 => x"fe921605",
			1404 => x"0600ca08",
			1405 => x"0e00a304",
			1406 => x"01311605",
			1407 => x"ff4e1605",
			1408 => x"ffaf1605",
			1409 => x"0f008004",
			1410 => x"fe7a16a1",
			1411 => x"0e00a544",
			1412 => x"00014730",
			1413 => x"0f00cd1c",
			1414 => x"0500340c",
			1415 => x"08001b04",
			1416 => x"fe9716a1",
			1417 => x"05002404",
			1418 => x"fea516a1",
			1419 => x"00db16a1",
			1420 => x"01001208",
			1421 => x"0c001804",
			1422 => x"008616a1",
			1423 => x"fe3c16a1",
			1424 => x"0c001c04",
			1425 => x"013516a1",
			1426 => x"ffda16a1",
			1427 => x"0600b708",
			1428 => x"0f00cf04",
			1429 => x"fe0616a1",
			1430 => x"fef416a1",
			1431 => x"07003f08",
			1432 => x"09001b04",
			1433 => x"fec616a1",
			1434 => x"01b916a1",
			1435 => x"fe8e16a1",
			1436 => x"07003308",
			1437 => x"02013f04",
			1438 => x"fec916a1",
			1439 => x"010b16a1",
			1440 => x"0c002208",
			1441 => x"05003604",
			1442 => x"01cc16a1",
			1443 => x"012216a1",
			1444 => x"feac16a1",
			1445 => x"02014704",
			1446 => x"fe6e16a1",
			1447 => x"ffea16a1",
			1448 => x"01000a04",
			1449 => x"feeb174d",
			1450 => x"05002e24",
			1451 => x"08002720",
			1452 => x"0000c704",
			1453 => x"ff42174d",
			1454 => x"08001d0c",
			1455 => x"00014208",
			1456 => x"05002504",
			1457 => x"0057174d",
			1458 => x"ff10174d",
			1459 => x"0090174d",
			1460 => x"0f00c008",
			1461 => x"0e008404",
			1462 => x"0094174d",
			1463 => x"ff3c174d",
			1464 => x"03002904",
			1465 => x"013e174d",
			1466 => x"007c174d",
			1467 => x"ff33174d",
			1468 => x"02011c14",
			1469 => x"0200fd08",
			1470 => x"0200f604",
			1471 => x"ff48174d",
			1472 => x"00f8174d",
			1473 => x"0a003604",
			1474 => x"fea2174d",
			1475 => x"04002904",
			1476 => x"009c174d",
			1477 => x"ff65174d",
			1478 => x"04002108",
			1479 => x"05003204",
			1480 => x"ffab174d",
			1481 => x"010c174d",
			1482 => x"00012c04",
			1483 => x"00bc174d",
			1484 => x"08002a08",
			1485 => x"0c001904",
			1486 => x"0083174d",
			1487 => x"ff46174d",
			1488 => x"03002d04",
			1489 => x"ff3c174d",
			1490 => x"00cc174d",
			1491 => x"0d002264",
			1492 => x"01001238",
			1493 => x"0b00130c",
			1494 => x"05002404",
			1495 => x"ff401819",
			1496 => x"08001b04",
			1497 => x"ffb61819",
			1498 => x"010c1819",
			1499 => x"08001f14",
			1500 => x"0300240c",
			1501 => x"0e007b04",
			1502 => x"ff121819",
			1503 => x"07002f04",
			1504 => x"00eb1819",
			1505 => x"ffb01819",
			1506 => x"04001504",
			1507 => x"00361819",
			1508 => x"feaf1819",
			1509 => x"0e008e10",
			1510 => x"05002e08",
			1511 => x"05002704",
			1512 => x"ff191819",
			1513 => x"00d31819",
			1514 => x"0d001a04",
			1515 => x"fe841819",
			1516 => x"00801819",
			1517 => x"0c001804",
			1518 => x"01211819",
			1519 => x"00081819",
			1520 => x"07003710",
			1521 => x"09002108",
			1522 => x"05002d04",
			1523 => x"00601819",
			1524 => x"ffbf1819",
			1525 => x"0f00b004",
			1526 => x"ff441819",
			1527 => x"015b1819",
			1528 => x"07003904",
			1529 => x"ff301819",
			1530 => x"0500380c",
			1531 => x"05003304",
			1532 => x"ffde1819",
			1533 => x"01001704",
			1534 => x"014a1819",
			1535 => x"ffcb1819",
			1536 => x"03003b08",
			1537 => x"01001804",
			1538 => x"feac1819",
			1539 => x"ffe41819",
			1540 => x"00701819",
			1541 => x"fece1819",
			1542 => x"0201495c",
			1543 => x"0600bb4c",
			1544 => x"0c00181c",
			1545 => x"08001d10",
			1546 => x"0b001308",
			1547 => x"09001a04",
			1548 => x"ffcd18d5",
			1549 => x"005e18d5",
			1550 => x"07003304",
			1551 => x"ff6918d5",
			1552 => x"002018d5",
			1553 => x"0000c704",
			1554 => x"ffb618d5",
			1555 => x"0f00c904",
			1556 => x"00ac18d5",
			1557 => x"000218d5",
			1558 => x"0a003b20",
			1559 => x"07003910",
			1560 => x"00012a08",
			1561 => x"00012104",
			1562 => x"ffa918d5",
			1563 => x"004718d5",
			1564 => x"08002404",
			1565 => x"ff1518d5",
			1566 => x"ffd018d5",
			1567 => x"08002708",
			1568 => x"0e009104",
			1569 => x"000218d5",
			1570 => x"007e18d5",
			1571 => x"08002d04",
			1572 => x"ff5a18d5",
			1573 => x"004f18d5",
			1574 => x"00013a0c",
			1575 => x"0f00bb08",
			1576 => x"02011704",
			1577 => x"ffd218d5",
			1578 => x"006c18d5",
			1579 => x"ff9b18d5",
			1580 => x"009d18d5",
			1581 => x"0f00d404",
			1582 => x"fff718d5",
			1583 => x"01001a04",
			1584 => x"ff4618d5",
			1585 => x"01001f04",
			1586 => x"000a18d5",
			1587 => x"fff018d5",
			1588 => x"007b18d5",
			1589 => x"05002714",
			1590 => x"07002908",
			1591 => x"07002804",
			1592 => x"ffe119e9",
			1593 => x"003319e9",
			1594 => x"04001e08",
			1595 => x"0e00a104",
			1596 => x"ff5c19e9",
			1597 => x"fffa19e9",
			1598 => x"000319e9",
			1599 => x"0c001824",
			1600 => x"02011b18",
			1601 => x"07002f14",
			1602 => x"08001f10",
			1603 => x"0000c008",
			1604 => x"02009a04",
			1605 => x"fff919e9",
			1606 => x"002f19e9",
			1607 => x"0e007c04",
			1608 => x"ffb019e9",
			1609 => x"000219e9",
			1610 => x"009019e9",
			1611 => x"ff9b19e9",
			1612 => x"08001c04",
			1613 => x"ffdf19e9",
			1614 => x"0600a904",
			1615 => x"001619e9",
			1616 => x"00c419e9",
			1617 => x"0d001a20",
			1618 => x"0b001608",
			1619 => x"03003204",
			1620 => x"004219e9",
			1621 => x"fff519e9",
			1622 => x"0a003708",
			1623 => x"09001e04",
			1624 => x"000619e9",
			1625 => x"ff4a19e9",
			1626 => x"0b001808",
			1627 => x"09001f04",
			1628 => x"fff919e9",
			1629 => x"003719e9",
			1630 => x"0a004f04",
			1631 => x"ffcf19e9",
			1632 => x"001419e9",
			1633 => x"02013720",
			1634 => x"0f00c510",
			1635 => x"0f00c108",
			1636 => x"0200fd04",
			1637 => x"005319e9",
			1638 => x"ffb419e9",
			1639 => x"07003e04",
			1640 => x"008b19e9",
			1641 => x"fff419e9",
			1642 => x"03003108",
			1643 => x"0600bc04",
			1644 => x"ff5b19e9",
			1645 => x"001719e9",
			1646 => x"00013c04",
			1647 => x"ffe319e9",
			1648 => x"005519e9",
			1649 => x"01001908",
			1650 => x"07004004",
			1651 => x"00c919e9",
			1652 => x"ffff19e9",
			1653 => x"0f00e208",
			1654 => x"0f00da04",
			1655 => x"fff819e9",
			1656 => x"ffad19e9",
			1657 => x"000e19e9",
			1658 => x"01000a04",
			1659 => x"fee21abf",
			1660 => x"05002e24",
			1661 => x"08002720",
			1662 => x"0000c704",
			1663 => x"ff381abf",
			1664 => x"08001d0c",
			1665 => x"07002c04",
			1666 => x"00821abf",
			1667 => x"0a002f04",
			1668 => x"ff2c1abf",
			1669 => x"00011abf",
			1670 => x"0f00c008",
			1671 => x"0e008404",
			1672 => x"00a61abf",
			1673 => x"ff301abf",
			1674 => x"03002904",
			1675 => x"014c1abf",
			1676 => x"00831abf",
			1677 => x"ff281abf",
			1678 => x"08002010",
			1679 => x"0c001604",
			1680 => x"00351abf",
			1681 => x"05003804",
			1682 => x"feb51abf",
			1683 => x"05004504",
			1684 => x"00351abf",
			1685 => x"ffd91abf",
			1686 => x"02012b1c",
			1687 => x"0c001c0c",
			1688 => x"08002304",
			1689 => x"ff6d1abf",
			1690 => x"09002304",
			1691 => x"00cf1abf",
			1692 => x"00191abf",
			1693 => x"04004108",
			1694 => x"07003704",
			1695 => x"ff811abf",
			1696 => x"fea21abf",
			1697 => x"04005404",
			1698 => x"008a1abf",
			1699 => x"ffef1abf",
			1700 => x"07003c08",
			1701 => x"0a003604",
			1702 => x"01551abf",
			1703 => x"003d1abf",
			1704 => x"05003808",
			1705 => x"01001904",
			1706 => x"00931abf",
			1707 => x"ff571abf",
			1708 => x"00015204",
			1709 => x"fef21abf",
			1710 => x"002e1abf",
			1711 => x"06009510",
			1712 => x"0f008004",
			1713 => x"fe621b41",
			1714 => x"0000d708",
			1715 => x"05002704",
			1716 => x"fe651b41",
			1717 => x"03e31b41",
			1718 => x"fe5d1b41",
			1719 => x"01000c10",
			1720 => x"0e009308",
			1721 => x"07002904",
			1722 => x"00761b41",
			1723 => x"fe521b41",
			1724 => x"00013a04",
			1725 => x"fe8b1b41",
			1726 => x"00d21b41",
			1727 => x"05003918",
			1728 => x"09002b14",
			1729 => x"0f00b104",
			1730 => x"03661b41",
			1731 => x"00014608",
			1732 => x"08001f04",
			1733 => x"feee1b41",
			1734 => x"01621b41",
			1735 => x"0c001d04",
			1736 => x"021a1b41",
			1737 => x"03531b41",
			1738 => x"fe601b41",
			1739 => x"0a004308",
			1740 => x"07003704",
			1741 => x"00bc1b41",
			1742 => x"fe571b41",
			1743 => x"03101b41",
			1744 => x"06009514",
			1745 => x"01000b10",
			1746 => x"0d001504",
			1747 => x"ff9b1bd5",
			1748 => x"05003308",
			1749 => x"0000b004",
			1750 => x"fffa1bd5",
			1751 => x"00b61bd5",
			1752 => x"ffec1bd5",
			1753 => x"fee81bd5",
			1754 => x"0f00b30c",
			1755 => x"0b001a08",
			1756 => x"0000f304",
			1757 => x"ffc61bd5",
			1758 => x"01081bd5",
			1759 => x"ff8f1bd5",
			1760 => x"0001220c",
			1761 => x"04001a08",
			1762 => x"07003104",
			1763 => x"00331bd5",
			1764 => x"ffd81bd5",
			1765 => x"fef01bd5",
			1766 => x"07004214",
			1767 => x"08001d08",
			1768 => x"00015104",
			1769 => x"ff061bd5",
			1770 => x"00711bd5",
			1771 => x"05002d04",
			1772 => x"00d11bd5",
			1773 => x"05003304",
			1774 => x"ffb21bd5",
			1775 => x"00451bd5",
			1776 => x"04002b04",
			1777 => x"ff271bd5",
			1778 => x"00014d04",
			1779 => x"ffb81bd5",
			1780 => x"004e1bd5",
			1781 => x"08001f24",
			1782 => x"0c001618",
			1783 => x"0d001308",
			1784 => x"01000c04",
			1785 => x"fe991c79",
			1786 => x"00651c79",
			1787 => x"07002e08",
			1788 => x"0000be04",
			1789 => x"ff7d1c79",
			1790 => x"016b1c79",
			1791 => x"0f00de04",
			1792 => x"fec21c79",
			1793 => x"ffeb1c79",
			1794 => x"09001b08",
			1795 => x"0a002c04",
			1796 => x"ff301c79",
			1797 => x"01071c79",
			1798 => x"fe751c79",
			1799 => x"05002704",
			1800 => x"fea21c79",
			1801 => x"0c00180c",
			1802 => x"0000c704",
			1803 => x"ff581c79",
			1804 => x"0600ad04",
			1805 => x"014b1c79",
			1806 => x"00801c79",
			1807 => x"0500330c",
			1808 => x"0b001a04",
			1809 => x"00631c79",
			1810 => x"03002c04",
			1811 => x"ffd41c79",
			1812 => x"fe741c79",
			1813 => x"05003404",
			1814 => x"01341c79",
			1815 => x"01001208",
			1816 => x"08002604",
			1817 => x"fe9f1c79",
			1818 => x"008d1c79",
			1819 => x"08002604",
			1820 => x"00c81c79",
			1821 => x"fffc1c79",
			1822 => x"0a003b2c",
			1823 => x"0a003828",
			1824 => x"0d002124",
			1825 => x"0201441c",
			1826 => x"0a003110",
			1827 => x"0d001b08",
			1828 => x"0d001604",
			1829 => x"ff7c1cfd",
			1830 => x"00411cfd",
			1831 => x"05002904",
			1832 => x"00531cfd",
			1833 => x"fee81cfd",
			1834 => x"03002904",
			1835 => x"01101cfd",
			1836 => x"02011804",
			1837 => x"ff2c1cfd",
			1838 => x"002b1cfd",
			1839 => x"0600ca04",
			1840 => x"010f1cfd",
			1841 => x"00241cfd",
			1842 => x"fed11cfd",
			1843 => x"febf1cfd",
			1844 => x"05003f08",
			1845 => x"0e008b04",
			1846 => x"ffd21cfd",
			1847 => x"01471cfd",
			1848 => x"0a004304",
			1849 => x"fef91cfd",
			1850 => x"0b001f08",
			1851 => x"08002004",
			1852 => x"ffd41cfd",
			1853 => x"00fc1cfd",
			1854 => x"ffa31cfd",
			1855 => x"02012e34",
			1856 => x"06009514",
			1857 => x"0f008004",
			1858 => x"cc671da1",
			1859 => x"0e006804",
			1860 => x"d2c41da1",
			1861 => x"0000d508",
			1862 => x"0e007204",
			1863 => x"ceb91da1",
			1864 => x"cc761da1",
			1865 => x"cc6a1da1",
			1866 => x"01000c04",
			1867 => x"cc6a1da1",
			1868 => x"06009d04",
			1869 => x"dac31da1",
			1870 => x"09002710",
			1871 => x"09001f08",
			1872 => x"07003004",
			1873 => x"cfc21da1",
			1874 => x"cc721da1",
			1875 => x"05003804",
			1876 => x"d7c61da1",
			1877 => x"cfe41da1",
			1878 => x"03003a04",
			1879 => x"cc6b1da1",
			1880 => x"ce991da1",
			1881 => x"07004018",
			1882 => x"08001c04",
			1883 => x"cc6d1da1",
			1884 => x"02013a0c",
			1885 => x"0c001804",
			1886 => x"e3721da1",
			1887 => x"01001404",
			1888 => x"d0421da1",
			1889 => x"dccc1da1",
			1890 => x"04002504",
			1891 => x"eba51da1",
			1892 => x"dc511da1",
			1893 => x"05003504",
			1894 => x"cfc21da1",
			1895 => x"cc6e1da1",
			1896 => x"01000c20",
			1897 => x"0f008108",
			1898 => x"06007304",
			1899 => x"ffd91e65",
			1900 => x"00531e65",
			1901 => x"0e009e14",
			1902 => x"0300230c",
			1903 => x"07002c08",
			1904 => x"03001f04",
			1905 => x"fff61e65",
			1906 => x"002e1e65",
			1907 => x"ffee1e65",
			1908 => x"07003704",
			1909 => x"ff041e65",
			1910 => x"fff81e65",
			1911 => x"00221e65",
			1912 => x"07003f30",
			1913 => x"0a003b1c",
			1914 => x"05003914",
			1915 => x"0d002110",
			1916 => x"08001d08",
			1917 => x"0b001304",
			1918 => x"002f1e65",
			1919 => x"ff681e65",
			1920 => x"0600b704",
			1921 => x"00311e65",
			1922 => x"00c51e65",
			1923 => x"ff6d1e65",
			1924 => x"07003004",
			1925 => x"00171e65",
			1926 => x"ff2b1e65",
			1927 => x"09002608",
			1928 => x"01001204",
			1929 => x"ffe71e65",
			1930 => x"00df1e65",
			1931 => x"0c002208",
			1932 => x"05005d04",
			1933 => x"ff6a1e65",
			1934 => x"00161e65",
			1935 => x"00971e65",
			1936 => x"0c002108",
			1937 => x"0f00d004",
			1938 => x"00091e65",
			1939 => x"ff2d1e65",
			1940 => x"0600c104",
			1941 => x"ffb21e65",
			1942 => x"03003104",
			1943 => x"00591e65",
			1944 => x"ffdc1e65",
			1945 => x"00013c3c",
			1946 => x"08001f14",
			1947 => x"0b001310",
			1948 => x"0c001304",
			1949 => x"ffd91f11",
			1950 => x"0b001204",
			1951 => x"fff71f11",
			1952 => x"01000704",
			1953 => x"fffb1f11",
			1954 => x"00551f11",
			1955 => x"ff5b1f11",
			1956 => x"0c001c18",
			1957 => x"0b001b14",
			1958 => x"0000d308",
			1959 => x"03002104",
			1960 => x"00251f11",
			1961 => x"ffad1f11",
			1962 => x"05003708",
			1963 => x"05002c04",
			1964 => x"fff51f11",
			1965 => x"009e1f11",
			1966 => x"fff21f11",
			1967 => x"ffb61f11",
			1968 => x"00012608",
			1969 => x"0f00bc04",
			1970 => x"ffa11f11",
			1971 => x"007d1f11",
			1972 => x"0600a904",
			1973 => x"00191f11",
			1974 => x"ff3d1f11",
			1975 => x"09002b18",
			1976 => x"01000a04",
			1977 => x"ffc11f11",
			1978 => x"0e00a510",
			1979 => x"08002008",
			1980 => x"0e009304",
			1981 => x"ffd81f11",
			1982 => x"00561f11",
			1983 => x"01001904",
			1984 => x"00991f11",
			1985 => x"00021f11",
			1986 => x"ffe11f11",
			1987 => x"ffa21f11",
			1988 => x"0f00a910",
			1989 => x"0f008004",
			1990 => x"fe641f95",
			1991 => x"0000d708",
			1992 => x"0d001504",
			1993 => x"fe601f95",
			1994 => x"02491f95",
			1995 => x"fe5f1f95",
			1996 => x"08001b04",
			1997 => x"fe681f95",
			1998 => x"0d002128",
			1999 => x"02013714",
			2000 => x"02013110",
			2001 => x"08001f08",
			2002 => x"0b001304",
			2003 => x"03171f95",
			2004 => x"fe581f95",
			2005 => x"0c001c04",
			2006 => x"01e41f95",
			2007 => x"00481f95",
			2008 => x"ff321f95",
			2009 => x"0800240c",
			2010 => x"0c001908",
			2011 => x"0a003104",
			2012 => x"01351f95",
			2013 => x"02551f95",
			2014 => x"ffc51f95",
			2015 => x"03003104",
			2016 => x"02e51f95",
			2017 => x"01701f95",
			2018 => x"01001804",
			2019 => x"00921f95",
			2020 => x"fe4e1f95",
			2021 => x"05002718",
			2022 => x"07002908",
			2023 => x"03002404",
			2024 => x"fff22069",
			2025 => x"00172069",
			2026 => x"03002108",
			2027 => x"03001f04",
			2028 => x"fff42069",
			2029 => x"00162069",
			2030 => x"0e00a104",
			2031 => x"ff802069",
			2032 => x"00052069",
			2033 => x"0c001824",
			2034 => x"02011b18",
			2035 => x"07002f10",
			2036 => x"08001d08",
			2037 => x"0000c004",
			2038 => x"00152069",
			2039 => x"ffcc2069",
			2040 => x"04002004",
			2041 => x"00522069",
			2042 => x"fffa2069",
			2043 => x"04001d04",
			2044 => x"00052069",
			2045 => x"ffb52069",
			2046 => x"01000a04",
			2047 => x"ffd82069",
			2048 => x"0600a904",
			2049 => x"000a2069",
			2050 => x"008b2069",
			2051 => x"0d001a10",
			2052 => x"01001208",
			2053 => x"0b001604",
			2054 => x"001e2069",
			2055 => x"ff572069",
			2056 => x"00013104",
			2057 => x"00462069",
			2058 => x"ffe92069",
			2059 => x"0b001b08",
			2060 => x"0a003804",
			2061 => x"006c2069",
			2062 => x"00032069",
			2063 => x"0c001e08",
			2064 => x"02013904",
			2065 => x"ff782069",
			2066 => x"00062069",
			2067 => x"01001708",
			2068 => x"05003804",
			2069 => x"00822069",
			2070 => x"ffe42069",
			2071 => x"0e009504",
			2072 => x"00172069",
			2073 => x"ffa92069",
			2074 => x"02012634",
			2075 => x"0f00b820",
			2076 => x"0f00a910",
			2077 => x"06007f0c",
			2078 => x"0f008004",
			2079 => x"ffca214d",
			2080 => x"05003404",
			2081 => x"0047214d",
			2082 => x"ffe7214d",
			2083 => x"ffa1214d",
			2084 => x"0b001b0c",
			2085 => x"01000e08",
			2086 => x"00010604",
			2087 => x"000c214d",
			2088 => x"ffd7214d",
			2089 => x"0090214d",
			2090 => x"ffc4214d",
			2091 => x"0b001c0c",
			2092 => x"04001908",
			2093 => x"07003004",
			2094 => x"0023214d",
			2095 => x"ffe6214d",
			2096 => x"ff49214d",
			2097 => x"00012604",
			2098 => x"0067214d",
			2099 => x"ffb3214d",
			2100 => x"0f00cd1c",
			2101 => x"0600a608",
			2102 => x"00013a04",
			2103 => x"ffb5214d",
			2104 => x"0020214d",
			2105 => x"04001e04",
			2106 => x"fff3214d",
			2107 => x"05003404",
			2108 => x"00a8214d",
			2109 => x"01001004",
			2110 => x"ffc8214d",
			2111 => x"01001704",
			2112 => x"0060214d",
			2113 => x"ffef214d",
			2114 => x"0201491c",
			2115 => x"0500330c",
			2116 => x"04002208",
			2117 => x"07002f04",
			2118 => x"fff8214d",
			2119 => x"ff81214d",
			2120 => x"000e214d",
			2121 => x"0d00210c",
			2122 => x"05003804",
			2123 => x"0067214d",
			2124 => x"09002704",
			2125 => x"fffe214d",
			2126 => x"ffba214d",
			2127 => x"ffae214d",
			2128 => x"07003d04",
			2129 => x"0058214d",
			2130 => x"0003214d",
			2131 => x"08001f28",
			2132 => x"0c00161c",
			2133 => x"0600990c",
			2134 => x"07002804",
			2135 => x"feff2201",
			2136 => x"05002404",
			2137 => x"ff752201",
			2138 => x"01a22201",
			2139 => x"0001510c",
			2140 => x"05003108",
			2141 => x"07002904",
			2142 => x"00302201",
			2143 => x"fe862201",
			2144 => x"00702201",
			2145 => x"008b2201",
			2146 => x"09001b08",
			2147 => x"0a002c04",
			2148 => x"ff292201",
			2149 => x"011b2201",
			2150 => x"fe712201",
			2151 => x"05002704",
			2152 => x"fe992201",
			2153 => x"0c00180c",
			2154 => x"0000c704",
			2155 => x"ff4e2201",
			2156 => x"0600ad04",
			2157 => x"015a2201",
			2158 => x"008e2201",
			2159 => x"05003310",
			2160 => x"0001460c",
			2161 => x"0200fd04",
			2162 => x"010b2201",
			2163 => x"03002904",
			2164 => x"ff4a2201",
			2165 => x"fe872201",
			2166 => x"00c52201",
			2167 => x"05003404",
			2168 => x"01472201",
			2169 => x"01001208",
			2170 => x"08002604",
			2171 => x"fe8d2201",
			2172 => x"00982201",
			2173 => x"0d001b04",
			2174 => x"01152201",
			2175 => x"00292201",
			2176 => x"00011f20",
			2177 => x"0f008c0c",
			2178 => x"0f008004",
			2179 => x"fe6122a5",
			2180 => x"08002204",
			2181 => x"fe5122a5",
			2182 => x"016422a5",
			2183 => x"0f008f04",
			2184 => x"04ad22a5",
			2185 => x"07002f08",
			2186 => x"09001d04",
			2187 => x"fe6622a5",
			2188 => x"028722a5",
			2189 => x"01001604",
			2190 => x"fe5322a5",
			2191 => x"ff8922a5",
			2192 => x"08001c04",
			2193 => x"fe6222a5",
			2194 => x"0d002128",
			2195 => x"00014614",
			2196 => x"03003810",
			2197 => x"0a003808",
			2198 => x"08001f04",
			2199 => x"ffce22a5",
			2200 => x"018422a5",
			2201 => x"01001604",
			2202 => x"fe3b22a5",
			2203 => x"ffd722a5",
			2204 => x"039f22a5",
			2205 => x"0e00a510",
			2206 => x"08002408",
			2207 => x"05003004",
			2208 => x"022e22a5",
			2209 => x"018822a5",
			2210 => x"05003504",
			2211 => x"03e722a5",
			2212 => x"024922a5",
			2213 => x"007122a5",
			2214 => x"01001804",
			2215 => x"00bb22a5",
			2216 => x"fe5222a5",
			2217 => x"0f008004",
			2218 => x"fe922301",
			2219 => x"0d002128",
			2220 => x"0d002020",
			2221 => x"0d001f1c",
			2222 => x"01000e0c",
			2223 => x"0b001608",
			2224 => x"08001c04",
			2225 => x"fe8c2301",
			2226 => x"00972301",
			2227 => x"fe702301",
			2228 => x"04002108",
			2229 => x"04001b04",
			2230 => x"00272301",
			2231 => x"011e2301",
			2232 => x"07003404",
			2233 => x"00d32301",
			2234 => x"ffb42301",
			2235 => x"fe772301",
			2236 => x"07003d04",
			2237 => x"ff432301",
			2238 => x"01892301",
			2239 => x"fe8e2301",
			2240 => x"0f00a90c",
			2241 => x"0f008004",
			2242 => x"fe5d238d",
			2243 => x"07002a04",
			2244 => x"0076238d",
			2245 => x"fe5b238d",
			2246 => x"08001c08",
			2247 => x"0f00af04",
			2248 => x"0101238d",
			2249 => x"fe5e238d",
			2250 => x"0700402c",
			2251 => x"02012614",
			2252 => x"08002710",
			2253 => x"01001008",
			2254 => x"0000fc04",
			2255 => x"0316238d",
			2256 => x"fe53238d",
			2257 => x"0d001c04",
			2258 => x"0331238d",
			2259 => x"fffb238d",
			2260 => x"fe57238d",
			2261 => x"0800200c",
			2262 => x"0b001504",
			2263 => x"0358238d",
			2264 => x"0d001704",
			2265 => x"0079238d",
			2266 => x"fe29238d",
			2267 => x"0600ac04",
			2268 => x"059d238d",
			2269 => x"08002704",
			2270 => x"0394238d",
			2271 => x"0100238d",
			2272 => x"05003504",
			2273 => x"ffee238d",
			2274 => x"fe5f238d",
			2275 => x"0d001a3c",
			2276 => x"0b001828",
			2277 => x"01000e18",
			2278 => x"0b001514",
			2279 => x"08001c04",
			2280 => x"fe992469",
			2281 => x"04001808",
			2282 => x"0600ae04",
			2283 => x"fec42469",
			2284 => x"00092469",
			2285 => x"0a002804",
			2286 => x"ff3c2469",
			2287 => x"01312469",
			2288 => x"fe732469",
			2289 => x"0e008808",
			2290 => x"0000c704",
			2291 => x"fede2469",
			2292 => x"013c2469",
			2293 => x"03002d04",
			2294 => x"fee62469",
			2295 => x"00af2469",
			2296 => x"0a004f0c",
			2297 => x"0f00b308",
			2298 => x"0e007a04",
			2299 => x"feda2469",
			2300 => x"00f12469",
			2301 => x"fe732469",
			2302 => x"07003304",
			2303 => x"00f92469",
			2304 => x"ffcb2469",
			2305 => x"0d001b0c",
			2306 => x"05003808",
			2307 => x"0a002c04",
			2308 => x"ffb42469",
			2309 => x"01f62469",
			2310 => x"003d2469",
			2311 => x"0900250c",
			2312 => x"03003108",
			2313 => x"05002e04",
			2314 => x"00fe2469",
			2315 => x"fe782469",
			2316 => x"00b32469",
			2317 => x"0e008604",
			2318 => x"fe982469",
			2319 => x"00012608",
			2320 => x"08002904",
			2321 => x"01e72469",
			2322 => x"ff2e2469",
			2323 => x"00013508",
			2324 => x"0f00be04",
			2325 => x"00172469",
			2326 => x"fe752469",
			2327 => x"0f00cd04",
			2328 => x"01842469",
			2329 => x"00422469",
			2330 => x"0a003b3c",
			2331 => x"05003a38",
			2332 => x"00014628",
			2333 => x"0f00ca1c",
			2334 => x"04002610",
			2335 => x"05003408",
			2336 => x"02012704",
			2337 => x"ffc424fd",
			2338 => x"00ab24fd",
			2339 => x"06009a04",
			2340 => x"002f24fd",
			2341 => x"fef824fd",
			2342 => x"08002608",
			2343 => x"04002a04",
			2344 => x"00f224fd",
			2345 => x"ffc824fd",
			2346 => x"ff4324fd",
			2347 => x"0a003104",
			2348 => x"ff1b24fd",
			2349 => x"02013004",
			2350 => x"ff4d24fd",
			2351 => x"002a24fd",
			2352 => x"0d001f0c",
			2353 => x"08002008",
			2354 => x"02013f04",
			2355 => x"ff7724fd",
			2356 => x"006924fd",
			2357 => x"010624fd",
			2358 => x"ff9d24fd",
			2359 => x"ff2224fd",
			2360 => x"0600b70c",
			2361 => x"00012a04",
			2362 => x"ffa724fd",
			2363 => x"01001704",
			2364 => x"00ef24fd",
			2365 => x"ffec24fd",
			2366 => x"ffa624fd",
			2367 => x"0e009c4c",
			2368 => x"04002628",
			2369 => x"04002424",
			2370 => x"0d001f20",
			2371 => x"01000c10",
			2372 => x"0f008108",
			2373 => x"03002904",
			2374 => x"ffed25b9",
			2375 => x"004425b9",
			2376 => x"0e009304",
			2377 => x"ff5325b9",
			2378 => x"001e25b9",
			2379 => x"0e008e08",
			2380 => x"06009e04",
			2381 => x"009425b9",
			2382 => x"ffb125b9",
			2383 => x"0e009404",
			2384 => x"00c525b9",
			2385 => x"000225b9",
			2386 => x"ff6225b9",
			2387 => x"ff4325b9",
			2388 => x"08002614",
			2389 => x"02011808",
			2390 => x"05003504",
			2391 => x"004b25b9",
			2392 => x"ff8d25b9",
			2393 => x"09002108",
			2394 => x"03003304",
			2395 => x"007c25b9",
			2396 => x"ff9d25b9",
			2397 => x"00fd25b9",
			2398 => x"0d002004",
			2399 => x"ff3f25b9",
			2400 => x"08002a04",
			2401 => x"ffdb25b9",
			2402 => x"00013404",
			2403 => x"fff425b9",
			2404 => x"00c625b9",
			2405 => x"01001a0c",
			2406 => x"0f00d404",
			2407 => x"001225b9",
			2408 => x"02014704",
			2409 => x"ff4825b9",
			2410 => x"ffd925b9",
			2411 => x"03002e04",
			2412 => x"003925b9",
			2413 => x"ffe525b9",
			2414 => x"0a002c08",
			2415 => x"02013904",
			2416 => x"ff91266d",
			2417 => x"0012266d",
			2418 => x"05002e1c",
			2419 => x"08001d10",
			2420 => x"05002708",
			2421 => x"0e009404",
			2422 => x"0002266d",
			2423 => x"ffcf266d",
			2424 => x"00014204",
			2425 => x"ffee266d",
			2426 => x"0021266d",
			2427 => x"03002e08",
			2428 => x"0000d604",
			2429 => x"fffb266d",
			2430 => x"0086266d",
			2431 => x"fff2266d",
			2432 => x"0d001a18",
			2433 => x"01001210",
			2434 => x"0c00180c",
			2435 => x"0f00c808",
			2436 => x"0f00c204",
			2437 => x"ffe0266d",
			2438 => x"004c266d",
			2439 => x"ffde266d",
			2440 => x"ff6e266d",
			2441 => x"0e008504",
			2442 => x"004a266d",
			2443 => x"ffe9266d",
			2444 => x"01001718",
			2445 => x"05003808",
			2446 => x"05003304",
			2447 => x"0001266d",
			2448 => x"007a266d",
			2449 => x"0a004308",
			2450 => x"08002404",
			2451 => x"002e266d",
			2452 => x"ff98266d",
			2453 => x"07004004",
			2454 => x"004b266d",
			2455 => x"fffa266d",
			2456 => x"0d001f04",
			2457 => x"001d266d",
			2458 => x"ff7f266d",
			2459 => x"07004054",
			2460 => x"0600a730",
			2461 => x"0f00b81c",
			2462 => x"0b001b18",
			2463 => x"0600950c",
			2464 => x"06007f08",
			2465 => x"07002904",
			2466 => x"ff942731",
			2467 => x"00922731",
			2468 => x"ff072731",
			2469 => x"01000e08",
			2470 => x"0000ff04",
			2471 => x"00452731",
			2472 => x"ff5c2731",
			2473 => x"01262731",
			2474 => x"ff092731",
			2475 => x"0c001508",
			2476 => x"00013404",
			2477 => x"ffe82731",
			2478 => x"00812731",
			2479 => x"04001d04",
			2480 => x"ffdf2731",
			2481 => x"04002804",
			2482 => x"feb82731",
			2483 => x"ffae2731",
			2484 => x"0600aa08",
			2485 => x"00013304",
			2486 => x"ffd12731",
			2487 => x"01302731",
			2488 => x"0e008e0c",
			2489 => x"0600ac04",
			2490 => x"007e2731",
			2491 => x"07002e04",
			2492 => x"00442731",
			2493 => x"fefd2731",
			2494 => x"04002c0c",
			2495 => x"04002808",
			2496 => x"04002304",
			2497 => x"006d2731",
			2498 => x"ff9b2731",
			2499 => x"00ed2731",
			2500 => x"ff492731",
			2501 => x"0c002104",
			2502 => x"fef02731",
			2503 => x"00014904",
			2504 => x"ff7e2731",
			2505 => x"02014104",
			2506 => x"00b42731",
			2507 => x"ffd42731",
			2508 => x"01001034",
			2509 => x"0b001520",
			2510 => x"00013c18",
			2511 => x"06009910",
			2512 => x"03002404",
			2513 => x"ffb6281d",
			2514 => x"0000be04",
			2515 => x"ffd3281d",
			2516 => x"01000704",
			2517 => x"fff9281d",
			2518 => x"009d281d",
			2519 => x"08001d04",
			2520 => x"ff62281d",
			2521 => x"0002281d",
			2522 => x"01000a04",
			2523 => x"ffab281d",
			2524 => x"00c8281d",
			2525 => x"0e008e0c",
			2526 => x"0c001608",
			2527 => x"05002a04",
			2528 => x"0022281d",
			2529 => x"ffe7281d",
			2530 => x"fef8281d",
			2531 => x"0c001804",
			2532 => x"0072281d",
			2533 => x"ff9a281d",
			2534 => x"0b001b18",
			2535 => x"0c001c14",
			2536 => x"03002d0c",
			2537 => x"0f00bc08",
			2538 => x"05002704",
			2539 => x"ffc2281d",
			2540 => x"00a0281d",
			2541 => x"ffd0281d",
			2542 => x"0b001904",
			2543 => x"004f281d",
			2544 => x"00f0281d",
			2545 => x"ffb8281d",
			2546 => x"09002508",
			2547 => x"04001d04",
			2548 => x"000d281d",
			2549 => x"ff33281d",
			2550 => x"0f00c310",
			2551 => x"0100150c",
			2552 => x"08002304",
			2553 => x"003a281d",
			2554 => x"05006304",
			2555 => x"ffca281d",
			2556 => x"002d281d",
			2557 => x"ff4d281d",
			2558 => x"09002b10",
			2559 => x"05003808",
			2560 => x"05003304",
			2561 => x"0005281d",
			2562 => x"00df281d",
			2563 => x"0c001f04",
			2564 => x"001f281d",
			2565 => x"ff89281d",
			2566 => x"ff61281d",
			2567 => x"0700404c",
			2568 => x"0f00a918",
			2569 => x"01000b0c",
			2570 => x"0b001508",
			2571 => x"03002404",
			2572 => x"fff728b9",
			2573 => x"003328b9",
			2574 => x"ffe128b9",
			2575 => x"03002108",
			2576 => x"03001d04",
			2577 => x"fff128b9",
			2578 => x"002028b9",
			2579 => x"ff7528b9",
			2580 => x"0f00cd20",
			2581 => x"00013c14",
			2582 => x"00013710",
			2583 => x"0c001c08",
			2584 => x"01000c04",
			2585 => x"ffc928b9",
			2586 => x"005a28b9",
			2587 => x"0e009104",
			2588 => x"ffa928b9",
			2589 => x"004a28b9",
			2590 => x"ffa328b9",
			2591 => x"01001008",
			2592 => x"0e008704",
			2593 => x"002d28b9",
			2594 => x"ffc528b9",
			2595 => x"00a128b9",
			2596 => x"00015710",
			2597 => x"0f00cf04",
			2598 => x"ff8628b9",
			2599 => x"04001d04",
			2600 => x"ff8a28b9",
			2601 => x"0a003404",
			2602 => x"005728b9",
			2603 => x"ffcb28b9",
			2604 => x"005d28b9",
			2605 => x"ff7928b9",
			2606 => x"02013750",
			2607 => x"0f00c538",
			2608 => x"0f00c22c",
			2609 => x"06009e18",
			2610 => x"0600950c",
			2611 => x"07002a08",
			2612 => x"07002904",
			2613 => x"ffb32985",
			2614 => x"00972985",
			2615 => x"ff2f2985",
			2616 => x"0c001c08",
			2617 => x"01000c04",
			2618 => x"ffc62985",
			2619 => x"00e62985",
			2620 => x"ff9f2985",
			2621 => x"05004810",
			2622 => x"0e008508",
			2623 => x"04002304",
			2624 => x"ff662985",
			2625 => x"00652985",
			2626 => x"07003304",
			2627 => x"ffe92985",
			2628 => x"fef22985",
			2629 => x"007c2985",
			2630 => x"04002004",
			2631 => x"ff942985",
			2632 => x"0e009304",
			2633 => x"00d42985",
			2634 => x"ffd52985",
			2635 => x"02012e04",
			2636 => x"fef02985",
			2637 => x"0800260c",
			2638 => x"00014208",
			2639 => x"0600af04",
			2640 => x"ffce2985",
			2641 => x"00c22985",
			2642 => x"ff592985",
			2643 => x"0600bb04",
			2644 => x"ff012985",
			2645 => x"000e2985",
			2646 => x"0c002214",
			2647 => x"0800220c",
			2648 => x"09001c08",
			2649 => x"08001b04",
			2650 => x"ffdf2985",
			2651 => x"00c22985",
			2652 => x"ff782985",
			2653 => x"07004004",
			2654 => x"00e72985",
			2655 => x"ffd02985",
			2656 => x"ff722985",
			2657 => x"0800275c",
			2658 => x"08001f24",
			2659 => x"02013418",
			2660 => x"0f008108",
			2661 => x"06007204",
			2662 => x"ffee2a69",
			2663 => x"001b2a69",
			2664 => x"0a002a0c",
			2665 => x"06009504",
			2666 => x"ffd52a69",
			2667 => x"06009d04",
			2668 => x"002c2a69",
			2669 => x"fff72a69",
			2670 => x"ff6c2a69",
			2671 => x"0e009a08",
			2672 => x"01000a04",
			2673 => x"fff32a69",
			2674 => x"00622a69",
			2675 => x"ffc72a69",
			2676 => x"0c00180c",
			2677 => x"05002504",
			2678 => x"ffdc2a69",
			2679 => x"0f008004",
			2680 => x"ffe72a69",
			2681 => x"00982a69",
			2682 => x"08002318",
			2683 => x"04002610",
			2684 => x"0d001b08",
			2685 => x"0600a204",
			2686 => x"00062a69",
			2687 => x"ff732a69",
			2688 => x"0d001d04",
			2689 => x"00122a69",
			2690 => x"fff52a69",
			2691 => x"00011d04",
			2692 => x"ffe62a69",
			2693 => x"004d2a69",
			2694 => x"0f00af04",
			2695 => x"ffcb2a69",
			2696 => x"0b001b08",
			2697 => x"07003704",
			2698 => x"00792a69",
			2699 => x"000f2a69",
			2700 => x"0600af04",
			2701 => x"ffbb2a69",
			2702 => x"003a2a69",
			2703 => x"04002108",
			2704 => x"08002a04",
			2705 => x"00282a69",
			2706 => x"ffd32a69",
			2707 => x"08002d08",
			2708 => x"03005304",
			2709 => x"ff5e2a69",
			2710 => x"00092a69",
			2711 => x"0e009504",
			2712 => x"00262a69",
			2713 => x"ffe52a69",
			2714 => x"05002404",
			2715 => x"feb72afd",
			2716 => x"0b00130c",
			2717 => x"08001b04",
			2718 => x"ffa92afd",
			2719 => x"0600b104",
			2720 => x"013d2afd",
			2721 => x"00542afd",
			2722 => x"08001f18",
			2723 => x"0f00d310",
			2724 => x"0500280c",
			2725 => x"06009b08",
			2726 => x"0000ce04",
			2727 => x"ffd62afd",
			2728 => x"00e82afd",
			2729 => x"ff172afd",
			2730 => x"fe832afd",
			2731 => x"0e009d04",
			2732 => x"00b32afd",
			2733 => x"ff2b2afd",
			2734 => x"0c00180c",
			2735 => x"0a002f08",
			2736 => x"03002604",
			2737 => x"013a2afd",
			2738 => x"ff3b2afd",
			2739 => x"016d2afd",
			2740 => x"0a003b0c",
			2741 => x"0a003808",
			2742 => x"0f00c004",
			2743 => x"ff5e2afd",
			2744 => x"002f2afd",
			2745 => x"fe9b2afd",
			2746 => x"0e009908",
			2747 => x"00012804",
			2748 => x"ff572afd",
			2749 => x"011d2afd",
			2750 => x"ff022afd",
			2751 => x"08002764",
			2752 => x"07003648",
			2753 => x"0c001828",
			2754 => x"0500240c",
			2755 => x"03002108",
			2756 => x"03001f04",
			2757 => x"ffe12be1",
			2758 => x"00192be1",
			2759 => x"ff792be1",
			2760 => x"05002e10",
			2761 => x"0f008c08",
			2762 => x"03002104",
			2763 => x"00362be1",
			2764 => x"ffa72be1",
			2765 => x"08001b04",
			2766 => x"ffdc2be1",
			2767 => x"00a72be1",
			2768 => x"04002004",
			2769 => x"ff852be1",
			2770 => x"0e008604",
			2771 => x"ffdb2be1",
			2772 => x"00672be1",
			2773 => x"08002310",
			2774 => x"05003808",
			2775 => x"04002604",
			2776 => x"ff092be1",
			2777 => x"00052be1",
			2778 => x"04002a04",
			2779 => x"004a2be1",
			2780 => x"ffd32be1",
			2781 => x"09002408",
			2782 => x"09002204",
			2783 => x"ffff2be1",
			2784 => x"007b2be1",
			2785 => x"0a003b04",
			2786 => x"ff912be1",
			2787 => x"000d2be1",
			2788 => x"0a00360c",
			2789 => x"0e008f04",
			2790 => x"ffed2be1",
			2791 => x"00014304",
			2792 => x"00d32be1",
			2793 => x"002d2be1",
			2794 => x"03003508",
			2795 => x"08002404",
			2796 => x"00132be1",
			2797 => x"ff612be1",
			2798 => x"0c001f04",
			2799 => x"00872be1",
			2800 => x"ffe62be1",
			2801 => x"02013708",
			2802 => x"0b001d04",
			2803 => x"00052be1",
			2804 => x"ff272be1",
			2805 => x"03002e04",
			2806 => x"004a2be1",
			2807 => x"ff8f2be1",
			2808 => x"08001c04",
			2809 => x"fe9e2c6d",
			2810 => x"00014734",
			2811 => x"0a003b24",
			2812 => x"0a003820",
			2813 => x"0f00c910",
			2814 => x"0e009008",
			2815 => x"0d001c04",
			2816 => x"003d2c6d",
			2817 => x"fe7b2c6d",
			2818 => x"00012204",
			2819 => x"ff212c6d",
			2820 => x"01702c6d",
			2821 => x"0d001c08",
			2822 => x"0600b704",
			2823 => x"fe732c6d",
			2824 => x"ffd32c6d",
			2825 => x"04002704",
			2826 => x"00ff2c6d",
			2827 => x"feae2c6d",
			2828 => x"fe852c6d",
			2829 => x"00012804",
			2830 => x"fef02c6d",
			2831 => x"00013d08",
			2832 => x"0600a904",
			2833 => x"01282c6d",
			2834 => x"fede2c6d",
			2835 => x"01832c6d",
			2836 => x"0700440c",
			2837 => x"0a003608",
			2838 => x"0a003104",
			2839 => x"00842c6d",
			2840 => x"01492c6d",
			2841 => x"ffcb2c6d",
			2842 => x"feed2c6d",
			2843 => x"0a002c1c",
			2844 => x"0000d304",
			2845 => x"fee12d39",
			2846 => x"06009908",
			2847 => x"0d001304",
			2848 => x"ff9a2d39",
			2849 => x"00d72d39",
			2850 => x"0400170c",
			2851 => x"07002e08",
			2852 => x"04001304",
			2853 => x"ff982d39",
			2854 => x"fff82d39",
			2855 => x"00512d39",
			2856 => x"fef62d39",
			2857 => x"03002a1c",
			2858 => x"01001618",
			2859 => x"00014614",
			2860 => x"07003010",
			2861 => x"00012808",
			2862 => x"06007404",
			2863 => x"ffc52d39",
			2864 => x"00d52d39",
			2865 => x"05002a04",
			2866 => x"ffd92d39",
			2867 => x"ff452d39",
			2868 => x"feb32d39",
			2869 => x"01292d39",
			2870 => x"01082d39",
			2871 => x"05003314",
			2872 => x"0b001810",
			2873 => x"0f00ce08",
			2874 => x"0d001404",
			2875 => x"ffd02d39",
			2876 => x"00cc2d39",
			2877 => x"07003404",
			2878 => x"ff392d39",
			2879 => x"00232d39",
			2880 => x"febd2d39",
			2881 => x"05003404",
			2882 => x"00fc2d39",
			2883 => x"0100120c",
			2884 => x"0e009008",
			2885 => x"0b001504",
			2886 => x"00712d39",
			2887 => x"feab2d39",
			2888 => x"003e2d39",
			2889 => x"02014008",
			2890 => x"05003804",
			2891 => x"00962d39",
			2892 => x"ffea2d39",
			2893 => x"fefb2d39",
			2894 => x"07004064",
			2895 => x"01001034",
			2896 => x"0b00151c",
			2897 => x"00013c14",
			2898 => x"0b00130c",
			2899 => x"0e009108",
			2900 => x"0000be04",
			2901 => x"ff8d2e1d",
			2902 => x"01052e1d",
			2903 => x"ff572e1d",
			2904 => x"09001d04",
			2905 => x"fecb2e1d",
			2906 => x"00632e1d",
			2907 => x"01000a04",
			2908 => x"ff362e1d",
			2909 => x"011f2e1d",
			2910 => x"0800220c",
			2911 => x"05002608",
			2912 => x"05002404",
			2913 => x"ffae2e1d",
			2914 => x"00642e1d",
			2915 => x"fe962e1d",
			2916 => x"05003408",
			2917 => x"01000e04",
			2918 => x"ff992e1d",
			2919 => x"01332e1d",
			2920 => x"fed42e1d",
			2921 => x"04001b10",
			2922 => x"0c001704",
			2923 => x"007b2e1d",
			2924 => x"04001608",
			2925 => x"04001504",
			2926 => x"fff92e1d",
			2927 => x"003b2e1d",
			2928 => x"fec52e1d",
			2929 => x"0f00ae08",
			2930 => x"08002204",
			2931 => x"00362e1d",
			2932 => x"fedc2e1d",
			2933 => x"03002c08",
			2934 => x"08002404",
			2935 => x"00432e1d",
			2936 => x"01402e1d",
			2937 => x"00012c08",
			2938 => x"08002604",
			2939 => x"012e2e1d",
			2940 => x"ff8a2e1d",
			2941 => x"02012604",
			2942 => x"fea32e1d",
			2943 => x"00252e1d",
			2944 => x"0c002104",
			2945 => x"feb02e1d",
			2946 => x"00014904",
			2947 => x"ff5d2e1d",
			2948 => x"00015004",
			2949 => x"01032e1d",
			2950 => x"ff992e1d",
			2951 => x"02013758",
			2952 => x"0f00cd48",
			2953 => x"05003424",
			2954 => x"08001f14",
			2955 => x"0b001308",
			2956 => x"08001b04",
			2957 => x"ffe72f01",
			2958 => x"003f2f01",
			2959 => x"01000e04",
			2960 => x"ff932f01",
			2961 => x"0d001504",
			2962 => x"fff02f01",
			2963 => x"00162f01",
			2964 => x"05002704",
			2965 => x"ffcd2f01",
			2966 => x"0f008004",
			2967 => x"ffe62f01",
			2968 => x"0b001904",
			2969 => x"00942f01",
			2970 => x"00182f01",
			2971 => x"0a003b18",
			2972 => x"07003d10",
			2973 => x"07003108",
			2974 => x"0e007d04",
			2975 => x"ffdb2f01",
			2976 => x"00302f01",
			2977 => x"07003904",
			2978 => x"ff4e2f01",
			2979 => x"fff22f01",
			2980 => x"0f00c404",
			2981 => x"002e2f01",
			2982 => x"fff92f01",
			2983 => x"00012804",
			2984 => x"ffdc2f01",
			2985 => x"01001704",
			2986 => x"00552f01",
			2987 => x"fff82f01",
			2988 => x"0e009a04",
			2989 => x"ff872f01",
			2990 => x"0600be08",
			2991 => x"05003804",
			2992 => x"00382f01",
			2993 => x"ffeb2f01",
			2994 => x"ffcf2f01",
			2995 => x"04002c18",
			2996 => x"0800200c",
			2997 => x"0b001508",
			2998 => x"01000a04",
			2999 => x"ffd62f01",
			3000 => x"00672f01",
			3001 => x"ff9d2f01",
			3002 => x"0b002108",
			3003 => x"07004004",
			3004 => x"00b12f01",
			3005 => x"00162f01",
			3006 => x"ffca2f01",
			3007 => x"ffcd2f01",
			3008 => x"0a002c1c",
			3009 => x"0000d304",
			3010 => x"fed82fd5",
			3011 => x"06009908",
			3012 => x"0f00aa04",
			3013 => x"ffe32fd5",
			3014 => x"010b2fd5",
			3015 => x"0400170c",
			3016 => x"07002e08",
			3017 => x"04001304",
			3018 => x"ff942fd5",
			3019 => x"fff42fd5",
			3020 => x"00502fd5",
			3021 => x"fee72fd5",
			3022 => x"03002a1c",
			3023 => x"01001618",
			3024 => x"00014614",
			3025 => x"07003010",
			3026 => x"00012808",
			3027 => x"06007404",
			3028 => x"ffc12fd5",
			3029 => x"00e22fd5",
			3030 => x"05002a04",
			3031 => x"ffd92fd5",
			3032 => x"ff3c2fd5",
			3033 => x"feac2fd5",
			3034 => x"01332fd5",
			3035 => x"011c2fd5",
			3036 => x"05003314",
			3037 => x"0b001810",
			3038 => x"0f00ce08",
			3039 => x"0d001404",
			3040 => x"ffcd2fd5",
			3041 => x"00d52fd5",
			3042 => x"07003404",
			3043 => x"ff2e2fd5",
			3044 => x"00252fd5",
			3045 => x"feb02fd5",
			3046 => x"05003404",
			3047 => x"01122fd5",
			3048 => x"01001210",
			3049 => x"0b001608",
			3050 => x"0a003404",
			3051 => x"ff3e2fd5",
			3052 => x"00f32fd5",
			3053 => x"09001e04",
			3054 => x"00562fd5",
			3055 => x"fec92fd5",
			3056 => x"02014008",
			3057 => x"05003804",
			3058 => x"00a42fd5",
			3059 => x"ffe32fd5",
			3060 => x"fef12fd5",
			3061 => x"07004060",
			3062 => x"0d001a30",
			3063 => x"0b001828",
			3064 => x"0400261c",
			3065 => x"05002e10",
			3066 => x"0200ea08",
			3067 => x"0b001504",
			3068 => x"fef830b1",
			3069 => x"005030b1",
			3070 => x"0d001204",
			3071 => x"ff9130b1",
			3072 => x"00aa30b1",
			3073 => x"03002f08",
			3074 => x"0e006304",
			3075 => x"009530b1",
			3076 => x"fedb30b1",
			3077 => x"005330b1",
			3078 => x"0e006f04",
			3079 => x"ffab30b1",
			3080 => x"01000a04",
			3081 => x"ffe030b1",
			3082 => x"010830b1",
			3083 => x"01001204",
			3084 => x"fec630b1",
			3085 => x"ffa230b1",
			3086 => x"0b001b0c",
			3087 => x"06009904",
			3088 => x"ff7430b1",
			3089 => x"0f00c404",
			3090 => x"011530b1",
			3091 => x"002730b1",
			3092 => x"03002a0c",
			3093 => x"01001608",
			3094 => x"0d001b04",
			3095 => x"001d30b1",
			3096 => x"ff7230b1",
			3097 => x"014130b1",
			3098 => x"0d00200c",
			3099 => x"05003304",
			3100 => x"fec130b1",
			3101 => x"0600b204",
			3102 => x"ff3030b1",
			3103 => x"006530b1",
			3104 => x"01001908",
			3105 => x"07003d04",
			3106 => x"ff8e30b1",
			3107 => x"011f30b1",
			3108 => x"ff3930b1",
			3109 => x"0c002104",
			3110 => x"fee330b1",
			3111 => x"00014904",
			3112 => x"ff7930b1",
			3113 => x"02014104",
			3114 => x"00bd30b1",
			3115 => x"ffd430b1",
			3116 => x"02012644",
			3117 => x"03003238",
			3118 => x"0a002d1c",
			3119 => x"08002614",
			3120 => x"09001c10",
			3121 => x"0b001508",
			3122 => x"0f00ae04",
			3123 => x"ffd131ad",
			3124 => x"000131ad",
			3125 => x"04001804",
			3126 => x"fff731ad",
			3127 => x"003131ad",
			3128 => x"ff8631ad",
			3129 => x"08002704",
			3130 => x"002f31ad",
			3131 => x"fff831ad",
			3132 => x"09002410",
			3133 => x"0e00910c",
			3134 => x"06007404",
			3135 => x"ffea31ad",
			3136 => x"00012a04",
			3137 => x"008831ad",
			3138 => x"ffff31ad",
			3139 => x"ffd131ad",
			3140 => x"0d002004",
			3141 => x"ff9531ad",
			3142 => x"04002904",
			3143 => x"fff931ad",
			3144 => x"003131ad",
			3145 => x"03004404",
			3146 => x"ff7131ad",
			3147 => x"05005004",
			3148 => x"001031ad",
			3149 => x"fff431ad",
			3150 => x"0600ac14",
			3151 => x"07003210",
			3152 => x"0c001504",
			3153 => x"003d31ad",
			3154 => x"0600a404",
			3155 => x"ffff31ad",
			3156 => x"05002d04",
			3157 => x"fffe31ad",
			3158 => x"ffb731ad",
			3159 => x"00a831ad",
			3160 => x"02013008",
			3161 => x"0c001804",
			3162 => x"fffe31ad",
			3163 => x"ff8931ad",
			3164 => x"0a002c04",
			3165 => x"ffaf31ad",
			3166 => x"03002e0c",
			3167 => x"0f00d304",
			3168 => x"ffeb31ad",
			3169 => x"01001704",
			3170 => x"00a931ad",
			3171 => x"fffe31ad",
			3172 => x"0a003708",
			3173 => x"0c001b04",
			3174 => x"000131ad",
			3175 => x"ff8c31ad",
			3176 => x"0600b904",
			3177 => x"005f31ad",
			3178 => x"ffe531ad",
			3179 => x"01000a04",
			3180 => x"ff083259",
			3181 => x"0201373c",
			3182 => x"0800272c",
			3183 => x"08001f10",
			3184 => x"01000e04",
			3185 => x"fee13259",
			3186 => x"0c001504",
			3187 => x"009c3259",
			3188 => x"03002404",
			3189 => x"00363259",
			3190 => x"ff5f3259",
			3191 => x"0d001b10",
			3192 => x"01001208",
			3193 => x"05003404",
			3194 => x"00983259",
			3195 => x"fed03259",
			3196 => x"09002104",
			3197 => x"ffef3259",
			3198 => x"012a3259",
			3199 => x"00012608",
			3200 => x"0f00b004",
			3201 => x"ff613259",
			3202 => x"00d03259",
			3203 => x"ff383259",
			3204 => x"0a003b08",
			3205 => x"0600bc04",
			3206 => x"fec53259",
			3207 => x"fff83259",
			3208 => x"02012c04",
			3209 => x"ff953259",
			3210 => x"00c63259",
			3211 => x"0c002214",
			3212 => x"0e00a510",
			3213 => x"08002008",
			3214 => x"0b001504",
			3215 => x"01123259",
			3216 => x"ff1a3259",
			3217 => x"03003104",
			3218 => x"01233259",
			3219 => x"005f3259",
			3220 => x"ffbe3259",
			3221 => x"ff413259",
			3222 => x"0b001f68",
			3223 => x"01001040",
			3224 => x"0b001524",
			3225 => x"04001a14",
			3226 => x"0d001410",
			3227 => x"0c001308",
			3228 => x"01000b04",
			3229 => x"ff793345",
			3230 => x"00003345",
			3231 => x"00012704",
			3232 => x"ffc63345",
			3233 => x"00973345",
			3234 => x"ff433345",
			3235 => x"0000be04",
			3236 => x"ffb23345",
			3237 => x"08001b04",
			3238 => x"ffc23345",
			3239 => x"0d001304",
			3240 => x"ffff3345",
			3241 => x"00df3345",
			3242 => x"0e009014",
			3243 => x"0d001a0c",
			3244 => x"05002608",
			3245 => x"0a002804",
			3246 => x"ffe63345",
			3247 => x"00403345",
			3248 => x"fed93345",
			3249 => x"09002304",
			3250 => x"00553345",
			3251 => x"ffa33345",
			3252 => x"0c001804",
			3253 => x"00733345",
			3254 => x"ff823345",
			3255 => x"0c00190c",
			3256 => x"08001d04",
			3257 => x"ffde3345",
			3258 => x"06007204",
			3259 => x"ffbe3345",
			3260 => x"00fd3345",
			3261 => x"09002204",
			3262 => x"ff183345",
			3263 => x"00011f0c",
			3264 => x"0200fd08",
			3265 => x"04001f04",
			3266 => x"00653345",
			3267 => x"ffcc3345",
			3268 => x"ff1b3345",
			3269 => x"07004208",
			3270 => x"05003904",
			3271 => x"00b33345",
			3272 => x"fff93345",
			3273 => x"ff613345",
			3274 => x"04002b04",
			3275 => x"fee73345",
			3276 => x"01001708",
			3277 => x"0d002004",
			3278 => x"ffe53345",
			3279 => x"00c53345",
			3280 => x"ffb33345",
			3281 => x"0f008004",
			3282 => x"fe6d33b9",
			3283 => x"08001b04",
			3284 => x"fe7633b9",
			3285 => x"07002a04",
			3286 => x"022f33b9",
			3287 => x"02012614",
			3288 => x"08002710",
			3289 => x"00012808",
			3290 => x"0f00aa04",
			3291 => x"ff1233b9",
			3292 => x"00d933b9",
			3293 => x"0d001704",
			3294 => x"00e933b9",
			3295 => x"fe6a33b9",
			3296 => x"fe6833b9",
			3297 => x"0a00310c",
			3298 => x"0f00cd04",
			3299 => x"018e33b9",
			3300 => x"0f00d304",
			3301 => x"fdfd33b9",
			3302 => x"006f33b9",
			3303 => x"04002108",
			3304 => x"08002004",
			3305 => x"ffd433b9",
			3306 => x"026733b9",
			3307 => x"08002a04",
			3308 => x"004f33b9",
			3309 => x"021533b9",
			3310 => x"0001566c",
			3311 => x"01001240",
			3312 => x"0b001310",
			3313 => x"0600b00c",
			3314 => x"0000be04",
			3315 => x"ff68349d",
			3316 => x"0d001204",
			3317 => x"ff8e349d",
			3318 => x"0172349d",
			3319 => x"ff19349d",
			3320 => x"0d001a18",
			3321 => x"0c00180c",
			3322 => x"08002008",
			3323 => x"01001004",
			3324 => x"ff22349d",
			3325 => x"00cc349d",
			3326 => x"00b8349d",
			3327 => x"0b001604",
			3328 => x"0044349d",
			3329 => x"04002004",
			3330 => x"ff1f349d",
			3331 => x"fe72349d",
			3332 => x"0500340c",
			3333 => x"08002304",
			3334 => x"ffb9349d",
			3335 => x"06002904",
			3336 => x"fff0349d",
			3337 => x"0171349d",
			3338 => x"08002204",
			3339 => x"fef5349d",
			3340 => x"01001004",
			3341 => x"ff12349d",
			3342 => x"008d349d",
			3343 => x"04001b0c",
			3344 => x"04001608",
			3345 => x"08002304",
			3346 => x"009e349d",
			3347 => x"fff2349d",
			3348 => x"fe9d349d",
			3349 => x"0b001b0c",
			3350 => x"09002104",
			3351 => x"ffd1349d",
			3352 => x"09002304",
			3353 => x"0171349d",
			3354 => x"0063349d",
			3355 => x"0f00c304",
			3356 => x"fe86349d",
			3357 => x"03002e08",
			3358 => x"04002304",
			3359 => x"015d349d",
			3360 => x"0001349d",
			3361 => x"0a003704",
			3362 => x"fe79349d",
			3363 => x"0089349d",
			3364 => x"0600ca04",
			3365 => x"0147349d",
			3366 => x"fff1349d",
			3367 => x"0001575c",
			3368 => x"0f00cd40",
			3369 => x"00013c30",
			3370 => x"05003420",
			3371 => x"0200ea10",
			3372 => x"0a002d08",
			3373 => x"0d001604",
			3374 => x"fec33561",
			3375 => x"fff13561",
			3376 => x"07002a04",
			3377 => x"01093561",
			3378 => x"ffe23561",
			3379 => x"0a002f08",
			3380 => x"01000c04",
			3381 => x"ff5e3561",
			3382 => x"01043561",
			3383 => x"0a003104",
			3384 => x"fee63561",
			3385 => x"00643561",
			3386 => x"01001204",
			3387 => x"fe983561",
			3388 => x"0c001c04",
			3389 => x"00b93561",
			3390 => x"07003d04",
			3391 => x"fee73561",
			3392 => x"009e3561",
			3393 => x"0100160c",
			3394 => x"04002508",
			3395 => x"01000c04",
			3396 => x"ff963561",
			3397 => x"00e33561",
			3398 => x"ffaf3561",
			3399 => x"015b3561",
			3400 => x"0f00cf04",
			3401 => x"fec43561",
			3402 => x"0e00a314",
			3403 => x"0c002210",
			3404 => x"05003308",
			3405 => x"00014604",
			3406 => x"feea3561",
			3407 => x"002a3561",
			3408 => x"05003804",
			3409 => x"00ec3561",
			3410 => x"ff933561",
			3411 => x"feed3561",
			3412 => x"fed83561",
			3413 => x"0600ca04",
			3414 => x"011c3561",
			3415 => x"001b3561",
			3416 => x"0201494c",
			3417 => x"03004644",
			3418 => x"05003a3c",
			3419 => x"08002020",
			3420 => x"0b001310",
			3421 => x"09001908",
			3422 => x"04002004",
			3423 => x"ff6935ff",
			3424 => x"000e35ff",
			3425 => x"04001a04",
			3426 => x"fff035ff",
			3427 => x"00bb35ff",
			3428 => x"0600b608",
			3429 => x"04002604",
			3430 => x"ff2b35ff",
			3431 => x"002435ff",
			3432 => x"0600bb04",
			3433 => x"006035ff",
			3434 => x"ff9035ff",
			3435 => x"0b00180c",
			3436 => x"0000c704",
			3437 => x"ffb935ff",
			3438 => x"00012504",
			3439 => x"003735ff",
			3440 => x"00bb35ff",
			3441 => x"09002508",
			3442 => x"07003604",
			3443 => x"fff435ff",
			3444 => x"ff0635ff",
			3445 => x"0b001c04",
			3446 => x"00dc35ff",
			3447 => x"ffd335ff",
			3448 => x"04002704",
			3449 => x"ffc335ff",
			3450 => x"fef035ff",
			3451 => x"0f009804",
			3452 => x"fff135ff",
			3453 => x"00b835ff",
			3454 => x"00ac35ff",
			3455 => x"0a003b24",
			3456 => x"0a003820",
			3457 => x"0300341c",
			3458 => x"0a003714",
			3459 => x"01001a0c",
			3460 => x"01001908",
			3461 => x"02013f04",
			3462 => x"ffef3669",
			3463 => x"00b53669",
			3464 => x"fe813669",
			3465 => x"01001d04",
			3466 => x"01a93669",
			3467 => x"fee73669",
			3468 => x"01001204",
			3469 => x"ff343669",
			3470 => x"01693669",
			3471 => x"fe8c3669",
			3472 => x"fe623669",
			3473 => x"00012804",
			3474 => x"feac3669",
			3475 => x"0600b70c",
			3476 => x"00013a08",
			3477 => x"0600a904",
			3478 => x"01793669",
			3479 => x"fec53669",
			3480 => x"01c63669",
			3481 => x"fecf3669",
			3482 => x"0200b704",
			3483 => x"feb036d5",
			3484 => x"07002a10",
			3485 => x"0d001308",
			3486 => x"07002404",
			3487 => x"005b36d5",
			3488 => x"ff3836d5",
			3489 => x"06007204",
			3490 => x"ff6d36d5",
			3491 => x"015436d5",
			3492 => x"0f00a904",
			3493 => x"fea636d5",
			3494 => x"0f00b308",
			3495 => x"0b001a04",
			3496 => x"012436d5",
			3497 => x"ff0136d5",
			3498 => x"00012208",
			3499 => x"07003004",
			3500 => x"001436d5",
			3501 => x"fe7b36d5",
			3502 => x"08002008",
			3503 => x"0b001504",
			3504 => x"005736d5",
			3505 => x"fece36d5",
			3506 => x"0b001804",
			3507 => x"013336d5",
			3508 => x"001236d5",
			3509 => x"0100102c",
			3510 => x"0b00151c",
			3511 => x"02013014",
			3512 => x"0400230c",
			3513 => x"0a002708",
			3514 => x"01000c04",
			3515 => x"ffda37a9",
			3516 => x"003937a9",
			3517 => x"ff7837a9",
			3518 => x"0a003104",
			3519 => x"005a37a9",
			3520 => x"ffe337a9",
			3521 => x"01000a04",
			3522 => x"ffb637a9",
			3523 => x"00aa37a9",
			3524 => x"0c001608",
			3525 => x"03002f04",
			3526 => x"002a37a9",
			3527 => x"ffec37a9",
			3528 => x"08002404",
			3529 => x"ff2437a9",
			3530 => x"001937a9",
			3531 => x"07003718",
			3532 => x"0b001b0c",
			3533 => x"0f00aa08",
			3534 => x"04001d04",
			3535 => x"001f37a9",
			3536 => x"ff8b37a9",
			3537 => x"00ad37a9",
			3538 => x"09002504",
			3539 => x"ff8737a9",
			3540 => x"05003504",
			3541 => x"002a37a9",
			3542 => x"fff837a9",
			3543 => x"0100160c",
			3544 => x"0a004308",
			3545 => x"0600b704",
			3546 => x"ff1c37a9",
			3547 => x"fffe37a9",
			3548 => x"006837a9",
			3549 => x"03002e0c",
			3550 => x"0d002108",
			3551 => x"00013604",
			3552 => x"001f37a9",
			3553 => x"00c437a9",
			3554 => x"ffa337a9",
			3555 => x"04002904",
			3556 => x"ff3637a9",
			3557 => x"05003a04",
			3558 => x"006837a9",
			3559 => x"03004604",
			3560 => x"ff8c37a9",
			3561 => x"004337a9",
			3562 => x"0f008c0c",
			3563 => x"0c001608",
			3564 => x"08001f04",
			3565 => x"fe6e3815",
			3566 => x"01cb3815",
			3567 => x"fe613815",
			3568 => x"01000a04",
			3569 => x"fe643815",
			3570 => x"0d002124",
			3571 => x"0a00431c",
			3572 => x"0b001610",
			3573 => x"05002408",
			3574 => x"0c001404",
			3575 => x"fe373815",
			3576 => x"002f3815",
			3577 => x"08001b04",
			3578 => x"fe963815",
			3579 => x"01e63815",
			3580 => x"01000e04",
			3581 => x"fe143815",
			3582 => x"03002e04",
			3583 => x"012f3815",
			3584 => x"000b3815",
			3585 => x"00010c04",
			3586 => x"fec63815",
			3587 => x"02bf3815",
			3588 => x"fe643815",
			3589 => x"0100102c",
			3590 => x"0b00151c",
			3591 => x"02013014",
			3592 => x"0400230c",
			3593 => x"0a002708",
			3594 => x"00011404",
			3595 => x"ffdd38e9",
			3596 => x"003738e9",
			3597 => x"ff7038e9",
			3598 => x"0a003104",
			3599 => x"005f38e9",
			3600 => x"ffe138e9",
			3601 => x"01000a04",
			3602 => x"ffb438e9",
			3603 => x"00b038e9",
			3604 => x"0c001608",
			3605 => x"03002f04",
			3606 => x"002b38e9",
			3607 => x"ffeb38e9",
			3608 => x"08002404",
			3609 => x"ff1638e9",
			3610 => x"001a38e9",
			3611 => x"07003714",
			3612 => x"0f00aa0c",
			3613 => x"03002108",
			3614 => x"07002604",
			3615 => x"ffea38e9",
			3616 => x"004038e9",
			3617 => x"ff7e38e9",
			3618 => x"01001204",
			3619 => x"001a38e9",
			3620 => x"00ce38e9",
			3621 => x"04002108",
			3622 => x"0d001f04",
			3623 => x"008638e9",
			3624 => x"ffab38e9",
			3625 => x"0400290c",
			3626 => x"08002d08",
			3627 => x"03002a04",
			3628 => x"ffe138e9",
			3629 => x"ff1638e9",
			3630 => x"004838e9",
			3631 => x"0d00200c",
			3632 => x"03003b08",
			3633 => x"01001804",
			3634 => x"ff6038e9",
			3635 => x"fffa38e9",
			3636 => x"005838e9",
			3637 => x"01001708",
			3638 => x"01001404",
			3639 => x"fff738e9",
			3640 => x"00c738e9",
			3641 => x"ffba38e9",
			3642 => x"01000c20",
			3643 => x"0f008108",
			3644 => x"06007304",
			3645 => x"ffda39ad",
			3646 => x"004f39ad",
			3647 => x"0e009e14",
			3648 => x"0300230c",
			3649 => x"07002c08",
			3650 => x"03001f04",
			3651 => x"fff639ad",
			3652 => x"002e39ad",
			3653 => x"ffef39ad",
			3654 => x"07003704",
			3655 => x"ff0d39ad",
			3656 => x"fff939ad",
			3657 => x"002239ad",
			3658 => x"07003f30",
			3659 => x"0a003b1c",
			3660 => x"05003914",
			3661 => x"0d002110",
			3662 => x"02013708",
			3663 => x"0f00ca04",
			3664 => x"004339ad",
			3665 => x"ff8a39ad",
			3666 => x"0600b504",
			3667 => x"ffcb39ad",
			3668 => x"00e439ad",
			3669 => x"ff7139ad",
			3670 => x"07003004",
			3671 => x"001539ad",
			3672 => x"ff3339ad",
			3673 => x"09002608",
			3674 => x"01001204",
			3675 => x"ffe839ad",
			3676 => x"00d439ad",
			3677 => x"0c002208",
			3678 => x"05005d04",
			3679 => x"ff7139ad",
			3680 => x"001639ad",
			3681 => x"009239ad",
			3682 => x"0c002108",
			3683 => x"0f00d004",
			3684 => x"000b39ad",
			3685 => x"ff3839ad",
			3686 => x"00014904",
			3687 => x"ffb339ad",
			3688 => x"02014204",
			3689 => x"006039ad",
			3690 => x"ffd339ad",
			3691 => x"0f00ae14",
			3692 => x"0f008004",
			3693 => x"fe5b3a51",
			3694 => x"0e006804",
			3695 => x"01ed3a51",
			3696 => x"06007f08",
			3697 => x"0c001a04",
			3698 => x"014b3a51",
			3699 => x"fe6e3a51",
			3700 => x"fe563a51",
			3701 => x"0d001f34",
			3702 => x"01000c10",
			3703 => x"08001c04",
			3704 => x"fe5e3a51",
			3705 => x"0b001508",
			3706 => x"0f00c704",
			3707 => x"fe873a51",
			3708 => x"035b3a51",
			3709 => x"fe3a3a51",
			3710 => x"00014618",
			3711 => x"08002610",
			3712 => x"08001f08",
			3713 => x"0c001504",
			3714 => x"03583a51",
			3715 => x"fee93a51",
			3716 => x"0f00ba04",
			3717 => x"05ca3a51",
			3718 => x"02ec3a51",
			3719 => x"05003604",
			3720 => x"00dc3a51",
			3721 => x"fe5f3a51",
			3722 => x"05003908",
			3723 => x"08002004",
			3724 => x"036e3a51",
			3725 => x"04933a51",
			3726 => x"01033a51",
			3727 => x"01001708",
			3728 => x"0d002004",
			3729 => x"fe5d3a51",
			3730 => x"02863a51",
			3731 => x"fe523a51",
			3732 => x"08002034",
			3733 => x"0b00130c",
			3734 => x"05002404",
			3735 => x"fed93b2d",
			3736 => x"08001b04",
			3737 => x"ff763b2d",
			3738 => x"015b3b2d",
			3739 => x"05002e18",
			3740 => x"01001010",
			3741 => x"0f00d80c",
			3742 => x"04002004",
			3743 => x"fe8a3b2d",
			3744 => x"07002d04",
			3745 => x"feec3b2d",
			3746 => x"007f3b2d",
			3747 => x"00a83b2d",
			3748 => x"0c001904",
			3749 => x"011c3b2d",
			3750 => x"ff123b2d",
			3751 => x"05003808",
			3752 => x"09001b04",
			3753 => x"ffdc3b2d",
			3754 => x"fe743b2d",
			3755 => x"05003a04",
			3756 => x"00bb3b2d",
			3757 => x"fed63b2d",
			3758 => x"0b001910",
			3759 => x"0500350c",
			3760 => x"04002208",
			3761 => x"05002a04",
			3762 => x"010b3b2d",
			3763 => x"00103b2d",
			3764 => x"01903b2d",
			3765 => x"00033b2d",
			3766 => x"01001210",
			3767 => x"0a003408",
			3768 => x"07003404",
			3769 => x"fefc3b2d",
			3770 => x"00cf3b2d",
			3771 => x"08002604",
			3772 => x"fe6f3b2d",
			3773 => x"00833b2d",
			3774 => x"04001d0c",
			3775 => x"01001408",
			3776 => x"04001504",
			3777 => x"fff63b2d",
			3778 => x"00673b2d",
			3779 => x"fe7a3b2d",
			3780 => x"0d001b04",
			3781 => x"010c3b2d",
			3782 => x"03002904",
			3783 => x"01103b2d",
			3784 => x"05003304",
			3785 => x"fe9f3b2d",
			3786 => x"002a3b2d",
			3787 => x"0f008c0c",
			3788 => x"0c001608",
			3789 => x"0d001504",
			3790 => x"fe643ba1",
			3791 => x"03bb3ba1",
			3792 => x"fe603ba1",
			3793 => x"01000a04",
			3794 => x"fe673ba1",
			3795 => x"0d002228",
			3796 => x"00014618",
			3797 => x"08001f08",
			3798 => x"0b001304",
			3799 => x"01c63ba1",
			3800 => x"fe543ba1",
			3801 => x"0b001908",
			3802 => x"09001d04",
			3803 => x"00513ba1",
			3804 => x"02273ba1",
			3805 => x"01001204",
			3806 => x"fe123ba1",
			3807 => x"00b33ba1",
			3808 => x"0e00a50c",
			3809 => x"08002004",
			3810 => x"00f53ba1",
			3811 => x"05003404",
			3812 => x"02143ba1",
			3813 => x"02d93ba1",
			3814 => x"ffee3ba1",
			3815 => x"fe533ba1",
			3816 => x"0f008c0c",
			3817 => x"0b001308",
			3818 => x"00009504",
			3819 => x"fe9a3c0d",
			3820 => x"03093c0d",
			3821 => x"fe623c0d",
			3822 => x"01000a04",
			3823 => x"fe673c0d",
			3824 => x"07002a04",
			3825 => x"02523c0d",
			3826 => x"07004420",
			3827 => x"01001010",
			3828 => x"0b001508",
			3829 => x"05002704",
			3830 => x"ff9e3c0d",
			3831 => x"01e23c0d",
			3832 => x"01000e04",
			3833 => x"fe303c0d",
			3834 => x"00133c0d",
			3835 => x"0c001908",
			3836 => x"04002004",
			3837 => x"00c33c0d",
			3838 => x"022d3c0d",
			3839 => x"00011f04",
			3840 => x"feea3c0d",
			3841 => x"00cc3c0d",
			3842 => x"fe6f3c0d",
			3843 => x"0a003b48",
			3844 => x"00014630",
			3845 => x"0f00ca20",
			3846 => x"0a00381c",
			3847 => x"04002610",
			3848 => x"04002108",
			3849 => x"02012704",
			3850 => x"ffc73cb9",
			3851 => x"00c63cb9",
			3852 => x"0f00b704",
			3853 => x"ffe23cb9",
			3854 => x"ff093cb9",
			3855 => x"08002608",
			3856 => x"03003404",
			3857 => x"01163cb9",
			3858 => x"ff913cb9",
			3859 => x"ff543cb9",
			3860 => x"ff243cb9",
			3861 => x"0a00370c",
			3862 => x"04001e08",
			3863 => x"0a003104",
			3864 => x"ff643cb9",
			3865 => x"005a3cb9",
			3866 => x"ff103cb9",
			3867 => x"00243cb9",
			3868 => x"0d001f10",
			3869 => x"0800200c",
			3870 => x"0b001508",
			3871 => x"0d001304",
			3872 => x"ffeb3cb9",
			3873 => x"00ac3cb9",
			3874 => x"ff7d3cb9",
			3875 => x"00e73cb9",
			3876 => x"04002704",
			3877 => x"ff633cb9",
			3878 => x"001e3cb9",
			3879 => x"0600b70c",
			3880 => x"00012a04",
			3881 => x"ffa43cb9",
			3882 => x"01001704",
			3883 => x"01013cb9",
			3884 => x"ffec3cb9",
			3885 => x"ffa23cb9",
			3886 => x"0a003b3c",
			3887 => x"05003a38",
			3888 => x"08002624",
			3889 => x"04002614",
			3890 => x"04002410",
			3891 => x"00013008",
			3892 => x"0f00b104",
			3893 => x"00563d5d",
			3894 => x"fee03d5d",
			3895 => x"08002204",
			3896 => x"ffe33d5d",
			3897 => x"00ce3d5d",
			3898 => x"fec33d5d",
			3899 => x"0300310c",
			3900 => x"02011808",
			3901 => x"01000c04",
			3902 => x"008d3d5d",
			3903 => x"ff313d5d",
			3904 => x"012f3d5d",
			3905 => x"ffec3d5d",
			3906 => x"0201370c",
			3907 => x"07003304",
			3908 => x"009e3d5d",
			3909 => x"0600bc04",
			3910 => x"fe8c3d5d",
			3911 => x"00043d5d",
			3912 => x"03002e04",
			3913 => x"00ed3d5d",
			3914 => x"ff243d5d",
			3915 => x"fecb3d5d",
			3916 => x"05003f08",
			3917 => x"0e008b04",
			3918 => x"ffd33d5d",
			3919 => x"01363d5d",
			3920 => x"0a004304",
			3921 => x"ff023d5d",
			3922 => x"0b001f08",
			3923 => x"08002004",
			3924 => x"ffd63d5d",
			3925 => x"00f23d5d",
			3926 => x"ffa83d5d",
			3927 => x"08002754",
			3928 => x"08001f20",
			3929 => x"02013414",
			3930 => x"0f008108",
			3931 => x"06007204",
			3932 => x"ffee3e31",
			3933 => x"001b3e31",
			3934 => x"0a002a08",
			3935 => x"0a002504",
			3936 => x"ffe73e31",
			3937 => x"00113e31",
			3938 => x"ff673e31",
			3939 => x"0e009a08",
			3940 => x"01000a04",
			3941 => x"fff33e31",
			3942 => x"00673e31",
			3943 => x"ffc43e31",
			3944 => x"0c00180c",
			3945 => x"05002504",
			3946 => x"ffdb3e31",
			3947 => x"0f008004",
			3948 => x"ffe73e31",
			3949 => x"00a03e31",
			3950 => x"08002318",
			3951 => x"04002610",
			3952 => x"0d001b08",
			3953 => x"0600a204",
			3954 => x"00053e31",
			3955 => x"ff6d3e31",
			3956 => x"0d001d04",
			3957 => x"00123e31",
			3958 => x"fff53e31",
			3959 => x"00011d04",
			3960 => x"ffe53e31",
			3961 => x"00503e31",
			3962 => x"0f00af04",
			3963 => x"ffc93e31",
			3964 => x"0c001f08",
			3965 => x"01001404",
			3966 => x"007a3e31",
			3967 => x"00173e31",
			3968 => x"ffdf3e31",
			3969 => x"04002108",
			3970 => x"08002a04",
			3971 => x"002a3e31",
			3972 => x"ffd33e31",
			3973 => x"08002d08",
			3974 => x"03005304",
			3975 => x"ff553e31",
			3976 => x"00093e31",
			3977 => x"0e009504",
			3978 => x"00273e31",
			3979 => x"ffe53e31",
			3980 => x"0f008c0c",
			3981 => x"0c001608",
			3982 => x"01001004",
			3983 => x"fe733ebd",
			3984 => x"01f53ebd",
			3985 => x"fe663ebd",
			3986 => x"01000a04",
			3987 => x"fe6e3ebd",
			3988 => x"0c001818",
			3989 => x"05002408",
			3990 => x"03002404",
			3991 => x"006a3ebd",
			3992 => x"fe523ebd",
			3993 => x"09001f0c",
			3994 => x"07002b04",
			3995 => x"021c3ebd",
			3996 => x"0b001604",
			3997 => x"00fc3ebd",
			3998 => x"fee43ebd",
			3999 => x"021d3ebd",
			4000 => x"0100120c",
			4001 => x"0d001a08",
			4002 => x"0b001804",
			4003 => x"ffeb3ebd",
			4004 => x"fe1b3ebd",
			4005 => x"014c3ebd",
			4006 => x"03002704",
			4007 => x"feaa3ebd",
			4008 => x"03002e08",
			4009 => x"02012b04",
			4010 => x"00243ebd",
			4011 => x"02773ebd",
			4012 => x"0b001b04",
			4013 => x"01483ebd",
			4014 => x"ff953ebd",
			4015 => x"0f008004",
			4016 => x"fe733f41",
			4017 => x"08001c0c",
			4018 => x"0a002708",
			4019 => x"09001a04",
			4020 => x"fed33f41",
			4021 => x"01c13f41",
			4022 => x"fe703f41",
			4023 => x"0c001714",
			4024 => x"05002404",
			4025 => x"ff343f41",
			4026 => x"07003008",
			4027 => x"0c001604",
			4028 => x"01ff3f41",
			4029 => x"01313f41",
			4030 => x"00012b04",
			4031 => x"fe903f41",
			4032 => x"012d3f41",
			4033 => x"04001e08",
			4034 => x"0f00c604",
			4035 => x"fdfb3f41",
			4036 => x"ffc23f41",
			4037 => x"08001f08",
			4038 => x"09002004",
			4039 => x"fe6f3f41",
			4040 => x"00363f41",
			4041 => x"0c001908",
			4042 => x"04002304",
			4043 => x"00d23f41",
			4044 => x"019e3f41",
			4045 => x"09002104",
			4046 => x"fe333f41",
			4047 => x"00873f41",
			4048 => x"06009514",
			4049 => x"01000b10",
			4050 => x"0b00150c",
			4051 => x"04002304",
			4052 => x"ffdf3fed",
			4053 => x"01000704",
			4054 => x"fffa3fed",
			4055 => x"00ab3fed",
			4056 => x"ffa83fed",
			4057 => x"fef13fed",
			4058 => x"0f00b30c",
			4059 => x"0b001a08",
			4060 => x"0000f304",
			4061 => x"ffc93fed",
			4062 => x"00fc3fed",
			4063 => x"ff963fed",
			4064 => x"0001220c",
			4065 => x"04001a08",
			4066 => x"07003104",
			4067 => x"00303fed",
			4068 => x"ffda3fed",
			4069 => x"fefa3fed",
			4070 => x"07004020",
			4071 => x"0600a710",
			4072 => x"04002608",
			4073 => x"02012f04",
			4074 => x"fedd3fed",
			4075 => x"00583fed",
			4076 => x"00012c04",
			4077 => x"00f33fed",
			4078 => x"ff6e3fed",
			4079 => x"0600a908",
			4080 => x"0e008904",
			4081 => x"ffda3fed",
			4082 => x"010d3fed",
			4083 => x"0b001a04",
			4084 => x"005f3fed",
			4085 => x"ffce3fed",
			4086 => x"0c002104",
			4087 => x"ff2c3fed",
			4088 => x"0d002104",
			4089 => x"004b3fed",
			4090 => x"ff933fed",
			4091 => x"00013c44",
			4092 => x"08001f14",
			4093 => x"0b001310",
			4094 => x"0c001304",
			4095 => x"ffd940a9",
			4096 => x"0b001204",
			4097 => x"fff740a9",
			4098 => x"01000704",
			4099 => x"fffb40a9",
			4100 => x"005140a9",
			4101 => x"ff6140a9",
			4102 => x"0c001c18",
			4103 => x"0b001b14",
			4104 => x"0000d308",
			4105 => x"03002104",
			4106 => x"002440a9",
			4107 => x"ffaf40a9",
			4108 => x"05003708",
			4109 => x"05002c04",
			4110 => x"fff740a9",
			4111 => x"009240a9",
			4112 => x"fff340a9",
			4113 => x"ffb740a9",
			4114 => x"00012608",
			4115 => x"0f00bc04",
			4116 => x"ffa340a9",
			4117 => x"007940a9",
			4118 => x"03003d0c",
			4119 => x"08002704",
			4120 => x"ff4340a9",
			4121 => x"0600a904",
			4122 => x"002940a9",
			4123 => x"ffc040a9",
			4124 => x"003840a9",
			4125 => x"09002b18",
			4126 => x"01000a04",
			4127 => x"ffc340a9",
			4128 => x"0e00a510",
			4129 => x"08002008",
			4130 => x"0b001504",
			4131 => x"009540a9",
			4132 => x"ff8540a9",
			4133 => x"01001904",
			4134 => x"008e40a9",
			4135 => x"000340a9",
			4136 => x"ffe340a9",
			4137 => x"ffa640a9",
			4138 => x"02012650",
			4139 => x"0c001c3c",
			4140 => x"0600951c",
			4141 => x"01000b10",
			4142 => x"0b00150c",
			4143 => x"03002404",
			4144 => x"fff541b5",
			4145 => x"0000d704",
			4146 => x"004341b5",
			4147 => x"fffb41b5",
			4148 => x"ffda41b5",
			4149 => x"03002108",
			4150 => x"03001d04",
			4151 => x"fff041b5",
			4152 => x"002841b5",
			4153 => x"ff5941b5",
			4154 => x"06009d0c",
			4155 => x"0f00b308",
			4156 => x"01000a04",
			4157 => x"fffb41b5",
			4158 => x"00ad41b5",
			4159 => x"ffe241b5",
			4160 => x"00012708",
			4161 => x"04001a04",
			4162 => x"fff641b5",
			4163 => x"ff6241b5",
			4164 => x"0600a204",
			4165 => x"ffc041b5",
			4166 => x"0f00c804",
			4167 => x"008141b5",
			4168 => x"ffed41b5",
			4169 => x"01001a0c",
			4170 => x"0a005404",
			4171 => x"ff5341b5",
			4172 => x"05007604",
			4173 => x"000b41b5",
			4174 => x"fffb41b5",
			4175 => x"0e009104",
			4176 => x"fff141b5",
			4177 => x"004441b5",
			4178 => x"0600ad14",
			4179 => x"0600a708",
			4180 => x"00013c04",
			4181 => x"ff9e41b5",
			4182 => x"003841b5",
			4183 => x"0f00c908",
			4184 => x"01000e04",
			4185 => x"001341b5",
			4186 => x"00e441b5",
			4187 => x"fff141b5",
			4188 => x"00014810",
			4189 => x"0d001c08",
			4190 => x"03002f04",
			4191 => x"ff3441b5",
			4192 => x"002541b5",
			4193 => x"05003804",
			4194 => x"004d41b5",
			4195 => x"ff9941b5",
			4196 => x"0100180c",
			4197 => x"02014408",
			4198 => x"08002204",
			4199 => x"ffcf41b5",
			4200 => x"004f41b5",
			4201 => x"00a741b5",
			4202 => x"01001a04",
			4203 => x"ffa041b5",
			4204 => x"001c41b5",
			4205 => x"0001333c",
			4206 => x"01001330",
			4207 => x"04002624",
			4208 => x"07003114",
			4209 => x"0200ea0c",
			4210 => x"0f008108",
			4211 => x"01001104",
			4212 => x"00214279",
			4213 => x"ffed4279",
			4214 => x"ffaf4279",
			4215 => x"01000c04",
			4216 => x"ffe54279",
			4217 => x"005f4279",
			4218 => x"0700360c",
			4219 => x"00010608",
			4220 => x"06009d04",
			4221 => x"00184279",
			4222 => x"ffea4279",
			4223 => x"ff714279",
			4224 => x"00194279",
			4225 => x"00011608",
			4226 => x"0a002f04",
			4227 => x"00134279",
			4228 => x"ffce4279",
			4229 => x"006d4279",
			4230 => x"0200fd08",
			4231 => x"0b001c04",
			4232 => x"00244279",
			4233 => x"fff34279",
			4234 => x"ff614279",
			4235 => x"05003920",
			4236 => x"09002b1c",
			4237 => x"0600a808",
			4238 => x"00013c04",
			4239 => x"ffbb4279",
			4240 => x"00194279",
			4241 => x"01000a04",
			4242 => x"ffd04279",
			4243 => x"05003508",
			4244 => x"00014604",
			4245 => x"002e4279",
			4246 => x"00954279",
			4247 => x"0d001d04",
			4248 => x"00214279",
			4249 => x"ffea4279",
			4250 => x"ffbe4279",
			4251 => x"03003a04",
			4252 => x"ff844279",
			4253 => x"003f4279",
			4254 => x"08001c04",
			4255 => x"fe984315",
			4256 => x"00014734",
			4257 => x"0a003b24",
			4258 => x"00012a14",
			4259 => x"01001a10",
			4260 => x"0e008808",
			4261 => x"0c001c04",
			4262 => x"00b34315",
			4263 => x"feba4315",
			4264 => x"02011904",
			4265 => x"fe754315",
			4266 => x"00384315",
			4267 => x"01934315",
			4268 => x"0f00c004",
			4269 => x"fe804315",
			4270 => x"0600ad04",
			4271 => x"00904315",
			4272 => x"0d001c04",
			4273 => x"fedb4315",
			4274 => x"00454315",
			4275 => x"00012804",
			4276 => x"fee64315",
			4277 => x"00013d08",
			4278 => x"0600a904",
			4279 => x"01384315",
			4280 => x"fed74315",
			4281 => x"01974315",
			4282 => x"0a00360c",
			4283 => x"01001808",
			4284 => x"01000e04",
			4285 => x"00724315",
			4286 => x"01624315",
			4287 => x"00164315",
			4288 => x"03003304",
			4289 => x"fedb4315",
			4290 => x"04002c04",
			4291 => x"01214315",
			4292 => x"ff574315",
			4293 => x"0a002c08",
			4294 => x"02013904",
			4295 => x"ff9743c1",
			4296 => x"001143c1",
			4297 => x"05002e1c",
			4298 => x"08001d10",
			4299 => x"05002708",
			4300 => x"0e009404",
			4301 => x"000243c1",
			4302 => x"ffd043c1",
			4303 => x"00014204",
			4304 => x"ffef43c1",
			4305 => x"002043c1",
			4306 => x"03002e08",
			4307 => x"0000d604",
			4308 => x"fffb43c1",
			4309 => x"007f43c1",
			4310 => x"fff243c1",
			4311 => x"0100172c",
			4312 => x"0d001a14",
			4313 => x"01001210",
			4314 => x"0c001608",
			4315 => x"01000a04",
			4316 => x"fff643c1",
			4317 => x"002b43c1",
			4318 => x"0e008e04",
			4319 => x"ff5d43c1",
			4320 => x"fffa43c1",
			4321 => x"002543c1",
			4322 => x"0b001b08",
			4323 => x"04002504",
			4324 => x"007f43c1",
			4325 => x"001043c1",
			4326 => x"0c001e08",
			4327 => x"0e008e04",
			4328 => x"000643c1",
			4329 => x"ff9243c1",
			4330 => x"05003804",
			4331 => x"007e43c1",
			4332 => x"ffe543c1",
			4333 => x"0d001f04",
			4334 => x"001a43c1",
			4335 => x"ff8343c1",
			4336 => x"09002544",
			4337 => x"0b001b38",
			4338 => x"02014330",
			4339 => x"0f00cb1c",
			4340 => x"0600a810",
			4341 => x"0600a308",
			4342 => x"01000e04",
			4343 => x"ff63449d",
			4344 => x"0074449d",
			4345 => x"02012d04",
			4346 => x"fea0449d",
			4347 => x"ffd4449d",
			4348 => x"00012704",
			4349 => x"fec9449d",
			4350 => x"0a003604",
			4351 => x"0181449d",
			4352 => x"0034449d",
			4353 => x"0001470c",
			4354 => x"0e009804",
			4355 => x"fe86449d",
			4356 => x"0f00d904",
			4357 => x"0009449d",
			4358 => x"fefe449d",
			4359 => x"03002d04",
			4360 => x"ff73449d",
			4361 => x"0098449d",
			4362 => x"0600c804",
			4363 => x"013e449d",
			4364 => x"0055449d",
			4365 => x"05002e08",
			4366 => x"05001e04",
			4367 => x"ffef449d",
			4368 => x"00cd449d",
			4369 => x"fe89449d",
			4370 => x"0500381c",
			4371 => x"07004418",
			4372 => x"0300270c",
			4373 => x"0d001b08",
			4374 => x"08002204",
			4375 => x"fffb449d",
			4376 => x"0012449d",
			4377 => x"fee2449d",
			4378 => x"0e008604",
			4379 => x"ff09449d",
			4380 => x"05003304",
			4381 => x"004e449d",
			4382 => x"014c449d",
			4383 => x"fedc449d",
			4384 => x"03004608",
			4385 => x"00014f04",
			4386 => x"fe97449d",
			4387 => x"008d449d",
			4388 => x"00010704",
			4389 => x"ffb5449d",
			4390 => x"012d449d",
			4391 => x"01001034",
			4392 => x"0b00172c",
			4393 => x"0e008d20",
			4394 => x"0b00140c",
			4395 => x"0d001304",
			4396 => x"ffc84591",
			4397 => x"0000be04",
			4398 => x"ffe94591",
			4399 => x"00a24591",
			4400 => x"0c001404",
			4401 => x"00264591",
			4402 => x"04002608",
			4403 => x"05002604",
			4404 => x"ffeb4591",
			4405 => x"ff244591",
			4406 => x"09001f04",
			4407 => x"ffeb4591",
			4408 => x"00304591",
			4409 => x"08001c04",
			4410 => x"ffa04591",
			4411 => x"00012704",
			4412 => x"ffa94591",
			4413 => x"00b34591",
			4414 => x"08002404",
			4415 => x"ff194591",
			4416 => x"00204591",
			4417 => x"0b001b18",
			4418 => x"0c001c14",
			4419 => x"03002d0c",
			4420 => x"0f00bc08",
			4421 => x"05002704",
			4422 => x"ffc54591",
			4423 => x"00944591",
			4424 => x"ffd14591",
			4425 => x"0b001904",
			4426 => x"004a4591",
			4427 => x"00e44591",
			4428 => x"ffbe4591",
			4429 => x"0e009114",
			4430 => x"03002a08",
			4431 => x"01001604",
			4432 => x"ffd74591",
			4433 => x"00794591",
			4434 => x"01001308",
			4435 => x"01001204",
			4436 => x"ffb74591",
			4437 => x"00254591",
			4438 => x"ff0c4591",
			4439 => x"0e009508",
			4440 => x"0a003804",
			4441 => x"00d64591",
			4442 => x"ffe14591",
			4443 => x"01001708",
			4444 => x"05003804",
			4445 => x"00804591",
			4446 => x"ffac4591",
			4447 => x"01001a04",
			4448 => x"ff2d4591",
			4449 => x"0f00d904",
			4450 => x"ffce4591",
			4451 => x"002f4591",
			4452 => x"0e009c50",
			4453 => x"04002628",
			4454 => x"04002424",
			4455 => x"0d001f20",
			4456 => x"01000c10",
			4457 => x"0f008108",
			4458 => x"03002904",
			4459 => x"ffed4655",
			4460 => x"00414655",
			4461 => x"0e009304",
			4462 => x"ff5a4655",
			4463 => x"001c4655",
			4464 => x"0e008e08",
			4465 => x"06009e04",
			4466 => x"008a4655",
			4467 => x"ffb54655",
			4468 => x"0e009404",
			4469 => x"00ba4655",
			4470 => x"ffff4655",
			4471 => x"ff694655",
			4472 => x"ff4c4655",
			4473 => x"08002618",
			4474 => x"0c001f14",
			4475 => x"00011608",
			4476 => x"05003504",
			4477 => x"002e4655",
			4478 => x"ffa54655",
			4479 => x"09002108",
			4480 => x"03003304",
			4481 => x"00794655",
			4482 => x"ff9d4655",
			4483 => x"010c4655",
			4484 => x"ffb44655",
			4485 => x"0d002004",
			4486 => x"ff4a4655",
			4487 => x"08002a04",
			4488 => x"ffdc4655",
			4489 => x"00013404",
			4490 => x"fff44655",
			4491 => x"00be4655",
			4492 => x"01001a0c",
			4493 => x"0f00d404",
			4494 => x"00104655",
			4495 => x"02014704",
			4496 => x"ff534655",
			4497 => x"ffdd4655",
			4498 => x"03002e04",
			4499 => x"00394655",
			4500 => x"ffe64655",
			4501 => x"08002030",
			4502 => x"02013f2c",
			4503 => x"06009e20",
			4504 => x"0e006f0c",
			4505 => x"0b001308",
			4506 => x"0b001204",
			4507 => x"ffef4749",
			4508 => x"001f4749",
			4509 => x"ffa84749",
			4510 => x"06009a0c",
			4511 => x"0a002a04",
			4512 => x"00504749",
			4513 => x"0b001704",
			4514 => x"fff44749",
			4515 => x"00044749",
			4516 => x"0f00b704",
			4517 => x"ffdb4749",
			4518 => x"00154749",
			4519 => x"04002608",
			4520 => x"07002a04",
			4521 => x"00064749",
			4522 => x"ff334749",
			4523 => x"000c4749",
			4524 => x"00174749",
			4525 => x"0b001b1c",
			4526 => x"02011c10",
			4527 => x"0600a00c",
			4528 => x"04002508",
			4529 => x"05002c04",
			4530 => x"fff74749",
			4531 => x"00764749",
			4532 => x"ffb74749",
			4533 => x"ff734749",
			4534 => x"05003908",
			4535 => x"0d001904",
			4536 => x"000f4749",
			4537 => x"00ae4749",
			4538 => x"00024749",
			4539 => x"0e009110",
			4540 => x"03002a08",
			4541 => x"08002704",
			4542 => x"ffe84749",
			4543 => x"00334749",
			4544 => x"0a005b04",
			4545 => x"ff484749",
			4546 => x"000a4749",
			4547 => x"0e009508",
			4548 => x"0a003804",
			4549 => x"00874749",
			4550 => x"fff94749",
			4551 => x"0100170c",
			4552 => x"0c001e04",
			4553 => x"ffbc4749",
			4554 => x"01001604",
			4555 => x"ffe74749",
			4556 => x"00744749",
			4557 => x"01001a04",
			4558 => x"ff704749",
			4559 => x"09002b04",
			4560 => x"00244749",
			4561 => x"ffe04749",
			4562 => x"08001c04",
			4563 => x"fe7447e5",
			4564 => x"0c001820",
			4565 => x"01001018",
			4566 => x"04002010",
			4567 => x"0b00150c",
			4568 => x"00012708",
			4569 => x"03002904",
			4570 => x"fe9347e5",
			4571 => x"fffb47e5",
			4572 => x"010b47e5",
			4573 => x"fe4f47e5",
			4574 => x"06009804",
			4575 => x"01b347e5",
			4576 => x"00cb47e5",
			4577 => x"0000c704",
			4578 => x"fede47e5",
			4579 => x"018147e5",
			4580 => x"0d001a14",
			4581 => x"01001210",
			4582 => x"0600b10c",
			4583 => x"03002708",
			4584 => x"0b001804",
			4585 => x"00e947e5",
			4586 => x"fedd47e5",
			4587 => x"fe4c47e5",
			4588 => x"ffde47e5",
			4589 => x"001447e5",
			4590 => x"0c002314",
			4591 => x"04001d04",
			4592 => x"fe5347e5",
			4593 => x"04002108",
			4594 => x"07003904",
			4595 => x"ffe347e5",
			4596 => x"01e347e5",
			4597 => x"08002404",
			4598 => x"013747e5",
			4599 => x"ffea47e5",
			4600 => x"fe8d47e5",
			4601 => x"01001028",
			4602 => x"07002a0c",
			4603 => x"0e007a08",
			4604 => x"07002904",
			4605 => x"ffd548b1",
			4606 => x"001448b1",
			4607 => x"003f48b1",
			4608 => x"08002418",
			4609 => x"0d001a10",
			4610 => x"06007f04",
			4611 => x"001048b1",
			4612 => x"03002104",
			4613 => x"001048b1",
			4614 => x"0e009f04",
			4615 => x"ff7148b1",
			4616 => x"fff848b1",
			4617 => x"03003304",
			4618 => x"ffdc48b1",
			4619 => x"002c48b1",
			4620 => x"001348b1",
			4621 => x"0c00190c",
			4622 => x"0b001508",
			4623 => x"05002804",
			4624 => x"000348b1",
			4625 => x"ffe448b1",
			4626 => x"006c48b1",
			4627 => x"09002204",
			4628 => x"ff9448b1",
			4629 => x"08002614",
			4630 => x"07003c0c",
			4631 => x"00012508",
			4632 => x"04001f04",
			4633 => x"001f48b1",
			4634 => x"ffd248b1",
			4635 => x"007548b1",
			4636 => x"00012804",
			4637 => x"001c48b1",
			4638 => x"ffc248b1",
			4639 => x"03002e0c",
			4640 => x"02013708",
			4641 => x"0a002d04",
			4642 => x"002748b1",
			4643 => x"ffaf48b1",
			4644 => x"005048b1",
			4645 => x"0a003b08",
			4646 => x"02011304",
			4647 => x"000e48b1",
			4648 => x"ff7a48b1",
			4649 => x"0600b704",
			4650 => x"003548b1",
			4651 => x"ffe848b1",
			4652 => x"05002714",
			4653 => x"07002908",
			4654 => x"07002804",
			4655 => x"ffe2498d",
			4656 => x"0031498d",
			4657 => x"04001e08",
			4658 => x"0e00a104",
			4659 => x"ff64498d",
			4660 => x"fffb498d",
			4661 => x"0003498d",
			4662 => x"0b001720",
			4663 => x"0300321c",
			4664 => x"08001d10",
			4665 => x"0001450c",
			4666 => x"0000c508",
			4667 => x"00009304",
			4668 => x"fffb498d",
			4669 => x"002d498d",
			4670 => x"ff87498d",
			4671 => x"0051498d",
			4672 => x"0000c704",
			4673 => x"ffee498d",
			4674 => x"0e009b04",
			4675 => x"00b4498d",
			4676 => x"fffa498d",
			4677 => x"ffc5498d",
			4678 => x"08002210",
			4679 => x"05002a04",
			4680 => x"003f498d",
			4681 => x"04002804",
			4682 => x"ff3e498d",
			4683 => x"09002204",
			4684 => x"0021498d",
			4685 => x"ffe3498d",
			4686 => x"0201371c",
			4687 => x"0a003b10",
			4688 => x"04002108",
			4689 => x"0e008604",
			4690 => x"ff9b498d",
			4691 => x"0063498d",
			4692 => x"08002404",
			4693 => x"000d498d",
			4694 => x"ff4a498d",
			4695 => x"00012804",
			4696 => x"ffda498d",
			4697 => x"07003f04",
			4698 => x"006d498d",
			4699 => x"fff4498d",
			4700 => x"01001908",
			4701 => x"03003104",
			4702 => x"00d4498d",
			4703 => x"000b498d",
			4704 => x"0f00e204",
			4705 => x"ffb6498d",
			4706 => x"000e498d",
			4707 => x"08002048",
			4708 => x"0b001314",
			4709 => x"0d001104",
			4710 => x"feb94a89",
			4711 => x"0e00910c",
			4712 => x"08001b04",
			4713 => x"ff954a89",
			4714 => x"06004b04",
			4715 => x"ffd44a89",
			4716 => x"01bc4a89",
			4717 => x"00064a89",
			4718 => x"05002e18",
			4719 => x"09001f10",
			4720 => x"0001470c",
			4721 => x"01000e04",
			4722 => x"fe844a89",
			4723 => x"0600a104",
			4724 => x"01524a89",
			4725 => x"feb34a89",
			4726 => x"008b4a89",
			4727 => x"04001e04",
			4728 => x"ff2b4a89",
			4729 => x"018e4a89",
			4730 => x"07003614",
			4731 => x"05003808",
			4732 => x"09001b04",
			4733 => x"ffcf4a89",
			4734 => x"fe564a89",
			4735 => x"0b001508",
			4736 => x"0a003704",
			4737 => x"00ed4a89",
			4738 => x"ffa34a89",
			4739 => x"fecf4a89",
			4740 => x"07003804",
			4741 => x"00c04a89",
			4742 => x"fef44a89",
			4743 => x"07003518",
			4744 => x"0c001c14",
			4745 => x"02012a10",
			4746 => x"0400260c",
			4747 => x"07002a08",
			4748 => x"00008f04",
			4749 => x"ffdb4a89",
			4750 => x"01504a89",
			4751 => x"ff8d4a89",
			4752 => x"015a4a89",
			4753 => x"01794a89",
			4754 => x"fe974a89",
			4755 => x"03002908",
			4756 => x"01001604",
			4757 => x"ff214a89",
			4758 => x"01734a89",
			4759 => x"05003304",
			4760 => x"fe9b4a89",
			4761 => x"02011904",
			4762 => x"fe6b4a89",
			4763 => x"09002508",
			4764 => x"03003304",
			4765 => x"ff594a89",
			4766 => x"007a4a89",
			4767 => x"05003804",
			4768 => x"01534a89",
			4769 => x"ffba4a89",
			4770 => x"01000a04",
			4771 => x"fefd4b25",
			4772 => x"02013f40",
			4773 => x"08001f14",
			4774 => x"0c00150c",
			4775 => x"07002c08",
			4776 => x"0d001304",
			4777 => x"ffe84b25",
			4778 => x"00d14b25",
			4779 => x"ff5d4b25",
			4780 => x"01001004",
			4781 => x"fed64b25",
			4782 => x"ffdd4b25",
			4783 => x"0800271c",
			4784 => x"05002e0c",
			4785 => x"05002704",
			4786 => x"ff554b25",
			4787 => x"0d001604",
			4788 => x"000f4b25",
			4789 => x"00ef4b25",
			4790 => x"03002f08",
			4791 => x"0f00bc04",
			4792 => x"009c4b25",
			4793 => x"ff244b25",
			4794 => x"01001204",
			4795 => x"ffc64b25",
			4796 => x"008a4b25",
			4797 => x"00013d04",
			4798 => x"feea4b25",
			4799 => x"0c002004",
			4800 => x"ff8e4b25",
			4801 => x"09002b04",
			4802 => x"00a24b25",
			4803 => x"ff7d4b25",
			4804 => x"0d002108",
			4805 => x"0e00a604",
			4806 => x"01244b25",
			4807 => x"ffe54b25",
			4808 => x"ff4a4b25",
			4809 => x"05002404",
			4810 => x"fec14bd9",
			4811 => x"05002e20",
			4812 => x"08001d0c",
			4813 => x"01000e08",
			4814 => x"00014604",
			4815 => x"fec14bd9",
			4816 => x"ffbf4bd9",
			4817 => x"00a74bd9",
			4818 => x"03002a10",
			4819 => x"0a002808",
			4820 => x"0d001704",
			4821 => x"00d84bd9",
			4822 => x"fefc4bd9",
			4823 => x"0f00c404",
			4824 => x"005f4bd9",
			4825 => x"014e4bd9",
			4826 => x"ff674bd9",
			4827 => x"08002018",
			4828 => x"0b001304",
			4829 => x"00e04bd9",
			4830 => x"0700360c",
			4831 => x"05003804",
			4832 => x"fe8c4bd9",
			4833 => x"04002a04",
			4834 => x"00684bd9",
			4835 => x"ff414bd9",
			4836 => x"07003804",
			4837 => x"008d4bd9",
			4838 => x"ff524bd9",
			4839 => x"0b001808",
			4840 => x"00012504",
			4841 => x"ffb14bd9",
			4842 => x"01004bd9",
			4843 => x"0d001a08",
			4844 => x"0600a704",
			4845 => x"fe994bd9",
			4846 => x"ffab4bd9",
			4847 => x"05003308",
			4848 => x"03002e04",
			4849 => x"fff64bd9",
			4850 => x"feaf4bd9",
			4851 => x"05003404",
			4852 => x"010f4bd9",
			4853 => x"00064bd9",
			4854 => x"08001c04",
			4855 => x"fe684c5d",
			4856 => x"0f008004",
			4857 => x"fe714c5d",
			4858 => x"0b001718",
			4859 => x"04001808",
			4860 => x"0d001404",
			4861 => x"00964c5d",
			4862 => x"fee64c5d",
			4863 => x"08001d04",
			4864 => x"ffdd4c5d",
			4865 => x"0d001708",
			4866 => x"0d001504",
			4867 => x"01264c5d",
			4868 => x"02144c5d",
			4869 => x"00c44c5d",
			4870 => x"08002210",
			4871 => x"0a004f0c",
			4872 => x"06009a08",
			4873 => x"0e007a04",
			4874 => x"feb84c5d",
			4875 => x"006a4c5d",
			4876 => x"fe314c5d",
			4877 => x"01234c5d",
			4878 => x"0d002210",
			4879 => x"02013708",
			4880 => x"0a003b04",
			4881 => x"000e4c5d",
			4882 => x"015c4c5d",
			4883 => x"05003904",
			4884 => x"01f44c5d",
			4885 => x"00024c5d",
			4886 => x"fe644c5d",
			4887 => x"07004064",
			4888 => x"08002030",
			4889 => x"0c001828",
			4890 => x"0400231c",
			4891 => x"01000e10",
			4892 => x"0f00d808",
			4893 => x"0b001304",
			4894 => x"001e4d41",
			4895 => x"fed74d41",
			4896 => x"09001904",
			4897 => x"ffab4d41",
			4898 => x"00ab4d41",
			4899 => x"06009504",
			4900 => x"ff8c4d41",
			4901 => x"0e009d04",
			4902 => x"009f4d41",
			4903 => x"ffea4d41",
			4904 => x"06007404",
			4905 => x"ffd24d41",
			4906 => x"05003904",
			4907 => x"00db4d41",
			4908 => x"ffee4d41",
			4909 => x"0b001604",
			4910 => x"003d4d41",
			4911 => x"fee84d41",
			4912 => x"00011f1c",
			4913 => x"0200fd14",
			4914 => x"0a002d0c",
			4915 => x"03002108",
			4916 => x"04001a04",
			4917 => x"ffe54d41",
			4918 => x"00744d41",
			4919 => x"ff374d41",
			4920 => x"05003404",
			4921 => x"00df4d41",
			4922 => x"ffbb4d41",
			4923 => x"0a003604",
			4924 => x"ff094d41",
			4925 => x"ffe04d41",
			4926 => x"04002004",
			4927 => x"ffde4d41",
			4928 => x"04002104",
			4929 => x"013c4d41",
			4930 => x"07003708",
			4931 => x"00013104",
			4932 => x"00d74d41",
			4933 => x"003d4d41",
			4934 => x"0b001e04",
			4935 => x"ff864d41",
			4936 => x"00854d41",
			4937 => x"0c002104",
			4938 => x"ff0e4d41",
			4939 => x"00014904",
			4940 => x"ff884d41",
			4941 => x"02014204",
			4942 => x"00854d41",
			4943 => x"ffbd4d41",
			4944 => x"08001b04",
			4945 => x"fe834ded",
			4946 => x"0b00130c",
			4947 => x"05002404",
			4948 => x"fea54ded",
			4949 => x"07002b04",
			4950 => x"02114ded",
			4951 => x"00c64ded",
			4952 => x"08002024",
			4953 => x"05002e14",
			4954 => x"04001d08",
			4955 => x"0f00d804",
			4956 => x"fe744ded",
			4957 => x"00a54ded",
			4958 => x"01000e08",
			4959 => x"0b001504",
			4960 => x"00b24ded",
			4961 => x"fe924ded",
			4962 => x"01654ded",
			4963 => x"07003608",
			4964 => x"09001c04",
			4965 => x"ff814ded",
			4966 => x"fe4a4ded",
			4967 => x"07003804",
			4968 => x"00d34ded",
			4969 => x"fea44ded",
			4970 => x"0c001808",
			4971 => x"0000c704",
			4972 => x"ff2b4ded",
			4973 => x"01694ded",
			4974 => x"04001d0c",
			4975 => x"04001608",
			4976 => x"0d001904",
			4977 => x"006b4ded",
			4978 => x"ff3c4ded",
			4979 => x"fe214ded",
			4980 => x"04002108",
			4981 => x"0e008604",
			4982 => x"fe5b4ded",
			4983 => x"017e4ded",
			4984 => x"07003404",
			4985 => x"010c4ded",
			4986 => x"ffd34ded",
			4987 => x"0f008004",
			4988 => x"fe6f4e61",
			4989 => x"08001b04",
			4990 => x"fe794e61",
			4991 => x"07002a04",
			4992 => x"01f84e61",
			4993 => x"02012614",
			4994 => x"08002710",
			4995 => x"0600a108",
			4996 => x"0f00aa04",
			4997 => x"ff214e61",
			4998 => x"01564e61",
			4999 => x"04002604",
			5000 => x"feee4e61",
			5001 => x"00fa4e61",
			5002 => x"fe6c4e61",
			5003 => x"0a00310c",
			5004 => x"03002a08",
			5005 => x"04001e04",
			5006 => x"ffcb4e61",
			5007 => x"015d4e61",
			5008 => x"feac4e61",
			5009 => x"04002108",
			5010 => x"08002004",
			5011 => x"ffd24e61",
			5012 => x"02384e61",
			5013 => x"08002a04",
			5014 => x"004c4e61",
			5015 => x"01c54e61",
			5016 => x"0201495c",
			5017 => x"0600bb4c",
			5018 => x"0c00181c",
			5019 => x"08001d10",
			5020 => x"0b001308",
			5021 => x"09001a04",
			5022 => x"ffcb4f1d",
			5023 => x"00614f1d",
			5024 => x"07003304",
			5025 => x"ff644f1d",
			5026 => x"00224f1d",
			5027 => x"0000c704",
			5028 => x"ffb44f1d",
			5029 => x"0f00c904",
			5030 => x"00b84f1d",
			5031 => x"00024f1d",
			5032 => x"0a003b20",
			5033 => x"07003910",
			5034 => x"00012a08",
			5035 => x"00012104",
			5036 => x"ffa44f1d",
			5037 => x"004a4f1d",
			5038 => x"08002404",
			5039 => x"ff094f1d",
			5040 => x"ffc74f1d",
			5041 => x"08002708",
			5042 => x"0e009104",
			5043 => x"00014f1d",
			5044 => x"00844f1d",
			5045 => x"08002d04",
			5046 => x"ff4f4f1d",
			5047 => x"00524f1d",
			5048 => x"00013a0c",
			5049 => x"0f00bb08",
			5050 => x"02011704",
			5051 => x"ffd14f1d",
			5052 => x"00704f1d",
			5053 => x"ff974f1d",
			5054 => x"00a54f1d",
			5055 => x"0f00d404",
			5056 => x"fff74f1d",
			5057 => x"01001a04",
			5058 => x"ff3f4f1d",
			5059 => x"01001f04",
			5060 => x"000b4f1d",
			5061 => x"fff04f1d",
			5062 => x"00814f1d",
			5063 => x"0d00226c",
			5064 => x"01001240",
			5065 => x"0c001824",
			5066 => x"01001020",
			5067 => x"0b001410",
			5068 => x"0d001208",
			5069 => x"05002804",
			5070 => x"ff214ff9",
			5071 => x"003d4ff9",
			5072 => x"0000be04",
			5073 => x"ff914ff9",
			5074 => x"00f94ff9",
			5075 => x"0e008e08",
			5076 => x"03002604",
			5077 => x"ffb24ff9",
			5078 => x"fe904ff9",
			5079 => x"0d001504",
			5080 => x"ff964ff9",
			5081 => x"01194ff9",
			5082 => x"00e44ff9",
			5083 => x"0d001a0c",
			5084 => x"0f00cc08",
			5085 => x"0b001604",
			5086 => x"00184ff9",
			5087 => x"fe844ff9",
			5088 => x"ffbc4ff9",
			5089 => x"09002408",
			5090 => x"03002704",
			5091 => x"ff834ff9",
			5092 => x"012c4ff9",
			5093 => x"07003f04",
			5094 => x"ff334ff9",
			5095 => x"005b4ff9",
			5096 => x"07003710",
			5097 => x"09002108",
			5098 => x"05002d04",
			5099 => x"006a4ff9",
			5100 => x"ffaf4ff9",
			5101 => x"0f00b004",
			5102 => x"ff394ff9",
			5103 => x"016e4ff9",
			5104 => x"05003810",
			5105 => x"0500360c",
			5106 => x"00014308",
			5107 => x"04002304",
			5108 => x"000c4ff9",
			5109 => x"fe904ff9",
			5110 => x"00f44ff9",
			5111 => x"01284ff9",
			5112 => x"03003b08",
			5113 => x"00014804",
			5114 => x"fea04ff9",
			5115 => x"fff14ff9",
			5116 => x"00ae4ff9",
			5117 => x"febf4ff9",
			5118 => x"08001c04",
			5119 => x"fe7850df",
			5120 => x"0c001824",
			5121 => x"05002408",
			5122 => x"08001d04",
			5123 => x"009f50df",
			5124 => x"fe9250df",
			5125 => x"01001014",
			5126 => x"0b001408",
			5127 => x"04001c04",
			5128 => x"00e750df",
			5129 => x"01bf50df",
			5130 => x"0e008e08",
			5131 => x"03002604",
			5132 => x"004650df",
			5133 => x"fe5750df",
			5134 => x"010150df",
			5135 => x"0000c704",
			5136 => x"ff0650df",
			5137 => x"018850df",
			5138 => x"0800221c",
			5139 => x"09001e08",
			5140 => x"08001d04",
			5141 => x"fef550df",
			5142 => x"00f450df",
			5143 => x"0a004f0c",
			5144 => x"03002708",
			5145 => x"03002404",
			5146 => x"fed450df",
			5147 => x"007450df",
			5148 => x"fe5350df",
			5149 => x"07003504",
			5150 => x"010650df",
			5151 => x"ff9250df",
			5152 => x"04001d10",
			5153 => x"0400160c",
			5154 => x"04001504",
			5155 => x"ff8450df",
			5156 => x"01001204",
			5157 => x"ffda50df",
			5158 => x"006a50df",
			5159 => x"fe4850df",
			5160 => x"05003710",
			5161 => x"0f00c008",
			5162 => x"0f00b304",
			5163 => x"013d50df",
			5164 => x"ff3d50df",
			5165 => x"05003304",
			5166 => x"002450df",
			5167 => x"014950df",
			5168 => x"0a003b08",
			5169 => x"00014804",
			5170 => x"fe6750df",
			5171 => x"002f50df",
			5172 => x"07003804",
			5173 => x"01a350df",
			5174 => x"ff9550df",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1711, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3455, initial_addr_3'length));
	end generate gen_rom_5;

	gen_rom_6: if SELECT_ROM = 6 generate
		bank <= (
			0 => x"0e00920c",
			1 => x"0d001008",
			2 => x"0d000f04",
			3 => x"fffa003d",
			4 => x"000f003d",
			5 => x"ffba003d",
			6 => x"0e009e08",
			7 => x"05002a04",
			8 => x"007a003d",
			9 => x"ffe9003d",
			10 => x"07003404",
			11 => x"ffc2003d",
			12 => x"07003804",
			13 => x"004a003d",
			14 => x"ffe5003d",
			15 => x"0e009b10",
			16 => x"0c001308",
			17 => x"04001b04",
			18 => x"00290081",
			19 => x"fffa0081",
			20 => x"04001404",
			21 => x"00030081",
			22 => x"ffa20081",
			23 => x"08001d08",
			24 => x"0600ca04",
			25 => x"00690081",
			26 => x"00000081",
			27 => x"0a003204",
			28 => x"ffd10081",
			29 => x"04002304",
			30 => x"00260081",
			31 => x"fff50081",
			32 => x"0e00920c",
			33 => x"0c001308",
			34 => x"0c001204",
			35 => x"fff400bd",
			36 => x"001f00bd",
			37 => x"ff8900bd",
			38 => x"01000a04",
			39 => x"ffe200bd",
			40 => x"0700380c",
			41 => x"05002e08",
			42 => x"07003304",
			43 => x"002e00bd",
			44 => x"009600bd",
			45 => x"ffe300bd",
			46 => x"ffc700bd",
			47 => x"0e00920c",
			48 => x"0c001308",
			49 => x"0c001204",
			50 => x"fffb0101",
			51 => x"00100101",
			52 => x"ffc30101",
			53 => x"0e00a410",
			54 => x"03002f0c",
			55 => x"07003608",
			56 => x"04001d04",
			57 => x"00770101",
			58 => x"00080101",
			59 => x"fff60101",
			60 => x"ffd80101",
			61 => x"03002e04",
			62 => x"ffc70101",
			63 => x"00300101",
			64 => x"0e009104",
			65 => x"fef0013d",
			66 => x"0e009408",
			67 => x"05002904",
			68 => x"012a013d",
			69 => x"ff95013d",
			70 => x"03002a08",
			71 => x"03002704",
			72 => x"000a013d",
			73 => x"ff29013d",
			74 => x"0c001504",
			75 => x"ffc5013d",
			76 => x"05002e04",
			77 => x"0131013d",
			78 => x"ff77013d",
			79 => x"01000a14",
			80 => x"0400140c",
			81 => x"08001d08",
			82 => x"07002a04",
			83 => x"ffff0191",
			84 => x"00340191",
			85 => x"fff70191",
			86 => x"05001f04",
			87 => x"00030191",
			88 => x"ffaa0191",
			89 => x"03002608",
			90 => x"0c001304",
			91 => x"001f0191",
			92 => x"ffc60191",
			93 => x"05002e0c",
			94 => x"0e00a408",
			95 => x"0f00bf04",
			96 => x"fff20191",
			97 => x"00860191",
			98 => x"fffd0191",
			99 => x"ffdf0191",
			100 => x"0600b10c",
			101 => x"0600ad04",
			102 => x"fe5f01dd",
			103 => x"0a002f04",
			104 => x"04a701dd",
			105 => x"fe6601dd",
			106 => x"05002d14",
			107 => x"09001804",
			108 => x"069801dd",
			109 => x"0001490c",
			110 => x"0600bb04",
			111 => x"06cc01dd",
			112 => x"0e00a304",
			113 => x"03da01dd",
			114 => x"022301dd",
			115 => x"fe0901dd",
			116 => x"02012104",
			117 => x"00a801dd",
			118 => x"fe5101dd",
			119 => x"0f00ca10",
			120 => x"0500250c",
			121 => x"04001804",
			122 => x"fff00231",
			123 => x"08001b04",
			124 => x"fffb0231",
			125 => x"004e0231",
			126 => x"ff7d0231",
			127 => x"0f00e314",
			128 => x"02012f10",
			129 => x"0d001508",
			130 => x"05002504",
			131 => x"00030231",
			132 => x"00b60231",
			133 => x"03002e04",
			134 => x"ffd10231",
			135 => x"ffff0231",
			136 => x"ffc00231",
			137 => x"03002e04",
			138 => x"ff9c0231",
			139 => x"00320231",
			140 => x"0b001310",
			141 => x"00011704",
			142 => x"ffc9028d",
			143 => x"01000704",
			144 => x"ffe3028d",
			145 => x"0c001404",
			146 => x"0070028d",
			147 => x"ffee028d",
			148 => x"02010b10",
			149 => x"04001808",
			150 => x"01000904",
			151 => x"0015028d",
			152 => x"ffc7028d",
			153 => x"0f00bc04",
			154 => x"ffea028d",
			155 => x"0060028d",
			156 => x"03002e04",
			157 => x"ff93028d",
			158 => x"08001d04",
			159 => x"002d028d",
			160 => x"03002f04",
			161 => x"000f028d",
			162 => x"ffd3028d",
			163 => x"0e009104",
			164 => x"fe7502c9",
			165 => x"07003818",
			166 => x"0700330c",
			167 => x"0b001304",
			168 => x"009b02c9",
			169 => x"05002704",
			170 => x"feea02c9",
			171 => x"00a102c9",
			172 => x"05002e08",
			173 => x"0d001404",
			174 => x"01a502c9",
			175 => x"00a002c9",
			176 => x"fee102c9",
			177 => x"fe9802c9",
			178 => x"0b001310",
			179 => x"00011704",
			180 => x"ffc10325",
			181 => x"01000704",
			182 => x"ffde0325",
			183 => x"0e009104",
			184 => x"ffff0325",
			185 => x"00a90325",
			186 => x"02010b0c",
			187 => x"08001c04",
			188 => x"ffc40325",
			189 => x"0f00bc04",
			190 => x"ffe90325",
			191 => x"006d0325",
			192 => x"04001704",
			193 => x"00030325",
			194 => x"01001208",
			195 => x"0a003604",
			196 => x"ff8e0325",
			197 => x"00080325",
			198 => x"08002304",
			199 => x"000f0325",
			200 => x"fff60325",
			201 => x"0f00d924",
			202 => x"07003214",
			203 => x"0d00140c",
			204 => x"0d001108",
			205 => x"0d000f04",
			206 => x"fffa0389",
			207 => x"000e0389",
			208 => x"ffa20389",
			209 => x"09001c04",
			210 => x"00180389",
			211 => x"fff60389",
			212 => x"0d001404",
			213 => x"00430389",
			214 => x"0a003204",
			215 => x"ffb50389",
			216 => x"04002004",
			217 => x"002e0389",
			218 => x"ffed0389",
			219 => x"02014708",
			220 => x"0600ca04",
			221 => x"005f0389",
			222 => x"00050389",
			223 => x"0600cb04",
			224 => x"ffd50389",
			225 => x"00040389",
			226 => x"0600ab04",
			227 => x"fe6303c5",
			228 => x"05002e18",
			229 => x"0b001308",
			230 => x"07002f04",
			231 => x"035603c5",
			232 => x"016d03c5",
			233 => x"03002604",
			234 => x"fe1d03c5",
			235 => x"07003204",
			236 => x"ffae03c5",
			237 => x"0d001504",
			238 => x"037f03c5",
			239 => x"00e003c5",
			240 => x"fe6103c5",
			241 => x"03002a24",
			242 => x"0b001314",
			243 => x"0f00d810",
			244 => x"0d001108",
			245 => x"01000a04",
			246 => x"fff70429",
			247 => x"00140429",
			248 => x"09001804",
			249 => x"00120429",
			250 => x"ff8d0429",
			251 => x"00610429",
			252 => x"0201060c",
			253 => x"0d001408",
			254 => x"08001d04",
			255 => x"ffe90429",
			256 => x"00650429",
			257 => x"ffde0429",
			258 => x"ff680429",
			259 => x"0200f704",
			260 => x"ffae0429",
			261 => x"05002e08",
			262 => x"0e008a04",
			263 => x"fffb0429",
			264 => x"00d80429",
			265 => x"ffcc0429",
			266 => x"0200f704",
			267 => x"ffa60475",
			268 => x"03002a1c",
			269 => x"07002f0c",
			270 => x"09001908",
			271 => x"05002704",
			272 => x"00520475",
			273 => x"fff80475",
			274 => x"ffe00475",
			275 => x"0600bd08",
			276 => x"00012704",
			277 => x"002c0475",
			278 => x"ffe90475",
			279 => x"04001d04",
			280 => x"ffa20475",
			281 => x"000c0475",
			282 => x"05002d04",
			283 => x"00960475",
			284 => x"ffd10475",
			285 => x"0600ab04",
			286 => x"fe6804c9",
			287 => x"00013010",
			288 => x"0700380c",
			289 => x"04001a08",
			290 => x"0600bd04",
			291 => x"018304c9",
			292 => x"007104c9",
			293 => x"025704c9",
			294 => x"fe6704c9",
			295 => x"0700300c",
			296 => x"09001904",
			297 => x"01d304c9",
			298 => x"00014404",
			299 => x"ffdb04c9",
			300 => x"fe3b04c9",
			301 => x"0e00ac08",
			302 => x"0600c504",
			303 => x"fe6d04c9",
			304 => x"fddb04c9",
			305 => x"00a004c9",
			306 => x"0600be2c",
			307 => x"08001c18",
			308 => x"09001808",
			309 => x"0d001104",
			310 => x"fff5053d",
			311 => x"0015053d",
			312 => x"0d001108",
			313 => x"04001804",
			314 => x"fff8053d",
			315 => x"0012053d",
			316 => x"0a003404",
			317 => x"ffa3053d",
			318 => x"000d053d",
			319 => x"01000b08",
			320 => x"0f00bf04",
			321 => x"fff3053d",
			322 => x"0041053d",
			323 => x"05002904",
			324 => x"ffc6053d",
			325 => x"05002b04",
			326 => x"0023053d",
			327 => x"fff2053d",
			328 => x"0b001304",
			329 => x"005f053d",
			330 => x"0f00e708",
			331 => x"05002e04",
			332 => x"0024053d",
			333 => x"fff4053d",
			334 => x"ffe0053d",
			335 => x"0600ab04",
			336 => x"fe650581",
			337 => x"0c00171c",
			338 => x"03002a10",
			339 => x"0b001304",
			340 => x"01770581",
			341 => x"0f00d508",
			342 => x"0a002d04",
			343 => x"fe7e0581",
			344 => x"01fa0581",
			345 => x"fe630581",
			346 => x"0e009604",
			347 => x"05df0581",
			348 => x"07003404",
			349 => x"00a00581",
			350 => x"023b0581",
			351 => x"fe6d0581",
			352 => x"0600ab04",
			353 => x"fe6605dd",
			354 => x"00013014",
			355 => x"03002a08",
			356 => x"0d001404",
			357 => x"015905dd",
			358 => x"fef605dd",
			359 => x"0d001504",
			360 => x"02d305dd",
			361 => x"0f00c704",
			362 => x"feb505dd",
			363 => x"00e205dd",
			364 => x"0700300c",
			365 => x"09001904",
			366 => x"01ff05dd",
			367 => x"00014404",
			368 => x"000b05dd",
			369 => x"fe2705dd",
			370 => x"0e00ac08",
			371 => x"0600c504",
			372 => x"fe6c05dd",
			373 => x"fd8405dd",
			374 => x"00b805dd",
			375 => x"0c001620",
			376 => x"07003218",
			377 => x"02010c04",
			378 => x"ff6b0641",
			379 => x"0f00e310",
			380 => x"0c00140c",
			381 => x"08001804",
			382 => x"ffda0641",
			383 => x"0e008a04",
			384 => x"fff80641",
			385 => x"00be0641",
			386 => x"ffbd0641",
			387 => x"ffbb0641",
			388 => x"0a002f04",
			389 => x"00110641",
			390 => x"00930641",
			391 => x"03002e04",
			392 => x"ff910641",
			393 => x"03003108",
			394 => x"0e009404",
			395 => x"fff70641",
			396 => x"002d0641",
			397 => x"0600c304",
			398 => x"ffd50641",
			399 => x"00010641",
			400 => x"0200f704",
			401 => x"fe82069d",
			402 => x"0001301c",
			403 => x"0d001510",
			404 => x"03002404",
			405 => x"febb069d",
			406 => x"05002d08",
			407 => x"0600ab04",
			408 => x"ffa0069d",
			409 => x"019d069d",
			410 => x"ff56069d",
			411 => x"0a003204",
			412 => x"fe75069d",
			413 => x"04002304",
			414 => x"0129069d",
			415 => x"ff4b069d",
			416 => x"0b001308",
			417 => x"05002704",
			418 => x"00bc069d",
			419 => x"fef8069d",
			420 => x"0600cc04",
			421 => x"fea0069d",
			422 => x"ffea069d",
			423 => x"0e008a04",
			424 => x"fe700701",
			425 => x"0d001518",
			426 => x"0001310c",
			427 => x"0000f804",
			428 => x"febe0701",
			429 => x"03002a04",
			430 => x"00c50701",
			431 => x"01d80701",
			432 => x"0b001304",
			433 => x"00c90701",
			434 => x"01000904",
			435 => x"ff270701",
			436 => x"fe1d0701",
			437 => x"0e00a00c",
			438 => x"0e009e08",
			439 => x"0e009c04",
			440 => x"fe910701",
			441 => x"00850701",
			442 => x"fd690701",
			443 => x"03002e04",
			444 => x"fe450701",
			445 => x"04002604",
			446 => x"01900701",
			447 => x"ff330701",
			448 => x"00013028",
			449 => x"05002310",
			450 => x"03002a0c",
			451 => x"09001808",
			452 => x"07002804",
			453 => x"fff00785",
			454 => x"00340785",
			455 => x"ff0f0785",
			456 => x"00680785",
			457 => x"05002e14",
			458 => x"01000b0c",
			459 => x"03002604",
			460 => x"ffb60785",
			461 => x"0f00bf04",
			462 => x"ffe10785",
			463 => x"01410785",
			464 => x"0600b104",
			465 => x"ff530785",
			466 => x"00840785",
			467 => x"ff5e0785",
			468 => x"07003014",
			469 => x"09001908",
			470 => x"05002704",
			471 => x"01050785",
			472 => x"ffac0785",
			473 => x"03002a04",
			474 => x"ff3d0785",
			475 => x"00013c04",
			476 => x"002f0785",
			477 => x"fff40785",
			478 => x"0e00ac04",
			479 => x"fee20785",
			480 => x"00300785",
			481 => x"03002a2c",
			482 => x"0900180c",
			483 => x"01000704",
			484 => x"ff550809",
			485 => x"03002104",
			486 => x"ffe60809",
			487 => x"014e0809",
			488 => x"0001120c",
			489 => x"07003304",
			490 => x"fef00809",
			491 => x"05002304",
			492 => x"ff850809",
			493 => x"01410809",
			494 => x"0b001308",
			495 => x"0f00cb04",
			496 => x"ff170809",
			497 => x"ffd60809",
			498 => x"04001e04",
			499 => x"fe780809",
			500 => x"04002004",
			501 => x"00410809",
			502 => x"ff4b0809",
			503 => x"0200f704",
			504 => x"fec30809",
			505 => x"00013008",
			506 => x"05002e04",
			507 => x"01860809",
			508 => x"ff280809",
			509 => x"01000e08",
			510 => x"0f00d004",
			511 => x"ff730809",
			512 => x"00b20809",
			513 => x"fede0809",
			514 => x"04001c2c",
			515 => x"0300240c",
			516 => x"09001708",
			517 => x"0000c204",
			518 => x"ffc70875",
			519 => x"00f30875",
			520 => x"fe990875",
			521 => x"0600bd18",
			522 => x"00012714",
			523 => x"0400180c",
			524 => x"04001508",
			525 => x"0d001704",
			526 => x"01040875",
			527 => x"ffdb0875",
			528 => x"fed50875",
			529 => x"0000f404",
			530 => x"ffb80875",
			531 => x"01b90875",
			532 => x"ffab0875",
			533 => x"07003304",
			534 => x"ff6a0875",
			535 => x"00c40875",
			536 => x"0e009b04",
			537 => x"fe920875",
			538 => x"05003204",
			539 => x"006e0875",
			540 => x"ff9b0875",
			541 => x"05002514",
			542 => x"03002608",
			543 => x"0c001304",
			544 => x"003708f9",
			545 => x"ffb108f9",
			546 => x"00011508",
			547 => x"01000b04",
			548 => x"000608f9",
			549 => x"fff708f9",
			550 => x"009108f9",
			551 => x"0f00e328",
			552 => x"0f00ca14",
			553 => x"01000908",
			554 => x"01000804",
			555 => x"fff108f9",
			556 => x"002208f9",
			557 => x"03002e04",
			558 => x"ff9508f9",
			559 => x"0a003204",
			560 => x"001d08f9",
			561 => x"ffe808f9",
			562 => x"0d001508",
			563 => x"00013d04",
			564 => x"009308f9",
			565 => x"ffe108f9",
			566 => x"0a003204",
			567 => x"ffbf08f9",
			568 => x"04002104",
			569 => x"002c08f9",
			570 => x"ffee08f9",
			571 => x"0a003404",
			572 => x"ffa008f9",
			573 => x"000608f9",
			574 => x"0f00bf04",
			575 => x"fe80093d",
			576 => x"01000804",
			577 => x"fe7a093d",
			578 => x"0d001204",
			579 => x"01b1093d",
			580 => x"00014910",
			581 => x"0700380c",
			582 => x"00011e04",
			583 => x"fffc093d",
			584 => x"0f00cc04",
			585 => x"fedc093d",
			586 => x"0140093d",
			587 => x"fea6093d",
			588 => x"0600cb04",
			589 => x"fe85093d",
			590 => x"ffc4093d",
			591 => x"01000b28",
			592 => x"0100080c",
			593 => x"04001004",
			594 => x"002309c1",
			595 => x"07003304",
			596 => x"ff9109c1",
			597 => x"fffe09c1",
			598 => x"08001804",
			599 => x"ffcd09c1",
			600 => x"0a00320c",
			601 => x"0f00bf04",
			602 => x"ffdf09c1",
			603 => x"03002604",
			604 => x"fff909c1",
			605 => x"00e409c1",
			606 => x"07003204",
			607 => x"ffa909c1",
			608 => x"08001f04",
			609 => x"004d09c1",
			610 => x"000009c1",
			611 => x"0a003214",
			612 => x"09001804",
			613 => x"003309c1",
			614 => x"09001c04",
			615 => x"ff4b09c1",
			616 => x"0b001608",
			617 => x"08001f04",
			618 => x"fff409c1",
			619 => x"002909c1",
			620 => x"ffec09c1",
			621 => x"05002f04",
			622 => x"005609c1",
			623 => x"ffd409c1",
			624 => x"00013030",
			625 => x"07003010",
			626 => x"0d001108",
			627 => x"07002b04",
			628 => x"fffb0a4d",
			629 => x"001a0a4d",
			630 => x"09001804",
			631 => x"000c0a4d",
			632 => x"ffb50a4d",
			633 => x"03002604",
			634 => x"ffd40a4d",
			635 => x"0d00150c",
			636 => x"01000a04",
			637 => x"fff10a4d",
			638 => x"0f00bf04",
			639 => x"ffee0a4d",
			640 => x"009f0a4d",
			641 => x"08001d04",
			642 => x"001f0a4d",
			643 => x"01001208",
			644 => x"0a003604",
			645 => x"ffc10a4d",
			646 => x"000a0a4d",
			647 => x"000c0a4d",
			648 => x"07003010",
			649 => x"09001908",
			650 => x"05002704",
			651 => x"00480a4d",
			652 => x"fff20a4d",
			653 => x"00013a04",
			654 => x"00080a4d",
			655 => x"ffd60a4d",
			656 => x"0e00ac04",
			657 => x"ff950a4d",
			658 => x"00110a4d",
			659 => x"05002518",
			660 => x"01000704",
			661 => x"ffbe0ae9",
			662 => x"00011508",
			663 => x"05002304",
			664 => x"ff8c0ae9",
			665 => x"005e0ae9",
			666 => x"03002608",
			667 => x"03002104",
			668 => x"ffeb0ae9",
			669 => x"00050ae9",
			670 => x"00d10ae9",
			671 => x"0a003118",
			672 => x"09001b0c",
			673 => x"0f00c208",
			674 => x"0f00bb04",
			675 => x"ffe00ae9",
			676 => x"002c0ae9",
			677 => x"ff470ae9",
			678 => x"05002a08",
			679 => x"05002804",
			680 => x"ffee0ae9",
			681 => x"004a0ae9",
			682 => x"ffe30ae9",
			683 => x"00013014",
			684 => x"0d001608",
			685 => x"0f00ca04",
			686 => x"ffd80ae9",
			687 => x"00c60ae9",
			688 => x"01001204",
			689 => x"ffb30ae9",
			690 => x"01001304",
			691 => x"00170ae9",
			692 => x"fff90ae9",
			693 => x"07003008",
			694 => x"0f00c704",
			695 => x"fff60ae9",
			696 => x"002b0ae9",
			697 => x"ff8b0ae9",
			698 => x"0200f704",
			699 => x"fe5b0b3d",
			700 => x"05002e24",
			701 => x"03002a18",
			702 => x"09001808",
			703 => x"01000704",
			704 => x"fe950b3d",
			705 => x"01cd0b3d",
			706 => x"0e009d0c",
			707 => x"00011304",
			708 => x"fd910b3d",
			709 => x"02012704",
			710 => x"ff990b3d",
			711 => x"fe570b3d",
			712 => x"fff00b3d",
			713 => x"00013108",
			714 => x"03002e04",
			715 => x"02890b3d",
			716 => x"01560b3d",
			717 => x"ff3d0b3d",
			718 => x"fe770b3d",
			719 => x"01000a10",
			720 => x"04001408",
			721 => x"08001904",
			722 => x"fff50bc9",
			723 => x"004f0bc9",
			724 => x"05002204",
			725 => x"00180bc9",
			726 => x"ff4d0bc9",
			727 => x"0f00e330",
			728 => x"0d001518",
			729 => x"0001060c",
			730 => x"05002408",
			731 => x"08001d04",
			732 => x"fffb0bc9",
			733 => x"00640bc9",
			734 => x"ff8e0bc9",
			735 => x"00013c08",
			736 => x"0e008a04",
			737 => x"fff60bc9",
			738 => x"01100bc9",
			739 => x"ffe20bc9",
			740 => x"0a00320c",
			741 => x"02011f04",
			742 => x"ff750bc9",
			743 => x"02012c04",
			744 => x"00150bc9",
			745 => x"fff20bc9",
			746 => x"04002108",
			747 => x"0e009204",
			748 => x"fffc0bc9",
			749 => x"004e0bc9",
			750 => x"ffce0bc9",
			751 => x"03002e04",
			752 => x"ff6b0bc9",
			753 => x"00610bc9",
			754 => x"0300260c",
			755 => x"09001808",
			756 => x"07002904",
			757 => x"ffe70c4d",
			758 => x"00580c4d",
			759 => x"fef70c4d",
			760 => x"01000a08",
			761 => x"05002504",
			762 => x"000a0c4d",
			763 => x"ff2b0c4d",
			764 => x"01000b14",
			765 => x"0a003208",
			766 => x"05002904",
			767 => x"01260c4d",
			768 => x"ffc60c4d",
			769 => x"07003204",
			770 => x"ff5d0c4d",
			771 => x"08002004",
			772 => x"00b00c4d",
			773 => x"fff80c4d",
			774 => x"04001708",
			775 => x"01000e04",
			776 => x"00040c4d",
			777 => x"00d00c4d",
			778 => x"02010b08",
			779 => x"02010004",
			780 => x"ff990c4d",
			781 => x"00db0c4d",
			782 => x"0a003204",
			783 => x"ff180c4d",
			784 => x"07003104",
			785 => x"003e0c4d",
			786 => x"ffae0c4d",
			787 => x"0e008a04",
			788 => x"fec50ca1",
			789 => x"03002404",
			790 => x"ff590ca1",
			791 => x"01000804",
			792 => x"fedd0ca1",
			793 => x"0d00150c",
			794 => x"0a003208",
			795 => x"04001a04",
			796 => x"016c0ca1",
			797 => x"00c50ca1",
			798 => x"ffe50ca1",
			799 => x"0e00a70c",
			800 => x"0a003204",
			801 => x"fe9b0ca1",
			802 => x"05003304",
			803 => x"01020ca1",
			804 => x"ff760ca1",
			805 => x"00015204",
			806 => x"01280ca1",
			807 => x"ffe00ca1",
			808 => x"0200f704",
			809 => x"ff380cfd",
			810 => x"02012f24",
			811 => x"07003820",
			812 => x"03002408",
			813 => x"09001804",
			814 => x"003a0cfd",
			815 => x"ff960cfd",
			816 => x"03002f0c",
			817 => x"01000804",
			818 => x"ffcc0cfd",
			819 => x"0a003204",
			820 => x"010d0cfd",
			821 => x"003b0cfd",
			822 => x"07003404",
			823 => x"ff870cfd",
			824 => x"03003304",
			825 => x"00660cfd",
			826 => x"fff00cfd",
			827 => x"ffaa0cfd",
			828 => x"0f00e904",
			829 => x"ff4e0cfd",
			830 => x"00130cfd",
			831 => x"0e009104",
			832 => x"fee60d71",
			833 => x"0e00950c",
			834 => x"0600ad04",
			835 => x"ff950d71",
			836 => x"00013a04",
			837 => x"01220d71",
			838 => x"ffcc0d71",
			839 => x"03002e18",
			840 => x"0e00a514",
			841 => x"0f00d80c",
			842 => x"0e009d08",
			843 => x"0f00d004",
			844 => x"ffc00d71",
			845 => x"ff2e0d71",
			846 => x"00860d71",
			847 => x"09001904",
			848 => x"00c20d71",
			849 => x"ffb20d71",
			850 => x"ff090d71",
			851 => x"0e00a00c",
			852 => x"0f00d108",
			853 => x"0e009b04",
			854 => x"ffbb0d71",
			855 => x"00760d71",
			856 => x"ff3d0d71",
			857 => x"04002304",
			858 => x"01290d71",
			859 => x"fff20d71",
			860 => x"0f00bf04",
			861 => x"fe840dcd",
			862 => x"09001804",
			863 => x"01960dcd",
			864 => x"03002608",
			865 => x"0d001304",
			866 => x"ff490dcd",
			867 => x"fe6a0dcd",
			868 => x"00013010",
			869 => x"0600ae04",
			870 => x"020a0dcd",
			871 => x"03002a04",
			872 => x"ff950dcd",
			873 => x"03002f04",
			874 => x"01640dcd",
			875 => x"ffb80dcd",
			876 => x"01000e0c",
			877 => x"00014908",
			878 => x"02012e04",
			879 => x"ff390dcd",
			880 => x"00f40dcd",
			881 => x"fea90dcd",
			882 => x"fe5f0dcd",
			883 => x"07003338",
			884 => x"09001708",
			885 => x"0a002104",
			886 => x"ffce0e59",
			887 => x"014d0e59",
			888 => x"05002314",
			889 => x"03002a10",
			890 => x"09001804",
			891 => x"001f0e59",
			892 => x"01000908",
			893 => x"01000804",
			894 => x"ffb60e59",
			895 => x"002f0e59",
			896 => x"fe6e0e59",
			897 => x"00850e59",
			898 => x"08001b04",
			899 => x"feb20e59",
			900 => x"0d001308",
			901 => x"05002804",
			902 => x"01790e59",
			903 => x"ff680e59",
			904 => x"0a002f08",
			905 => x"08001c04",
			906 => x"ffe50e59",
			907 => x"fea30e59",
			908 => x"0d001404",
			909 => x"ff130e59",
			910 => x"00ef0e59",
			911 => x"0c001604",
			912 => x"013c0e59",
			913 => x"0d001608",
			914 => x"01000a04",
			915 => x"ff6c0e59",
			916 => x"00e20e59",
			917 => x"febf0e59",
			918 => x"01000804",
			919 => x"fed20ee7",
			920 => x"0d001210",
			921 => x"0500280c",
			922 => x"08001804",
			923 => x"ffc00ee7",
			924 => x"0e007b04",
			925 => x"fff40ee7",
			926 => x"01680ee7",
			927 => x"ff8d0ee7",
			928 => x"07003320",
			929 => x"01000908",
			930 => x"04001c04",
			931 => x"010d0ee7",
			932 => x"ffcf0ee7",
			933 => x"09001b0c",
			934 => x"00012604",
			935 => x"fe770ee7",
			936 => x"00013c04",
			937 => x"00110ee7",
			938 => x"ff380ee7",
			939 => x"0b001508",
			940 => x"03002a04",
			941 => x"ffbe0ee7",
			942 => x"00ea0ee7",
			943 => x"ff1f0ee7",
			944 => x"07003810",
			945 => x"01000a04",
			946 => x"ff040ee7",
			947 => x"0a002d04",
			948 => x"ff2a0ee7",
			949 => x"00013004",
			950 => x"01200ee7",
			951 => x"ff620ee7",
			952 => x"fec20ee7",
			953 => x"0e00920c",
			954 => x"0c001308",
			955 => x"0c001204",
			956 => x"fffb0f21",
			957 => x"00100f21",
			958 => x"ffc50f21",
			959 => x"0e00a40c",
			960 => x"03002f08",
			961 => x"07003604",
			962 => x"006c0f21",
			963 => x"fff60f21",
			964 => x"ffda0f21",
			965 => x"03002e04",
			966 => x"ffca0f21",
			967 => x"002f0f21",
			968 => x"0e009b10",
			969 => x"0c001308",
			970 => x"04001b04",
			971 => x"00280f65",
			972 => x"fffa0f65",
			973 => x"04001404",
			974 => x"00030f65",
			975 => x"ffa50f65",
			976 => x"08001d08",
			977 => x"0600ca04",
			978 => x"00660f65",
			979 => x"00010f65",
			980 => x"0a003204",
			981 => x"ffd30f65",
			982 => x"04002304",
			983 => x"00260f65",
			984 => x"fff50f65",
			985 => x"0e00920c",
			986 => x"0c001308",
			987 => x"0c001204",
			988 => x"fff40fa1",
			989 => x"001f0fa1",
			990 => x"ff8e0fa1",
			991 => x"0b001304",
			992 => x"00790fa1",
			993 => x"02010b04",
			994 => x"00670fa1",
			995 => x"03002e04",
			996 => x"ff6c0fa1",
			997 => x"0e00a104",
			998 => x"ffb80fa1",
			999 => x"00710fa1",
			1000 => x"0e009204",
			1001 => x"ffaf0fdd",
			1002 => x"0500280c",
			1003 => x"00011d04",
			1004 => x"fff20fdd",
			1005 => x"0b001304",
			1006 => x"00950fdd",
			1007 => x"ffff0fdd",
			1008 => x"03002e08",
			1009 => x"0a003404",
			1010 => x"ffb70fdd",
			1011 => x"00000fdd",
			1012 => x"0d001804",
			1013 => x"002b0fdd",
			1014 => x"ffed0fdd",
			1015 => x"0200f704",
			1016 => x"ffa21019",
			1017 => x"03002a14",
			1018 => x"09001808",
			1019 => x"01000704",
			1020 => x"ffde1019",
			1021 => x"004f1019",
			1022 => x"00012408",
			1023 => x"07003304",
			1024 => x"ffd01019",
			1025 => x"00321019",
			1026 => x"ffa21019",
			1027 => x"05002d04",
			1028 => x"009d1019",
			1029 => x"ffd01019",
			1030 => x"00014920",
			1031 => x"0e00910c",
			1032 => x"0c001308",
			1033 => x"0d000f04",
			1034 => x"fff71065",
			1035 => x"003b1065",
			1036 => x"ff681065",
			1037 => x"00011e08",
			1038 => x"0e009504",
			1039 => x"00781065",
			1040 => x"ffb01065",
			1041 => x"0f00e108",
			1042 => x"09001c04",
			1043 => x"00f31065",
			1044 => x"ffdc1065",
			1045 => x"00041065",
			1046 => x"0f00e904",
			1047 => x"ff641065",
			1048 => x"001b1065",
			1049 => x"0c001624",
			1050 => x"03002a14",
			1051 => x"09001808",
			1052 => x"0600a804",
			1053 => x"ffe710b9",
			1054 => x"00d410b9",
			1055 => x"07003308",
			1056 => x"0d001104",
			1057 => x"002810b9",
			1058 => x"ff2010b9",
			1059 => x"005210b9",
			1060 => x"00013108",
			1061 => x"05002e04",
			1062 => x"011e10b9",
			1063 => x"ffe410b9",
			1064 => x"09001a04",
			1065 => x"ffba10b9",
			1066 => x"002e10b9",
			1067 => x"0f00e404",
			1068 => x"ff3c10b9",
			1069 => x"000c10b9",
			1070 => x"0e00920c",
			1071 => x"0c001308",
			1072 => x"0c001204",
			1073 => x"fffa110d",
			1074 => x"000c110d",
			1075 => x"ffc1110d",
			1076 => x"0f00e318",
			1077 => x"0d001408",
			1078 => x"07003204",
			1079 => x"0007110d",
			1080 => x"006b110d",
			1081 => x"0a003208",
			1082 => x"0e009604",
			1083 => x"000c110d",
			1084 => x"ffa3110d",
			1085 => x"04002104",
			1086 => x"0043110d",
			1087 => x"ffef110d",
			1088 => x"0f00ea04",
			1089 => x"ffb7110d",
			1090 => x"001e110d",
			1091 => x"0e009204",
			1092 => x"fe611141",
			1093 => x"07003814",
			1094 => x"0e00a410",
			1095 => x"05002e0c",
			1096 => x"07003308",
			1097 => x"09001904",
			1098 => x"02271141",
			1099 => x"00421141",
			1100 => x"03881141",
			1101 => x"fe691141",
			1102 => x"007a1141",
			1103 => x"fe5d1141",
			1104 => x"0f00ca10",
			1105 => x"0400140c",
			1106 => x"01000908",
			1107 => x"01000804",
			1108 => x"ffe2118d",
			1109 => x"008f118d",
			1110 => x"ff92118d",
			1111 => x"fea9118d",
			1112 => x"09001804",
			1113 => x"00e2118d",
			1114 => x"00014910",
			1115 => x"0700380c",
			1116 => x"07003408",
			1117 => x"05002704",
			1118 => x"ff7c118d",
			1119 => x"00c2118d",
			1120 => x"00d5118d",
			1121 => x"ff1e118d",
			1122 => x"fee0118d",
			1123 => x"0b001310",
			1124 => x"00011704",
			1125 => x"ffc311e9",
			1126 => x"01000704",
			1127 => x"ffdf11e9",
			1128 => x"0e009104",
			1129 => x"000011e9",
			1130 => x"00a211e9",
			1131 => x"02010b0c",
			1132 => x"08001c04",
			1133 => x"ffc511e9",
			1134 => x"0f00bc04",
			1135 => x"ffea11e9",
			1136 => x"006a11e9",
			1137 => x"04001704",
			1138 => x"000311e9",
			1139 => x"01001208",
			1140 => x"0a003604",
			1141 => x"ff9311e9",
			1142 => x"000811e9",
			1143 => x"08002304",
			1144 => x"000e11e9",
			1145 => x"fff711e9",
			1146 => x"0e009104",
			1147 => x"fe611225",
			1148 => x"05002e18",
			1149 => x"0d001510",
			1150 => x"0e00a10c",
			1151 => x"00010604",
			1152 => x"00ed1225",
			1153 => x"02012e04",
			1154 => x"06821225",
			1155 => x"03d81225",
			1156 => x"01d81225",
			1157 => x"0a002f04",
			1158 => x"fdca1225",
			1159 => x"019d1225",
			1160 => x"fe581225",
			1161 => x"03002a20",
			1162 => x"0b00130c",
			1163 => x"00011d04",
			1164 => x"ff381281",
			1165 => x"0e009104",
			1166 => x"ff7c1281",
			1167 => x"00c31281",
			1168 => x"00011210",
			1169 => x"07003304",
			1170 => x"ff851281",
			1171 => x"04001804",
			1172 => x"ffd31281",
			1173 => x"07003504",
			1174 => x"00e01281",
			1175 => x"fff21281",
			1176 => x"fed41281",
			1177 => x"05002e0c",
			1178 => x"00013108",
			1179 => x"0f00c104",
			1180 => x"ffec1281",
			1181 => x"01001281",
			1182 => x"ffde1281",
			1183 => x"ff4f1281",
			1184 => x"0e008a04",
			1185 => x"fe7412d5",
			1186 => x"0d001514",
			1187 => x"03002a0c",
			1188 => x"09001a08",
			1189 => x"05002404",
			1190 => x"00c112d5",
			1191 => x"ffc512d5",
			1192 => x"fe6f12d5",
			1193 => x"00013104",
			1194 => x"01f012d5",
			1195 => x"fefc12d5",
			1196 => x"0e00a008",
			1197 => x"02010b04",
			1198 => x"ffc212d5",
			1199 => x"fdfe12d5",
			1200 => x"03002e04",
			1201 => x"fe6c12d5",
			1202 => x"00014604",
			1203 => x"017012d5",
			1204 => x"ff4312d5",
			1205 => x"04001c28",
			1206 => x"0700331c",
			1207 => x"07002f10",
			1208 => x"03002304",
			1209 => x"fec01339",
			1210 => x"09001908",
			1211 => x"0e008a04",
			1212 => x"ffca1339",
			1213 => x"01941339",
			1214 => x"ff401339",
			1215 => x"05002708",
			1216 => x"00011b04",
			1217 => x"fe301339",
			1218 => x"ff841339",
			1219 => x"00b31339",
			1220 => x"07003808",
			1221 => x"0a002d04",
			1222 => x"ff111339",
			1223 => x"014f1339",
			1224 => x"feb61339",
			1225 => x"0e009b04",
			1226 => x"fe8c1339",
			1227 => x"05003204",
			1228 => x"00761339",
			1229 => x"ff941339",
			1230 => x"0f00bf04",
			1231 => x"fe681385",
			1232 => x"00013018",
			1233 => x"05002304",
			1234 => x"ff0d1385",
			1235 => x"0d001508",
			1236 => x"03002a04",
			1237 => x"011f1385",
			1238 => x"028f1385",
			1239 => x"02011f08",
			1240 => x"0a003204",
			1241 => x"fd8e1385",
			1242 => x"01271385",
			1243 => x"01661385",
			1244 => x"05002204",
			1245 => x"012c1385",
			1246 => x"05002704",
			1247 => x"ffc31385",
			1248 => x"fe5b1385",
			1249 => x"03002a28",
			1250 => x"09001a1c",
			1251 => x"0d001314",
			1252 => x"0c001308",
			1253 => x"00011d04",
			1254 => x"ff6e13f1",
			1255 => x"007b13f1",
			1256 => x"00011e08",
			1257 => x"05002504",
			1258 => x"fff813f1",
			1259 => x"003613f1",
			1260 => x"ff2d13f1",
			1261 => x"03002404",
			1262 => x"ff9813f1",
			1263 => x"00b413f1",
			1264 => x"0d001308",
			1265 => x"04001e04",
			1266 => x"ffd513f1",
			1267 => x"003313f1",
			1268 => x"ff1913f1",
			1269 => x"0200f704",
			1270 => x"ff6213f1",
			1271 => x"05002e08",
			1272 => x"00013104",
			1273 => x"010313f1",
			1274 => x"ffec13f1",
			1275 => x"ff8913f1",
			1276 => x"0600ab04",
			1277 => x"fe691435",
			1278 => x"05002e1c",
			1279 => x"03002a14",
			1280 => x"0b001308",
			1281 => x"0600bf04",
			1282 => x"00061435",
			1283 => x"01631435",
			1284 => x"0f00d708",
			1285 => x"08001c04",
			1286 => x"fe3b1435",
			1287 => x"01d81435",
			1288 => x"fe161435",
			1289 => x"0f00d404",
			1290 => x"02a31435",
			1291 => x"01181435",
			1292 => x"fe761435",
			1293 => x"0b001314",
			1294 => x"00011704",
			1295 => x"ff0014b1",
			1296 => x"05002708",
			1297 => x"01000804",
			1298 => x"000914b1",
			1299 => x"015c14b1",
			1300 => x"0c001404",
			1301 => x"003d14b1",
			1302 => x"ff7d14b1",
			1303 => x"02010b10",
			1304 => x"08001c08",
			1305 => x"00010604",
			1306 => x"ff1014b1",
			1307 => x"008814b1",
			1308 => x"0f00bf04",
			1309 => x"ff7514b1",
			1310 => x"013414b1",
			1311 => x"03002e10",
			1312 => x"04001e08",
			1313 => x"01000904",
			1314 => x"ffd814b1",
			1315 => x"fee714b1",
			1316 => x"0600bf04",
			1317 => x"ff7914b1",
			1318 => x"005b14b1",
			1319 => x"0e00a104",
			1320 => x"ff2814b1",
			1321 => x"00014804",
			1322 => x"00d714b1",
			1323 => x"fff014b1",
			1324 => x"05002518",
			1325 => x"07003210",
			1326 => x"07002f0c",
			1327 => x"0b001308",
			1328 => x"0600ab04",
			1329 => x"fff8152d",
			1330 => x"005c152d",
			1331 => x"ffdd152d",
			1332 => x"ffb7152d",
			1333 => x"03002604",
			1334 => x"ffeb152d",
			1335 => x"0074152d",
			1336 => x"0f00ca0c",
			1337 => x"01000908",
			1338 => x"01000804",
			1339 => x"ffec152d",
			1340 => x"0020152d",
			1341 => x"ff85152d",
			1342 => x"0f00e314",
			1343 => x"0d001508",
			1344 => x"00013d04",
			1345 => x"0099152d",
			1346 => x"ffdc152d",
			1347 => x"0a003204",
			1348 => x"ffc3152d",
			1349 => x"0a003404",
			1350 => x"001d152d",
			1351 => x"ffff152d",
			1352 => x"0a003404",
			1353 => x"ffa6152d",
			1354 => x"0006152d",
			1355 => x"0f00ca10",
			1356 => x"0400140c",
			1357 => x"01000908",
			1358 => x"01000804",
			1359 => x"ffe31589",
			1360 => x"008e1589",
			1361 => x"ff981589",
			1362 => x"feb41589",
			1363 => x"09001804",
			1364 => x"00d71589",
			1365 => x"00014918",
			1366 => x"03002a0c",
			1367 => x"05002504",
			1368 => x"fef11589",
			1369 => x"0d001404",
			1370 => x"00d11589",
			1371 => x"ff391589",
			1372 => x"07003404",
			1373 => x"ffdc1589",
			1374 => x"04002204",
			1375 => x"01301589",
			1376 => x"ffb41589",
			1377 => x"fee91589",
			1378 => x"0e008a04",
			1379 => x"fe7215ed",
			1380 => x"0d001518",
			1381 => x"0001310c",
			1382 => x"00011708",
			1383 => x"09001b04",
			1384 => x"fffd15ed",
			1385 => x"019b15ed",
			1386 => x"017f15ed",
			1387 => x"0b001304",
			1388 => x"00b915ed",
			1389 => x"01000904",
			1390 => x"ff2b15ed",
			1391 => x"fe2e15ed",
			1392 => x"0e00a00c",
			1393 => x"02010b04",
			1394 => x"ff9215ed",
			1395 => x"0a002f04",
			1396 => x"fd7215ed",
			1397 => x"fe9515ed",
			1398 => x"03002e04",
			1399 => x"fe5c15ed",
			1400 => x"04002604",
			1401 => x"018515ed",
			1402 => x"ff3f15ed",
			1403 => x"0e009d28",
			1404 => x"0900180c",
			1405 => x"04001408",
			1406 => x"07002704",
			1407 => x"fffa1671",
			1408 => x"00491671",
			1409 => x"ffee1671",
			1410 => x"0d00110c",
			1411 => x"03002c08",
			1412 => x"03002704",
			1413 => x"fff71671",
			1414 => x"002b1671",
			1415 => x"fff31671",
			1416 => x"03002e08",
			1417 => x"0f00d804",
			1418 => x"ff461671",
			1419 => x"fff31671",
			1420 => x"03002f04",
			1421 => x"002b1671",
			1422 => x"ffdd1671",
			1423 => x"0f00e314",
			1424 => x"0d001504",
			1425 => x"00ac1671",
			1426 => x"0f00d204",
			1427 => x"00261671",
			1428 => x"0f00dd08",
			1429 => x"0a003704",
			1430 => x"ffa11671",
			1431 => x"00041671",
			1432 => x"00121671",
			1433 => x"03002e04",
			1434 => x"ffa61671",
			1435 => x"00451671",
			1436 => x"0600ab04",
			1437 => x"fe6716bd",
			1438 => x"05002e20",
			1439 => x"0001310c",
			1440 => x"02010004",
			1441 => x"005116bd",
			1442 => x"0e009e04",
			1443 => x"036916bd",
			1444 => x"014a16bd",
			1445 => x"04001504",
			1446 => x"01f016bd",
			1447 => x"07003008",
			1448 => x"0b001404",
			1449 => x"013a16bd",
			1450 => x"fe4916bd",
			1451 => x"05002a04",
			1452 => x"fd9016bd",
			1453 => x"fe8816bd",
			1454 => x"fe6a16bd",
			1455 => x"07003320",
			1456 => x"0d00120c",
			1457 => x"01000804",
			1458 => x"ffb31739",
			1459 => x"07002904",
			1460 => x"fff51739",
			1461 => x"00961739",
			1462 => x"09001804",
			1463 => x"00291739",
			1464 => x"04001a04",
			1465 => x"ff591739",
			1466 => x"04001c04",
			1467 => x"00331739",
			1468 => x"05002504",
			1469 => x"00041739",
			1470 => x"ffcd1739",
			1471 => x"0001301c",
			1472 => x"0700350c",
			1473 => x"05002e08",
			1474 => x"0a002d04",
			1475 => x"fff81739",
			1476 => x"00c71739",
			1477 => x"ffec1739",
			1478 => x"03002e04",
			1479 => x"ffc41739",
			1480 => x"08001d04",
			1481 => x"fff81739",
			1482 => x"04002504",
			1483 => x"002c1739",
			1484 => x"fffb1739",
			1485 => x"ffc11739",
			1486 => x"0200f704",
			1487 => x"fe7a179d",
			1488 => x"0001301c",
			1489 => x"0d001510",
			1490 => x"03002404",
			1491 => x"feb2179d",
			1492 => x"05002e08",
			1493 => x"0600ab04",
			1494 => x"ff8f179d",
			1495 => x"01aa179d",
			1496 => x"ff38179d",
			1497 => x"0a003204",
			1498 => x"fe64179d",
			1499 => x"04002304",
			1500 => x"0136179d",
			1501 => x"ff41179d",
			1502 => x"05002304",
			1503 => x"00c2179d",
			1504 => x"0d001408",
			1505 => x"03002604",
			1506 => x"ffbd179d",
			1507 => x"fe81179d",
			1508 => x"05002a04",
			1509 => x"00d0179d",
			1510 => x"fef2179d",
			1511 => x"0f00bf04",
			1512 => x"fe6717f9",
			1513 => x"00013014",
			1514 => x"05002304",
			1515 => x"feea17f9",
			1516 => x"03002f0c",
			1517 => x"0600ad04",
			1518 => x"06ae17f9",
			1519 => x"07003704",
			1520 => x"01fd17f9",
			1521 => x"fe7c17f9",
			1522 => x"ff1117f9",
			1523 => x"05002204",
			1524 => x"015a17f9",
			1525 => x"0700300c",
			1526 => x"08001b04",
			1527 => x"fe5f17f9",
			1528 => x"0b001404",
			1529 => x"018317f9",
			1530 => x"fee417f9",
			1531 => x"0e00ac04",
			1532 => x"fe2817f9",
			1533 => x"009717f9",
			1534 => x"03002a30",
			1535 => x"0900180c",
			1536 => x"01000704",
			1537 => x"ff6d1895",
			1538 => x"0600a604",
			1539 => x"ffec1895",
			1540 => x"01301895",
			1541 => x"0200ee10",
			1542 => x"09001a0c",
			1543 => x"04001908",
			1544 => x"07002b04",
			1545 => x"fff81895",
			1546 => x"00ff1895",
			1547 => x"ffea1895",
			1548 => x"ff871895",
			1549 => x"0b001308",
			1550 => x"0d001204",
			1551 => x"00f81895",
			1552 => x"ff7c1895",
			1553 => x"08001f04",
			1554 => x"fe931895",
			1555 => x"00012604",
			1556 => x"00a91895",
			1557 => x"ffd31895",
			1558 => x"03002f14",
			1559 => x"00013108",
			1560 => x"0f00c104",
			1561 => x"ffbe1895",
			1562 => x"016b1895",
			1563 => x"01000e08",
			1564 => x"0f00d004",
			1565 => x"ffad1895",
			1566 => x"00941895",
			1567 => x"ff2e1895",
			1568 => x"0e00a004",
			1569 => x"fed71895",
			1570 => x"00014804",
			1571 => x"00ce1895",
			1572 => x"ffed1895",
			1573 => x"03002a30",
			1574 => x"0900180c",
			1575 => x"01000704",
			1576 => x"ff711931",
			1577 => x"0600a604",
			1578 => x"ffed1931",
			1579 => x"01261931",
			1580 => x"0500230c",
			1581 => x"01000908",
			1582 => x"01000804",
			1583 => x"ffe31931",
			1584 => x"001f1931",
			1585 => x"febd1931",
			1586 => x"00012110",
			1587 => x"0d00140c",
			1588 => x"03002604",
			1589 => x"ff421931",
			1590 => x"04001d04",
			1591 => x"01541931",
			1592 => x"ff791931",
			1593 => x"ff211931",
			1594 => x"0c001404",
			1595 => x"00071931",
			1596 => x"febe1931",
			1597 => x"03002f14",
			1598 => x"00013108",
			1599 => x"0f00c104",
			1600 => x"ffc11931",
			1601 => x"01631931",
			1602 => x"01000e08",
			1603 => x"0f00d004",
			1604 => x"ffb21931",
			1605 => x"008d1931",
			1606 => x"ff3a1931",
			1607 => x"0e00a004",
			1608 => x"fee31931",
			1609 => x"00014804",
			1610 => x"00c61931",
			1611 => x"ffee1931",
			1612 => x"01000a0c",
			1613 => x"05002208",
			1614 => x"03002304",
			1615 => x"ffb919bd",
			1616 => x"009419bd",
			1617 => x"ff2819bd",
			1618 => x"01000b18",
			1619 => x"04001508",
			1620 => x"04001004",
			1621 => x"006d19bd",
			1622 => x"ff8619bd",
			1623 => x"04001b04",
			1624 => x"012819bd",
			1625 => x"07003204",
			1626 => x"ffcb19bd",
			1627 => x"08001f04",
			1628 => x"002d19bd",
			1629 => x"000019bd",
			1630 => x"0400160c",
			1631 => x"0d001304",
			1632 => x"ffcb19bd",
			1633 => x"0b001504",
			1634 => x"00b819bd",
			1635 => x"ffd719bd",
			1636 => x"0500290c",
			1637 => x"05002508",
			1638 => x"05002304",
			1639 => x"ffe119bd",
			1640 => x"002b19bd",
			1641 => x"ff2619bd",
			1642 => x"00011d08",
			1643 => x"0e008c04",
			1644 => x"ffd919bd",
			1645 => x"00df19bd",
			1646 => x"ff5419bd",
			1647 => x"0e008a04",
			1648 => x"fead1a01",
			1649 => x"0700381c",
			1650 => x"03002404",
			1651 => x"ff271a01",
			1652 => x"01000804",
			1653 => x"febb1a01",
			1654 => x"07002f04",
			1655 => x"01791a01",
			1656 => x"00013008",
			1657 => x"00011f04",
			1658 => x"002f1a01",
			1659 => x"01531a01",
			1660 => x"01000e04",
			1661 => x"ffdd1a01",
			1662 => x"febf1a01",
			1663 => x"feaa1a01",
			1664 => x"0f00bf04",
			1665 => x"fe881a55",
			1666 => x"09001804",
			1667 => x"01901a55",
			1668 => x"03002608",
			1669 => x"0d001304",
			1670 => x"ff611a55",
			1671 => x"fe751a55",
			1672 => x"00013010",
			1673 => x"0600ae04",
			1674 => x"01de1a55",
			1675 => x"0c001504",
			1676 => x"ffac1a55",
			1677 => x"00011d04",
			1678 => x"01901a55",
			1679 => x"ffd71a55",
			1680 => x"01000e08",
			1681 => x"0b001404",
			1682 => x"005d1a55",
			1683 => x"feb21a55",
			1684 => x"fe6f1a55",
			1685 => x"01000a14",
			1686 => x"04001408",
			1687 => x"02011204",
			1688 => x"ffce1ae9",
			1689 => x"00861ae9",
			1690 => x"05002208",
			1691 => x"05001f04",
			1692 => x"00071ae9",
			1693 => x"fff71ae9",
			1694 => x"ff1e1ae9",
			1695 => x"0d001208",
			1696 => x"07002a04",
			1697 => x"ffdc1ae9",
			1698 => x"00f51ae9",
			1699 => x"07003318",
			1700 => x"09001b0c",
			1701 => x"07002f08",
			1702 => x"0c001304",
			1703 => x"00861ae9",
			1704 => x"ffb61ae9",
			1705 => x"ff2f1ae9",
			1706 => x"04001c08",
			1707 => x"07003004",
			1708 => x"ffee1ae9",
			1709 => x"00961ae9",
			1710 => x"ffbf1ae9",
			1711 => x"07003814",
			1712 => x"0d001608",
			1713 => x"00012a04",
			1714 => x"010b1ae9",
			1715 => x"000f1ae9",
			1716 => x"01001204",
			1717 => x"ff851ae9",
			1718 => x"05002f04",
			1719 => x"002e1ae9",
			1720 => x"fff11ae9",
			1721 => x"ff791ae9",
			1722 => x"0e008a04",
			1723 => x"fe6d1b45",
			1724 => x"0d001204",
			1725 => x"01841b45",
			1726 => x"00014920",
			1727 => x"0d001614",
			1728 => x"07003208",
			1729 => x"00013304",
			1730 => x"ff181b45",
			1731 => x"014b1b45",
			1732 => x"01000a04",
			1733 => x"ffb81b45",
			1734 => x"00012504",
			1735 => x"02711b45",
			1736 => x"007a1b45",
			1737 => x"0a003108",
			1738 => x"0f00d004",
			1739 => x"fefd1b45",
			1740 => x"00f21b45",
			1741 => x"fe4f1b45",
			1742 => x"0600cb04",
			1743 => x"fe551b45",
			1744 => x"00061b45",
			1745 => x"0f00bf04",
			1746 => x"fe931ba9",
			1747 => x"01000808",
			1748 => x"03002404",
			1749 => x"009e1ba9",
			1750 => x"fe911ba9",
			1751 => x"03002408",
			1752 => x"07002e04",
			1753 => x"ffa61ba9",
			1754 => x"fe8f1ba9",
			1755 => x"0d001510",
			1756 => x"0a00320c",
			1757 => x"04001d08",
			1758 => x"0f00df04",
			1759 => x"01ad1ba9",
			1760 => x"00b61ba9",
			1761 => x"febc1ba9",
			1762 => x"ffff1ba9",
			1763 => x"0f00e60c",
			1764 => x"0a003204",
			1765 => x"fe5d1ba9",
			1766 => x"04002104",
			1767 => x"01111ba9",
			1768 => x"ff111ba9",
			1769 => x"01221ba9",
			1770 => x"01000808",
			1771 => x"07003304",
			1772 => x"ff831c2d",
			1773 => x"fffd1c2d",
			1774 => x"0200fb10",
			1775 => x"05002408",
			1776 => x"05002204",
			1777 => x"ffe81c2d",
			1778 => x"00621c2d",
			1779 => x"01000904",
			1780 => x"002d1c2d",
			1781 => x"ff5c1c2d",
			1782 => x"0f00e324",
			1783 => x"0d001510",
			1784 => x"00013c0c",
			1785 => x"05002e08",
			1786 => x"03002404",
			1787 => x"fff31c2d",
			1788 => x"010b1c2d",
			1789 => x"ffef1c2d",
			1790 => x"ffda1c2d",
			1791 => x"02010b08",
			1792 => x"00010f04",
			1793 => x"fffa1c2d",
			1794 => x"002f1c2d",
			1795 => x"0f00de08",
			1796 => x"01001204",
			1797 => x"ff7b1c2d",
			1798 => x"00071c2d",
			1799 => x"00151c2d",
			1800 => x"03002e04",
			1801 => x"ff921c2d",
			1802 => x"005e1c2d",
			1803 => x"01000a18",
			1804 => x"0400140c",
			1805 => x"08001d08",
			1806 => x"07002904",
			1807 => x"fff41ce9",
			1808 => x"00911ce9",
			1809 => x"ffe41ce9",
			1810 => x"05002208",
			1811 => x"05002104",
			1812 => x"fffc1ce9",
			1813 => x"00001ce9",
			1814 => x"ff2d1ce9",
			1815 => x"01000b18",
			1816 => x"04001508",
			1817 => x"04001004",
			1818 => x"006b1ce9",
			1819 => x"ffbc1ce9",
			1820 => x"04001b04",
			1821 => x"01001ce9",
			1822 => x"07003204",
			1823 => x"ffdf1ce9",
			1824 => x"08002004",
			1825 => x"00151ce9",
			1826 => x"fffb1ce9",
			1827 => x"0700341c",
			1828 => x"05002914",
			1829 => x"04001408",
			1830 => x"07002b04",
			1831 => x"fff81ce9",
			1832 => x"00421ce9",
			1833 => x"05002508",
			1834 => x"05002304",
			1835 => x"ffe11ce9",
			1836 => x"00271ce9",
			1837 => x"ff3a1ce9",
			1838 => x"04001e04",
			1839 => x"00581ce9",
			1840 => x"ffdc1ce9",
			1841 => x"07003610",
			1842 => x"0d001804",
			1843 => x"00b71ce9",
			1844 => x"03002e04",
			1845 => x"ffad1ce9",
			1846 => x"03003304",
			1847 => x"00541ce9",
			1848 => x"fffb1ce9",
			1849 => x"ff8f1ce9",
			1850 => x"0900180c",
			1851 => x"01000704",
			1852 => x"ff691d67",
			1853 => x"0f00c604",
			1854 => x"ffbe1d67",
			1855 => x"014a1d67",
			1856 => x"02012f30",
			1857 => x"0d001208",
			1858 => x"01000a04",
			1859 => x"ff7c1d67",
			1860 => x"01401d67",
			1861 => x"07003214",
			1862 => x"0001330c",
			1863 => x"03002e04",
			1864 => x"fe8e1d67",
			1865 => x"0b001504",
			1866 => x"00e71d67",
			1867 => x"ff891d67",
			1868 => x"0e008604",
			1869 => x"fff51d67",
			1870 => x"00d61d67",
			1871 => x"0d001404",
			1872 => x"00dd1d67",
			1873 => x"0a003208",
			1874 => x"02011f04",
			1875 => x"fe8d1d67",
			1876 => x"01011d67",
			1877 => x"04002204",
			1878 => x"013d1d67",
			1879 => x"ff641d67",
			1880 => x"feb91d67",
			1881 => x"0600bc10",
			1882 => x"0e009104",
			1883 => x"c00d1da1",
			1884 => x"09001b04",
			1885 => x"e1d41da1",
			1886 => x"09001d04",
			1887 => x"c87d1da1",
			1888 => x"c0121da1",
			1889 => x"09001c08",
			1890 => x"03002a04",
			1891 => x"e7a71da1",
			1892 => x"fd7b1da1",
			1893 => x"02013204",
			1894 => x"c49b1da1",
			1895 => x"c0171da1",
			1896 => x"0e009204",
			1897 => x"fe621dcd",
			1898 => x"0c001710",
			1899 => x"0e00a40c",
			1900 => x"07003308",
			1901 => x"0f00dc04",
			1902 => x"00db1dcd",
			1903 => x"020d1dcd",
			1904 => x"02ea1dcd",
			1905 => x"004b1dcd",
			1906 => x"fe6c1dcd",
			1907 => x"0e00920c",
			1908 => x"0d001008",
			1909 => x"0d000f04",
			1910 => x"fffa1e11",
			1911 => x"000e1e11",
			1912 => x"ffbc1e11",
			1913 => x"0e009e08",
			1914 => x"05002a04",
			1915 => x"00741e11",
			1916 => x"ffe91e11",
			1917 => x"07003404",
			1918 => x"ffc71e11",
			1919 => x"03002a04",
			1920 => x"ffeb1e11",
			1921 => x"05002f04",
			1922 => x"005b1e11",
			1923 => x"fff21e11",
			1924 => x"0e00920c",
			1925 => x"0d001008",
			1926 => x"03002904",
			1927 => x"fff01e5d",
			1928 => x"00331e5d",
			1929 => x"ff611e5d",
			1930 => x"0700330c",
			1931 => x"07002f04",
			1932 => x"00801e5d",
			1933 => x"05002704",
			1934 => x"ff861e5d",
			1935 => x"004c1e5d",
			1936 => x"0c001604",
			1937 => x"00b41e5d",
			1938 => x"04001e04",
			1939 => x"ffa51e5d",
			1940 => x"04002204",
			1941 => x"00361e5d",
			1942 => x"ffe71e5d",
			1943 => x"01000a14",
			1944 => x"0400140c",
			1945 => x"08001d08",
			1946 => x"07002904",
			1947 => x"fffc1eb1",
			1948 => x"00371eb1",
			1949 => x"fff71eb1",
			1950 => x"05001f04",
			1951 => x"00031eb1",
			1952 => x"ffa71eb1",
			1953 => x"03002608",
			1954 => x"0c001304",
			1955 => x"00201eb1",
			1956 => x"ffc41eb1",
			1957 => x"05002e0c",
			1958 => x"0e00a408",
			1959 => x"0f00bf04",
			1960 => x"fff11eb1",
			1961 => x"008d1eb1",
			1962 => x"fffe1eb1",
			1963 => x"ffde1eb1",
			1964 => x"04001710",
			1965 => x"02011308",
			1966 => x"03002a04",
			1967 => x"ffb71f0d",
			1968 => x"00151f0d",
			1969 => x"03002304",
			1970 => x"ffe81f0d",
			1971 => x"00971f0d",
			1972 => x"02010b10",
			1973 => x"07003104",
			1974 => x"ffde1f0d",
			1975 => x"0a002d04",
			1976 => x"fff01f0d",
			1977 => x"04002104",
			1978 => x"00731f0d",
			1979 => x"fff71f0d",
			1980 => x"0b001308",
			1981 => x"0a002f04",
			1982 => x"ffea1f0d",
			1983 => x"00201f0d",
			1984 => x"05002504",
			1985 => x"00011f0d",
			1986 => x"ff7b1f0d",
			1987 => x"00013018",
			1988 => x"0f00bf04",
			1989 => x"ff8e1f61",
			1990 => x"05002304",
			1991 => x"ffb61f61",
			1992 => x"0d001508",
			1993 => x"0f00ca04",
			1994 => x"00371f61",
			1995 => x"00d71f61",
			1996 => x"0a003204",
			1997 => x"ffb91f61",
			1998 => x"001a1f61",
			1999 => x"0700300c",
			2000 => x"0b001408",
			2001 => x"0600bb04",
			2002 => x"ffdd1f61",
			2003 => x"00a31f61",
			2004 => x"ffa41f61",
			2005 => x"0e00ac04",
			2006 => x"ff321f61",
			2007 => x"002d1f61",
			2008 => x"0f00ca14",
			2009 => x"05002508",
			2010 => x"03002704",
			2011 => x"ffee1fbd",
			2012 => x"00491fbd",
			2013 => x"03002e04",
			2014 => x"ff791fbd",
			2015 => x"03003104",
			2016 => x"00191fbd",
			2017 => x"ffe21fbd",
			2018 => x"0f00e314",
			2019 => x"02012f10",
			2020 => x"0d001508",
			2021 => x"05002504",
			2022 => x"00041fbd",
			2023 => x"00b11fbd",
			2024 => x"03002e04",
			2025 => x"ffd21fbd",
			2026 => x"00001fbd",
			2027 => x"ffc11fbd",
			2028 => x"03002e04",
			2029 => x"ffa21fbd",
			2030 => x"00311fbd",
			2031 => x"0e009104",
			2032 => x"fe731ff9",
			2033 => x"07003818",
			2034 => x"0700330c",
			2035 => x"0b001304",
			2036 => x"00aa1ff9",
			2037 => x"05002704",
			2038 => x"fed21ff9",
			2039 => x"00b81ff9",
			2040 => x"0d001404",
			2041 => x"01aa1ff9",
			2042 => x"0a003204",
			2043 => x"ff7f1ff9",
			2044 => x"018b1ff9",
			2045 => x"fe911ff9",
			2046 => x"0e00920c",
			2047 => x"0d001008",
			2048 => x"01000904",
			2049 => x"ffb2204d",
			2050 => x"00ea204d",
			2051 => x"fea4204d",
			2052 => x"0f00e318",
			2053 => x"08001c08",
			2054 => x"0f00d804",
			2055 => x"ff15204d",
			2056 => x"0117204d",
			2057 => x"0d001604",
			2058 => x"0134204d",
			2059 => x"01001204",
			2060 => x"fef9204d",
			2061 => x"01001404",
			2062 => x"0076204d",
			2063 => x"ffaf204d",
			2064 => x"05002504",
			2065 => x"002e204d",
			2066 => x"feab204d",
			2067 => x"0f00d924",
			2068 => x"07003214",
			2069 => x"0d00140c",
			2070 => x"0d001108",
			2071 => x"0d000f04",
			2072 => x"fffa20b1",
			2073 => x"000e20b1",
			2074 => x"ff9e20b1",
			2075 => x"09001c04",
			2076 => x"001920b1",
			2077 => x"fff620b1",
			2078 => x"0d001404",
			2079 => x"004520b1",
			2080 => x"0a003204",
			2081 => x"ffb320b1",
			2082 => x"04002004",
			2083 => x"002f20b1",
			2084 => x"ffed20b1",
			2085 => x"02014708",
			2086 => x"0600ca04",
			2087 => x"006320b1",
			2088 => x"000520b1",
			2089 => x"0600cb04",
			2090 => x"ffd420b1",
			2091 => x"000420b1",
			2092 => x"0e009104",
			2093 => x"fe6120ed",
			2094 => x"05002e18",
			2095 => x"0d001510",
			2096 => x"0e00a10c",
			2097 => x"00010604",
			2098 => x"00dc20ed",
			2099 => x"02012e04",
			2100 => x"050820ed",
			2101 => x"031020ed",
			2102 => x"018c20ed",
			2103 => x"0a002f04",
			2104 => x"fdce20ed",
			2105 => x"016720ed",
			2106 => x"fe5b20ed",
			2107 => x"0e009d28",
			2108 => x"0900180c",
			2109 => x"04001408",
			2110 => x"07002704",
			2111 => x"fffa2159",
			2112 => x"00472159",
			2113 => x"ffee2159",
			2114 => x"0d00110c",
			2115 => x"03002c08",
			2116 => x"03002704",
			2117 => x"fff72159",
			2118 => x"002b2159",
			2119 => x"fff32159",
			2120 => x"03002e08",
			2121 => x"0f00d804",
			2122 => x"ff502159",
			2123 => x"fff52159",
			2124 => x"03002f04",
			2125 => x"002a2159",
			2126 => x"ffde2159",
			2127 => x"0f00e308",
			2128 => x"0d001704",
			2129 => x"00962159",
			2130 => x"ffc52159",
			2131 => x"0600ce04",
			2132 => x"ff9f2159",
			2133 => x"00372159",
			2134 => x"0c001624",
			2135 => x"0700321c",
			2136 => x"09001808",
			2137 => x"0e008404",
			2138 => x"ffe621ad",
			2139 => x"00cf21ad",
			2140 => x"0d001108",
			2141 => x"02011304",
			2142 => x"007821ad",
			2143 => x"ffef21ad",
			2144 => x"01000908",
			2145 => x"03002a04",
			2146 => x"ffd621ad",
			2147 => x"002c21ad",
			2148 => x"ff3421ad",
			2149 => x"00012604",
			2150 => x"00f121ad",
			2151 => x"001621ad",
			2152 => x"0f00e404",
			2153 => x"ff4621ad",
			2154 => x"000b21ad",
			2155 => x"0e00920c",
			2156 => x"0c001308",
			2157 => x"0c001204",
			2158 => x"ffe82209",
			2159 => x"00492209",
			2160 => x"ff522209",
			2161 => x"0e00a41c",
			2162 => x"03002f14",
			2163 => x"0200f704",
			2164 => x"ffdd2209",
			2165 => x"00014908",
			2166 => x"07003604",
			2167 => x"00d12209",
			2168 => x"ffea2209",
			2169 => x"00015504",
			2170 => x"ffce2209",
			2171 => x"00142209",
			2172 => x"0e00a004",
			2173 => x"ff7c2209",
			2174 => x"001f2209",
			2175 => x"03002e04",
			2176 => x"ff9d2209",
			2177 => x"00592209",
			2178 => x"0e008a04",
			2179 => x"fe762255",
			2180 => x"00013018",
			2181 => x"05002304",
			2182 => x"ff132255",
			2183 => x"0d001508",
			2184 => x"03002a04",
			2185 => x"00d32255",
			2186 => x"01d72255",
			2187 => x"0a003204",
			2188 => x"fee42255",
			2189 => x"0e009604",
			2190 => x"ff412255",
			2191 => x"01192255",
			2192 => x"07003008",
			2193 => x"09001904",
			2194 => x"01432255",
			2195 => x"fecb2255",
			2196 => x"fe492255",
			2197 => x"03002a28",
			2198 => x"09001a1c",
			2199 => x"0d001314",
			2200 => x"05002208",
			2201 => x"0a002504",
			2202 => x"fff022c1",
			2203 => x"006422c1",
			2204 => x"05002504",
			2205 => x"ff4522c1",
			2206 => x"00013504",
			2207 => x"003222c1",
			2208 => x"ffac22c1",
			2209 => x"03002404",
			2210 => x"ff9e22c1",
			2211 => x"00a822c1",
			2212 => x"0d001308",
			2213 => x"04001e04",
			2214 => x"ffd622c1",
			2215 => x"003122c1",
			2216 => x"ff2222c1",
			2217 => x"0200f704",
			2218 => x"ff6922c1",
			2219 => x"05002e08",
			2220 => x"00013104",
			2221 => x"00fa22c1",
			2222 => x"ffef22c1",
			2223 => x"ff8f22c1",
			2224 => x"0600b620",
			2225 => x"0500250c",
			2226 => x"03002708",
			2227 => x"0c001304",
			2228 => x"00042345",
			2229 => x"ffe52345",
			2230 => x"00422345",
			2231 => x"01000908",
			2232 => x"01000804",
			2233 => x"ffea2345",
			2234 => x"00202345",
			2235 => x"0f00cb04",
			2236 => x"ff802345",
			2237 => x"0f00cd04",
			2238 => x"000c2345",
			2239 => x"fff82345",
			2240 => x"0e00a418",
			2241 => x"0001490c",
			2242 => x"03002f08",
			2243 => x"07003604",
			2244 => x"00962345",
			2245 => x"fff82345",
			2246 => x"ffda2345",
			2247 => x"0e009b04",
			2248 => x"ffd22345",
			2249 => x"0e00a004",
			2250 => x"00142345",
			2251 => x"ffea2345",
			2252 => x"03002c04",
			2253 => x"ff902345",
			2254 => x"0e00a604",
			2255 => x"ffe32345",
			2256 => x"005a2345",
			2257 => x"0e008a04",
			2258 => x"fe6f2399",
			2259 => x"00013018",
			2260 => x"0e008d04",
			2261 => x"03622399",
			2262 => x"0f00cb0c",
			2263 => x"0f00c208",
			2264 => x"0f00bf04",
			2265 => x"feac2399",
			2266 => x"02432399",
			2267 => x"fe4b2399",
			2268 => x"03002a04",
			2269 => x"008d2399",
			2270 => x"01b92399",
			2271 => x"07003008",
			2272 => x"0e009804",
			2273 => x"fe712399",
			2274 => x"016b2399",
			2275 => x"0e00ab04",
			2276 => x"fe2c2399",
			2277 => x"00102399",
			2278 => x"0600ab04",
			2279 => x"fe6323dd",
			2280 => x"05002e1c",
			2281 => x"0b001308",
			2282 => x"07002f04",
			2283 => x"03e823dd",
			2284 => x"019d23dd",
			2285 => x"03002604",
			2286 => x"fe1023dd",
			2287 => x"00013108",
			2288 => x"02010b04",
			2289 => x"03b723dd",
			2290 => x"01c623dd",
			2291 => x"0e009304",
			2292 => x"fe5523dd",
			2293 => x"fffd23dd",
			2294 => x"fe5e23dd",
			2295 => x"03002a28",
			2296 => x"09001708",
			2297 => x"08001804",
			2298 => x"fffb2449",
			2299 => x"00442449",
			2300 => x"0200ee08",
			2301 => x"0b001404",
			2302 => x"00472449",
			2303 => x"fff12449",
			2304 => x"0b00130c",
			2305 => x"05002504",
			2306 => x"ffbc2449",
			2307 => x"0a002d04",
			2308 => x"fffb2449",
			2309 => x"003f2449",
			2310 => x"08001f04",
			2311 => x"ff622449",
			2312 => x"08002204",
			2313 => x"00222449",
			2314 => x"fffc2449",
			2315 => x"0200f704",
			2316 => x"ffb02449",
			2317 => x"05002e08",
			2318 => x"0e008a04",
			2319 => x"fffb2449",
			2320 => x"00cf2449",
			2321 => x"ffce2449",
			2322 => x"0b001314",
			2323 => x"00011704",
			2324 => x"ff0c24cd",
			2325 => x"05002708",
			2326 => x"01000804",
			2327 => x"000e24cd",
			2328 => x"015424cd",
			2329 => x"0a002f04",
			2330 => x"ff8224cd",
			2331 => x"003724cd",
			2332 => x"02010b14",
			2333 => x"0200f70c",
			2334 => x"05002408",
			2335 => x"03002704",
			2336 => x"ffc424cd",
			2337 => x"00e424cd",
			2338 => x"ff0524cd",
			2339 => x"04002104",
			2340 => x"012624cd",
			2341 => x"ffcf24cd",
			2342 => x"03002e10",
			2343 => x"0e00a50c",
			2344 => x"0e009b04",
			2345 => x"ff1424cd",
			2346 => x"01001904",
			2347 => x"00a024cd",
			2348 => x"fffa24cd",
			2349 => x"fedf24cd",
			2350 => x"0e00a104",
			2351 => x"ff3324cd",
			2352 => x"00014804",
			2353 => x"00cf24cd",
			2354 => x"fff024cd",
			2355 => x"0c001628",
			2356 => x"07003320",
			2357 => x"08001d18",
			2358 => x"02010a08",
			2359 => x"03002a04",
			2360 => x"ff722541",
			2361 => x"002d2541",
			2362 => x"01000704",
			2363 => x"ffb02541",
			2364 => x"08001804",
			2365 => x"ffe62541",
			2366 => x"0b001304",
			2367 => x"00b22541",
			2368 => x"00132541",
			2369 => x"04002004",
			2370 => x"ff6c2541",
			2371 => x"00072541",
			2372 => x"04001604",
			2373 => x"00202541",
			2374 => x"00992541",
			2375 => x"03002e04",
			2376 => x"ff8d2541",
			2377 => x"03003108",
			2378 => x"0e009404",
			2379 => x"fff72541",
			2380 => x"002d2541",
			2381 => x"0600c304",
			2382 => x"ffd42541",
			2383 => x"00012541",
			2384 => x"0f00bf04",
			2385 => x"fe65259d",
			2386 => x"00013018",
			2387 => x"03002604",
			2388 => x"fef6259d",
			2389 => x"0d001508",
			2390 => x"00012304",
			2391 => x"0307259d",
			2392 => x"01a7259d",
			2393 => x"03002e04",
			2394 => x"fe39259d",
			2395 => x"00012a04",
			2396 => x"0009259d",
			2397 => x"0193259d",
			2398 => x"04001504",
			2399 => x"01cd259d",
			2400 => x"07003008",
			2401 => x"0c001404",
			2402 => x"012e259d",
			2403 => x"fe59259d",
			2404 => x"05002a04",
			2405 => x"fdb4259d",
			2406 => x"fe69259d",
			2407 => x"05002514",
			2408 => x"03002608",
			2409 => x"0c001304",
			2410 => x"003a2621",
			2411 => x"ffaf2621",
			2412 => x"00011508",
			2413 => x"01000b04",
			2414 => x"00062621",
			2415 => x"fff72621",
			2416 => x"00972621",
			2417 => x"0f00e328",
			2418 => x"0f00ca14",
			2419 => x"01000908",
			2420 => x"01000804",
			2421 => x"fff12621",
			2422 => x"00242621",
			2423 => x"03002e04",
			2424 => x"ff912621",
			2425 => x"0a003204",
			2426 => x"001d2621",
			2427 => x"ffe72621",
			2428 => x"0d001508",
			2429 => x"00013d04",
			2430 => x"00982621",
			2431 => x"ffe02621",
			2432 => x"0a003204",
			2433 => x"ffbc2621",
			2434 => x"04002104",
			2435 => x"002c2621",
			2436 => x"ffee2621",
			2437 => x"0a003404",
			2438 => x"ff9c2621",
			2439 => x"00062621",
			2440 => x"0e00920c",
			2441 => x"0d001008",
			2442 => x"03002904",
			2443 => x"fff12685",
			2444 => x"00332685",
			2445 => x"ff672685",
			2446 => x"03002604",
			2447 => x"ffda2685",
			2448 => x"03002f18",
			2449 => x"0e00a410",
			2450 => x"04001d04",
			2451 => x"00ce2685",
			2452 => x"08001f04",
			2453 => x"ffb52685",
			2454 => x"07003b04",
			2455 => x"00422685",
			2456 => x"fffc2685",
			2457 => x"0d001604",
			2458 => x"00172685",
			2459 => x"ffbb2685",
			2460 => x"0e00a004",
			2461 => x"ff832685",
			2462 => x"00014604",
			2463 => x"00532685",
			2464 => x"fffb2685",
			2465 => x"01000b28",
			2466 => x"0100080c",
			2467 => x"04001004",
			2468 => x"00252709",
			2469 => x"07003304",
			2470 => x"ff8d2709",
			2471 => x"fffe2709",
			2472 => x"08001804",
			2473 => x"ffcb2709",
			2474 => x"0a00320c",
			2475 => x"0f00bf04",
			2476 => x"ffde2709",
			2477 => x"03002604",
			2478 => x"fffb2709",
			2479 => x"00ec2709",
			2480 => x"07003204",
			2481 => x"ffa52709",
			2482 => x"08001f04",
			2483 => x"00502709",
			2484 => x"00002709",
			2485 => x"0a003214",
			2486 => x"09001804",
			2487 => x"00332709",
			2488 => x"09001c04",
			2489 => x"ff422709",
			2490 => x"0b001608",
			2491 => x"08001f04",
			2492 => x"fff32709",
			2493 => x"002a2709",
			2494 => x"ffeb2709",
			2495 => x"05002f04",
			2496 => x"00572709",
			2497 => x"ffd22709",
			2498 => x"00013030",
			2499 => x"07003010",
			2500 => x"0d001108",
			2501 => x"07002b04",
			2502 => x"fffb2795",
			2503 => x"001a2795",
			2504 => x"09001804",
			2505 => x"000c2795",
			2506 => x"ffb22795",
			2507 => x"03002604",
			2508 => x"ffd32795",
			2509 => x"0d00150c",
			2510 => x"01000a04",
			2511 => x"fff02795",
			2512 => x"0f00bf04",
			2513 => x"ffed2795",
			2514 => x"00a62795",
			2515 => x"08001d04",
			2516 => x"00202795",
			2517 => x"01001208",
			2518 => x"0a003604",
			2519 => x"ffbf2795",
			2520 => x"000a2795",
			2521 => x"000c2795",
			2522 => x"07003010",
			2523 => x"09001908",
			2524 => x"05002704",
			2525 => x"004a2795",
			2526 => x"fff22795",
			2527 => x"00013a04",
			2528 => x"00082795",
			2529 => x"ffd52795",
			2530 => x"0e00ac04",
			2531 => x"ff912795",
			2532 => x"00112795",
			2533 => x"05002518",
			2534 => x"01000704",
			2535 => x"ffbb2831",
			2536 => x"00011508",
			2537 => x"05002304",
			2538 => x"ff872831",
			2539 => x"005d2831",
			2540 => x"03002608",
			2541 => x"03002104",
			2542 => x"ffeb2831",
			2543 => x"00062831",
			2544 => x"00d72831",
			2545 => x"0a003118",
			2546 => x"09001b0c",
			2547 => x"0f00c208",
			2548 => x"0f00bb04",
			2549 => x"ffde2831",
			2550 => x"002b2831",
			2551 => x"ff3e2831",
			2552 => x"05002a08",
			2553 => x"05002804",
			2554 => x"ffee2831",
			2555 => x"004a2831",
			2556 => x"ffe22831",
			2557 => x"00013014",
			2558 => x"0d001608",
			2559 => x"0f00ca04",
			2560 => x"ffd72831",
			2561 => x"00cc2831",
			2562 => x"01001204",
			2563 => x"ffaf2831",
			2564 => x"01001304",
			2565 => x"00172831",
			2566 => x"fff92831",
			2567 => x"07003008",
			2568 => x"0f00c704",
			2569 => x"fff52831",
			2570 => x"002c2831",
			2571 => x"ff862831",
			2572 => x"0200f704",
			2573 => x"fe572885",
			2574 => x"05002e24",
			2575 => x"03002a18",
			2576 => x"09001808",
			2577 => x"01000704",
			2578 => x"fe812885",
			2579 => x"01db2885",
			2580 => x"0e009d0c",
			2581 => x"0a002f08",
			2582 => x"02012704",
			2583 => x"fefb2885",
			2584 => x"fe4f2885",
			2585 => x"fd012885",
			2586 => x"ffde2885",
			2587 => x"00013108",
			2588 => x"03002e04",
			2589 => x"02a82885",
			2590 => x"01702885",
			2591 => x"ff362885",
			2592 => x"fe742885",
			2593 => x"0e008a04",
			2594 => x"feb528c9",
			2595 => x"0700381c",
			2596 => x"03002404",
			2597 => x"ff3a28c9",
			2598 => x"01000804",
			2599 => x"fec428c9",
			2600 => x"07002f04",
			2601 => x"017028c9",
			2602 => x"07003308",
			2603 => x"0f00d204",
			2604 => x"00bf28c9",
			2605 => x"ff6328c9",
			2606 => x"0c001604",
			2607 => x"011628c9",
			2608 => x"ffc628c9",
			2609 => x"feb928c9",
			2610 => x"0f00bf04",
			2611 => x"fe8d292d",
			2612 => x"00013018",
			2613 => x"05002304",
			2614 => x"ff24292d",
			2615 => x"0d001508",
			2616 => x"00012604",
			2617 => x"016e292d",
			2618 => x"0054292d",
			2619 => x"0a003204",
			2620 => x"fef2292d",
			2621 => x"00012b04",
			2622 => x"00dd292d",
			2623 => x"ffe1292d",
			2624 => x"05002204",
			2625 => x"00dc292d",
			2626 => x"0e00ac10",
			2627 => x"0700300c",
			2628 => x"0d001204",
			2629 => x"fea4292d",
			2630 => x"0b001404",
			2631 => x"010a292d",
			2632 => x"ff7a292d",
			2633 => x"fe6a292d",
			2634 => x"008c292d",
			2635 => x"0f00bf04",
			2636 => x"fe7c2979",
			2637 => x"01000804",
			2638 => x"fe732979",
			2639 => x"0d001204",
			2640 => x"01cc2979",
			2641 => x"00014914",
			2642 => x"0d001304",
			2643 => x"ff4b2979",
			2644 => x"0d001508",
			2645 => x"0a003104",
			2646 => x"00692979",
			2647 => x"01c92979",
			2648 => x"0e00a004",
			2649 => x"fe942979",
			2650 => x"009a2979",
			2651 => x"0600cb04",
			2652 => x"fe7b2979",
			2653 => x"ffba2979",
			2654 => x"0200f704",
			2655 => x"ff2f29d5",
			2656 => x"02012f24",
			2657 => x"07003820",
			2658 => x"03002408",
			2659 => x"09001804",
			2660 => x"003c29d5",
			2661 => x"ff9029d5",
			2662 => x"03002f0c",
			2663 => x"01000804",
			2664 => x"ffca29d5",
			2665 => x"0e008a04",
			2666 => x"ffdc29d5",
			2667 => x"00ee29d5",
			2668 => x"07003404",
			2669 => x"ff7f29d5",
			2670 => x"03003304",
			2671 => x"006a29d5",
			2672 => x"ffef29d5",
			2673 => x"ffa629d5",
			2674 => x"0f00e904",
			2675 => x"ff4429d5",
			2676 => x"001129d5",
			2677 => x"0900180c",
			2678 => x"01000704",
			2679 => x"ff6a2a49",
			2680 => x"0f00c604",
			2681 => x"ffc02a49",
			2682 => x"01432a49",
			2683 => x"02012f2c",
			2684 => x"0d001208",
			2685 => x"0c001404",
			2686 => x"01372a49",
			2687 => x"ff832a49",
			2688 => x"07003314",
			2689 => x"03002908",
			2690 => x"00013204",
			2691 => x"fe9f2a49",
			2692 => x"00712a49",
			2693 => x"03002f08",
			2694 => x"01000d04",
			2695 => x"00f22a49",
			2696 => x"ff522a49",
			2697 => x"fef12a49",
			2698 => x"0700380c",
			2699 => x"01000a04",
			2700 => x"ff332a49",
			2701 => x"0d001604",
			2702 => x"01022a49",
			2703 => x"ffca2a49",
			2704 => x"fefa2a49",
			2705 => x"fec12a49",
			2706 => x"0300260c",
			2707 => x"09001808",
			2708 => x"07002904",
			2709 => x"ffe62ad5",
			2710 => x"005c2ad5",
			2711 => x"feec2ad5",
			2712 => x"01000a08",
			2713 => x"05002504",
			2714 => x"000d2ad5",
			2715 => x"ff1f2ad5",
			2716 => x"01000b14",
			2717 => x"0a003208",
			2718 => x"05002904",
			2719 => x"01302ad5",
			2720 => x"ffc22ad5",
			2721 => x"07003204",
			2722 => x"ff512ad5",
			2723 => x"08002004",
			2724 => x"00ba2ad5",
			2725 => x"fff82ad5",
			2726 => x"04001708",
			2727 => x"01000e04",
			2728 => x"00052ad5",
			2729 => x"00d92ad5",
			2730 => x"02010b08",
			2731 => x"02010004",
			2732 => x"ff932ad5",
			2733 => x"00e52ad5",
			2734 => x"07003108",
			2735 => x"00013504",
			2736 => x"ffb22ad5",
			2737 => x"003e2ad5",
			2738 => x"01001204",
			2739 => x"ff082ad5",
			2740 => x"fff42ad5",
			2741 => x"07003338",
			2742 => x"09001708",
			2743 => x"0d000f04",
			2744 => x"fffa2b81",
			2745 => x"00662b81",
			2746 => x"0d001420",
			2747 => x"0d001214",
			2748 => x"0a00310c",
			2749 => x"03002908",
			2750 => x"04001004",
			2751 => x"00042b81",
			2752 => x"ffb92b81",
			2753 => x"00152b81",
			2754 => x"0a003204",
			2755 => x"00332b81",
			2756 => x"fffc2b81",
			2757 => x"05002208",
			2758 => x"05001f04",
			2759 => x"fff42b81",
			2760 => x"000d2b81",
			2761 => x"ff632b81",
			2762 => x"0a002f08",
			2763 => x"04001404",
			2764 => x"00072b81",
			2765 => x"ffc32b81",
			2766 => x"04001d04",
			2767 => x"004f2b81",
			2768 => x"fff22b81",
			2769 => x"0001301c",
			2770 => x"0700350c",
			2771 => x"05002e08",
			2772 => x"0a002d04",
			2773 => x"fff82b81",
			2774 => x"00c02b81",
			2775 => x"ffec2b81",
			2776 => x"03002e04",
			2777 => x"ffc62b81",
			2778 => x"08001d04",
			2779 => x"fff82b81",
			2780 => x"04002504",
			2781 => x"002b2b81",
			2782 => x"fffb2b81",
			2783 => x"ffc22b81",
			2784 => x"01000804",
			2785 => x"fede2c07",
			2786 => x"0d00120c",
			2787 => x"05002808",
			2788 => x"0e008904",
			2789 => x"ffc32c07",
			2790 => x"015e2c07",
			2791 => x"ff952c07",
			2792 => x"07003320",
			2793 => x"01000908",
			2794 => x"04001c04",
			2795 => x"01052c07",
			2796 => x"ffd12c07",
			2797 => x"09001b0c",
			2798 => x"00012604",
			2799 => x"fe812c07",
			2800 => x"00013c04",
			2801 => x"00062c07",
			2802 => x"ff432c07",
			2803 => x"0b001508",
			2804 => x"03002a04",
			2805 => x"ffbf2c07",
			2806 => x"00e32c07",
			2807 => x"ff272c07",
			2808 => x"07003810",
			2809 => x"01000a04",
			2810 => x"ff102c07",
			2811 => x"0a002d04",
			2812 => x"ff382c07",
			2813 => x"00013004",
			2814 => x"01122c07",
			2815 => x"ff702c07",
			2816 => x"fed12c07",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(953, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1881, initial_addr_3'length));
	end generate gen_rom_6;

	gen_rom_7: if SELECT_ROM = 7 generate
		bank <= (
			0 => x"02010224",
			1 => x"0000fa1c",
			2 => x"01000504",
			3 => x"fe9d005d",
			4 => x"0e006d10",
			5 => x"0600780c",
			6 => x"0000d008",
			7 => x"07002d04",
			8 => x"fff5005d",
			9 => x"00da005d",
			10 => x"fea6005d",
			11 => x"00c5005d",
			12 => x"0b001404",
			13 => x"00fc005d",
			14 => x"fe80005d",
			15 => x"0e007404",
			16 => x"0131005d",
			17 => x"ff98005d",
			18 => x"01000608",
			19 => x"0d001304",
			20 => x"ff60005d",
			21 => x"007f005d",
			22 => x"fe9e005d",
			23 => x"06008628",
			24 => x"0000dd20",
			25 => x"0f00891c",
			26 => x"06007514",
			27 => x"0600700c",
			28 => x"06006d08",
			29 => x"0000b904",
			30 => x"001d00c1",
			31 => x"ff1200c1",
			32 => x"011300c1",
			33 => x"04003b04",
			34 => x"ff0100c1",
			35 => x"000c00c1",
			36 => x"0000d504",
			37 => x"00fb00c1",
			38 => x"003e00c1",
			39 => x"ff1000c1",
			40 => x"07002d04",
			41 => x"00f500c1",
			42 => x"ff7400c1",
			43 => x"01000808",
			44 => x"0b001604",
			45 => x"ff4a00c1",
			46 => x"008c00c1",
			47 => x"fed200c1",
			48 => x"0e007228",
			49 => x"04004720",
			50 => x"0400431c",
			51 => x"0c001308",
			52 => x"08001804",
			53 => x"004f0115",
			54 => x"01a50115",
			55 => x"04001704",
			56 => x"fe890115",
			57 => x"03003e08",
			58 => x"0a004204",
			59 => x"00270115",
			60 => x"014d0115",
			61 => x"04003e04",
			62 => x"fe910115",
			63 => x"00d60115",
			64 => x"fe3e0115",
			65 => x"07002f04",
			66 => x"01db0115",
			67 => x"fea70115",
			68 => x"fe6f0115",
			69 => x"0200ac38",
			70 => x"0e005228",
			71 => x"00008118",
			72 => x"0c001910",
			73 => x"08001604",
			74 => x"ffe801e1",
			75 => x"05000c04",
			76 => x"fff201e1",
			77 => x"01000704",
			78 => x"ffff01e1",
			79 => x"006501e1",
			80 => x"01001604",
			81 => x"ffdf01e1",
			82 => x"000101e1",
			83 => x"01000b08",
			84 => x"0e004d04",
			85 => x"ff9501e1",
			86 => x"fff701e1",
			87 => x"0e004804",
			88 => x"fffd01e1",
			89 => x"002501e1",
			90 => x"0d00190c",
			91 => x"08001b08",
			92 => x"06006204",
			93 => x"ffdf01e1",
			94 => x"001901e1",
			95 => x"009e01e1",
			96 => x"ffd301e1",
			97 => x"0e00650c",
			98 => x"01001208",
			99 => x"0000b904",
			100 => x"000201e1",
			101 => x"ff8901e1",
			102 => x"000c01e1",
			103 => x"06008618",
			104 => x"08001f10",
			105 => x"08001b08",
			106 => x"08001904",
			107 => x"002501e1",
			108 => x"ffcf01e1",
			109 => x"03003e04",
			110 => x"008001e1",
			111 => x"fff501e1",
			112 => x"0f007704",
			113 => x"000f01e1",
			114 => x"ffd201e1",
			115 => x"01000408",
			116 => x"05002e04",
			117 => x"fff801e1",
			118 => x"002201e1",
			119 => x"ffb501e1",
			120 => x"06008d38",
			121 => x"0500120c",
			122 => x"04000504",
			123 => x"00710255",
			124 => x"01000e04",
			125 => x"fe2c0255",
			126 => x"fffb0255",
			127 => x"08001814",
			128 => x"06006510",
			129 => x"06005c0c",
			130 => x"05001b04",
			131 => x"003c0255",
			132 => x"00009904",
			133 => x"fe950255",
			134 => x"ff460255",
			135 => x"00f00255",
			136 => x"fe720255",
			137 => x"0c001508",
			138 => x"08001b04",
			139 => x"00690255",
			140 => x"01750255",
			141 => x"05002504",
			142 => x"fe830255",
			143 => x"06008a08",
			144 => x"06008604",
			145 => x"002a0255",
			146 => x"fe850255",
			147 => x"01b50255",
			148 => x"fe800255",
			149 => x"05004338",
			150 => x"0b001730",
			151 => x"08001b10",
			152 => x"0c001104",
			153 => x"004a0311",
			154 => x"0f009e04",
			155 => x"ff5e0311",
			156 => x"03003104",
			157 => x"ffe90311",
			158 => x"00300311",
			159 => x"0d001618",
			160 => x"0d00130c",
			161 => x"02005c04",
			162 => x"002f0311",
			163 => x"0e006804",
			164 => x"ffc40311",
			165 => x"00120311",
			166 => x"01000904",
			167 => x"fff50311",
			168 => x"06008104",
			169 => x"00b00311",
			170 => x"fffc0311",
			171 => x"0000eb04",
			172 => x"ffc60311",
			173 => x"00290311",
			174 => x"08001904",
			175 => x"00060311",
			176 => x"ff660311",
			177 => x"0a00451c",
			178 => x"0b00180c",
			179 => x"03003908",
			180 => x"09001e04",
			181 => x"ffae0311",
			182 => x"00850311",
			183 => x"ff950311",
			184 => x"01000704",
			185 => x"ffe30311",
			186 => x"07003008",
			187 => x"03003a04",
			188 => x"00260311",
			189 => x"00a70311",
			190 => x"fff30311",
			191 => x"07002e04",
			192 => x"ff940311",
			193 => x"09002504",
			194 => x"003a0311",
			195 => x"ffdc0311",
			196 => x"0000be3c",
			197 => x"0e005a2c",
			198 => x"08001d20",
			199 => x"0a003614",
			200 => x"0e00480c",
			201 => x"07001604",
			202 => x"005d03f5",
			203 => x"01000a04",
			204 => x"ff7603f5",
			205 => x"000b03f5",
			206 => x"05002804",
			207 => x"000a03f5",
			208 => x"008503f5",
			209 => x"03003d08",
			210 => x"0c001704",
			211 => x"ffff03f5",
			212 => x"ff5403f5",
			213 => x"002903f5",
			214 => x"04002708",
			215 => x"0b001704",
			216 => x"007503f5",
			217 => x"ff7703f5",
			218 => x"009803f5",
			219 => x"08001908",
			220 => x"0000af04",
			221 => x"ffa003f5",
			222 => x"001403f5",
			223 => x"08001f04",
			224 => x"00d203f5",
			225 => x"ffe403f5",
			226 => x"0e006510",
			227 => x"0100120c",
			228 => x"07002c04",
			229 => x"ff2c03f5",
			230 => x"07002e04",
			231 => x"000203f5",
			232 => x"ffe703f5",
			233 => x"002603f5",
			234 => x"0e006d14",
			235 => x"08001b08",
			236 => x"0b001704",
			237 => x"ff7103f5",
			238 => x"001b03f5",
			239 => x"0f007b08",
			240 => x"06006f04",
			241 => x"002003f5",
			242 => x"ffc403f5",
			243 => x"00ba03f5",
			244 => x"01000408",
			245 => x"0b001404",
			246 => x"003f03f5",
			247 => x"fff303f5",
			248 => x"05004a04",
			249 => x"ff5203f5",
			250 => x"05004f04",
			251 => x"002c03f5",
			252 => x"ffe703f5",
			253 => x"06008d38",
			254 => x"0c001b28",
			255 => x"01000508",
			256 => x"0e006804",
			257 => x"fe530469",
			258 => x"017d0469",
			259 => x"0a00451c",
			260 => x"0200aa10",
			261 => x"0e005108",
			262 => x"00009e04",
			263 => x"010e0469",
			264 => x"fe4c0469",
			265 => x"0f006804",
			266 => x"02040469",
			267 => x"00f10469",
			268 => x"0e005c04",
			269 => x"fe1b0469",
			270 => x"0a003604",
			271 => x"ffba0469",
			272 => x"01c20469",
			273 => x"fe670469",
			274 => x"05004704",
			275 => x"fe4c0469",
			276 => x"0000c808",
			277 => x"0e005f04",
			278 => x"00330469",
			279 => x"01cb0469",
			280 => x"fe6c0469",
			281 => x"fe650469",
			282 => x"0200bb44",
			283 => x"05002214",
			284 => x"0c001308",
			285 => x"00004904",
			286 => x"07ab051d",
			287 => x"032e051d",
			288 => x"0c001404",
			289 => x"01b8051d",
			290 => x"0c001504",
			291 => x"ff7f051d",
			292 => x"fe48051d",
			293 => x"08001b10",
			294 => x"0d001308",
			295 => x"04003604",
			296 => x"fe48051d",
			297 => x"0026051d",
			298 => x"05004404",
			299 => x"ff4e051d",
			300 => x"0489051d",
			301 => x"0b001c1c",
			302 => x"01000a10",
			303 => x"0e004d08",
			304 => x"0a002d04",
			305 => x"040a051d",
			306 => x"fe39051d",
			307 => x"0000ae04",
			308 => x"0692051d",
			309 => x"016c051d",
			310 => x"03003a08",
			311 => x"0000a204",
			312 => x"06dd051d",
			313 => x"022f051d",
			314 => x"0975051d",
			315 => x"fe4f051d",
			316 => x"0e007214",
			317 => x"0f008e10",
			318 => x"0a002c04",
			319 => x"010b051d",
			320 => x"0a004808",
			321 => x"04003d04",
			322 => x"fe4b051d",
			323 => x"01e4051d",
			324 => x"fe4a051d",
			325 => x"0320051d",
			326 => x"fe49051d",
			327 => x"0200bb44",
			328 => x"05002110",
			329 => x"0c00140c",
			330 => x"08001604",
			331 => x"fe2105d9",
			332 => x"0c001104",
			333 => x"038005d9",
			334 => x"028905d9",
			335 => x"fe5405d9",
			336 => x"01000918",
			337 => x"0d00130c",
			338 => x"03003508",
			339 => x"08001904",
			340 => x"fe5a05d9",
			341 => x"017805d9",
			342 => x"fe3105d9",
			343 => x"05004404",
			344 => x"ffd805d9",
			345 => x"0000ad04",
			346 => x"033a05d9",
			347 => x"006b05d9",
			348 => x"0c001e18",
			349 => x"0c001608",
			350 => x"01000c04",
			351 => x"046705d9",
			352 => x"034e05d9",
			353 => x"05003708",
			354 => x"0b001704",
			355 => x"025a05d9",
			356 => x"fe9205d9",
			357 => x"0e005a04",
			358 => x"025905d9",
			359 => x"041a05d9",
			360 => x"fe5805d9",
			361 => x"0e007218",
			362 => x"0f007d08",
			363 => x"0000c704",
			364 => x"ffa805d9",
			365 => x"fe5105d9",
			366 => x"07002f0c",
			367 => x"08001b08",
			368 => x"0c001804",
			369 => x"fe4905d9",
			370 => x"023505d9",
			371 => x"03ba05d9",
			372 => x"fe5505d9",
			373 => x"fe5305d9",
			374 => x"0000be3c",
			375 => x"0e005a2c",
			376 => x"08001d20",
			377 => x"0a003614",
			378 => x"05002d0c",
			379 => x"0c001104",
			380 => x"007206b5",
			381 => x"01000d04",
			382 => x"ff6a06b5",
			383 => x"000b06b5",
			384 => x"09001c04",
			385 => x"000306b5",
			386 => x"007e06b5",
			387 => x"03003d08",
			388 => x"0c001704",
			389 => x"fffc06b5",
			390 => x"ff4406b5",
			391 => x"002906b5",
			392 => x"04002708",
			393 => x"0b001704",
			394 => x"007706b5",
			395 => x"ff7006b5",
			396 => x"00a006b5",
			397 => x"08001908",
			398 => x"0000af04",
			399 => x"ff9c06b5",
			400 => x"001306b5",
			401 => x"08001f04",
			402 => x"00db06b5",
			403 => x"ffe106b5",
			404 => x"0100040c",
			405 => x"0e006c04",
			406 => x"ffe006b5",
			407 => x"00012504",
			408 => x"007406b5",
			409 => x"fff906b5",
			410 => x"04001808",
			411 => x"0000e104",
			412 => x"004906b5",
			413 => x"ffe906b5",
			414 => x"01000608",
			415 => x"06007a04",
			416 => x"004806b5",
			417 => x"ff9006b5",
			418 => x"0600700c",
			419 => x"06006e08",
			420 => x"0e006204",
			421 => x"ff7d06b5",
			422 => x"001206b5",
			423 => x"007006b5",
			424 => x"06007e04",
			425 => x"ff2806b5",
			426 => x"06008604",
			427 => x"005306b5",
			428 => x"ff7506b5",
			429 => x"00009e34",
			430 => x"0500432c",
			431 => x"0b001518",
			432 => x"0800190c",
			433 => x"00003d04",
			434 => x"00a00781",
			435 => x"0d001104",
			436 => x"fe910781",
			437 => x"ffeb0781",
			438 => x"04001204",
			439 => x"004f0781",
			440 => x"02007a04",
			441 => x"01720781",
			442 => x"00ab0781",
			443 => x"0d001508",
			444 => x"01000b04",
			445 => x"fe7d0781",
			446 => x"ffda0781",
			447 => x"0e003d04",
			448 => x"feb60781",
			449 => x"05003204",
			450 => x"ff3f0781",
			451 => x"00e50781",
			452 => x"0c001804",
			453 => x"ff5c0781",
			454 => x"016c0781",
			455 => x"0400472c",
			456 => x"0e005108",
			457 => x"08002204",
			458 => x"fe5c0781",
			459 => x"007a0781",
			460 => x"0000ad0c",
			461 => x"05003e04",
			462 => x"ff410781",
			463 => x"0e005704",
			464 => x"001a0781",
			465 => x"017e0781",
			466 => x"0e005b08",
			467 => x"0b001b04",
			468 => x"fe490781",
			469 => x"00270781",
			470 => x"06007008",
			471 => x"01000904",
			472 => x"ff5e0781",
			473 => x"00cf0781",
			474 => x"06007804",
			475 => x"fe7d0781",
			476 => x"ffd80781",
			477 => x"03004904",
			478 => x"011a0781",
			479 => x"fef40781",
			480 => x"08001d50",
			481 => x"0e005b2c",
			482 => x"00009e18",
			483 => x"0e004d14",
			484 => x"0b001208",
			485 => x"00004904",
			486 => x"00a50885",
			487 => x"ffe50885",
			488 => x"01000a04",
			489 => x"ff230885",
			490 => x"0b001504",
			491 => x"00560885",
			492 => x"ff970885",
			493 => x"008f0885",
			494 => x"0a004210",
			495 => x"0700280c",
			496 => x"03003408",
			497 => x"07002504",
			498 => x"ffc30885",
			499 => x"00a60885",
			500 => x"ff750885",
			501 => x"ff0f0885",
			502 => x"002d0885",
			503 => x"0500380c",
			504 => x"01000b04",
			505 => x"ff050885",
			506 => x"07002a04",
			507 => x"00930885",
			508 => x"ff8a0885",
			509 => x"03003e0c",
			510 => x"08001804",
			511 => x"ffab0885",
			512 => x"02010204",
			513 => x"00ec0885",
			514 => x"ffd60885",
			515 => x"0000d008",
			516 => x"03004404",
			517 => x"007b0885",
			518 => x"ffaa0885",
			519 => x"ff440885",
			520 => x"0600651c",
			521 => x"0d001b14",
			522 => x"05001e0c",
			523 => x"00003908",
			524 => x"05001904",
			525 => x"fffa0885",
			526 => x"00080885",
			527 => x"ffd40885",
			528 => x"0b001a04",
			529 => x"01070885",
			530 => x"00050885",
			531 => x"04002804",
			532 => x"ff9c0885",
			533 => x"000f0885",
			534 => x"0a002c08",
			535 => x"0a002a04",
			536 => x"ffce0885",
			537 => x"00c80885",
			538 => x"0f007208",
			539 => x"0b002104",
			540 => x"00420885",
			541 => x"fffb0885",
			542 => x"05005904",
			543 => x"ff1a0885",
			544 => x"ffe00885",
			545 => x"0e007250",
			546 => x"0c001b3c",
			547 => x"01000b28",
			548 => x"0e005210",
			549 => x"0b001204",
			550 => x"01720931",
			551 => x"05001c04",
			552 => x"fe460931",
			553 => x"07002004",
			554 => x"01540931",
			555 => x"ff1d0931",
			556 => x"0d00130c",
			557 => x"0b001608",
			558 => x"04002b04",
			559 => x"ff7e0931",
			560 => x"02310931",
			561 => x"fe3e0931",
			562 => x"0b001604",
			563 => x"ff4e0931",
			564 => x"0a003b04",
			565 => x"02690931",
			566 => x"011e0931",
			567 => x"0f00650c",
			568 => x"05001304",
			569 => x"ffd40931",
			570 => x"04001304",
			571 => x"015b0931",
			572 => x"02190931",
			573 => x"08001f04",
			574 => x"01190931",
			575 => x"ff680931",
			576 => x"05004708",
			577 => x"05003a04",
			578 => x"fe5f0931",
			579 => x"fdf50931",
			580 => x"0000c808",
			581 => x"0e005f04",
			582 => x"00be0931",
			583 => x"022f0931",
			584 => x"fe650931",
			585 => x"0000bc04",
			586 => x"00bd0931",
			587 => x"fe600931",
			588 => x"07002f34",
			589 => x"0e007230",
			590 => x"00002504",
			591 => x"fe6009ad",
			592 => x"0800180c",
			593 => x"01000908",
			594 => x"0d001304",
			595 => x"fe4d09ad",
			596 => x"002309ad",
			597 => x"005e09ad",
			598 => x"0c001610",
			599 => x"01000908",
			600 => x"00008904",
			601 => x"019b09ad",
			602 => x"fefc09ad",
			603 => x"05002c04",
			604 => x"01fd09ad",
			605 => x"029309ad",
			606 => x"05003708",
			607 => x"0b001604",
			608 => x"00e409ad",
			609 => x"fe8809ad",
			610 => x"0d001704",
			611 => x"00ed09ad",
			612 => x"024909ad",
			613 => x"fe5d09ad",
			614 => x"0c001408",
			615 => x"00012a04",
			616 => x"011609ad",
			617 => x"fe8f09ad",
			618 => x"fe5d09ad",
			619 => x"0000b548",
			620 => x"08001914",
			621 => x"00003304",
			622 => x"00850aa1",
			623 => x"0100060c",
			624 => x"0b001508",
			625 => x"0a001b04",
			626 => x"003b0aa1",
			627 => x"ff4c0aa1",
			628 => x"00750aa1",
			629 => x"ff3d0aa1",
			630 => x"0700271c",
			631 => x"0c001608",
			632 => x"04001204",
			633 => x"00130aa1",
			634 => x"010a0aa1",
			635 => x"01000d0c",
			636 => x"04003408",
			637 => x"09001d04",
			638 => x"ffe30aa1",
			639 => x"fef20aa1",
			640 => x"00180aa1",
			641 => x"0e003704",
			642 => x"ffd50aa1",
			643 => x"00b40aa1",
			644 => x"0d001910",
			645 => x"01000708",
			646 => x"0c001b04",
			647 => x"005a0aa1",
			648 => x"ff610aa1",
			649 => x"0e005204",
			650 => x"ffe10aa1",
			651 => x"01440aa1",
			652 => x"01001604",
			653 => x"ff490aa1",
			654 => x"00140aa1",
			655 => x"06006b10",
			656 => x"0d001704",
			657 => x"feeb0aa1",
			658 => x"04004008",
			659 => x"0d001a04",
			660 => x"00710aa1",
			661 => x"fff60aa1",
			662 => x"ff940aa1",
			663 => x"06007008",
			664 => x"0000cb04",
			665 => x"01010aa1",
			666 => x"ffbe0aa1",
			667 => x"0100060c",
			668 => x"08001804",
			669 => x"ff800aa1",
			670 => x"0e007204",
			671 => x"00aa0aa1",
			672 => x"ffac0aa1",
			673 => x"06007804",
			674 => x"fec70aa1",
			675 => x"08001f08",
			676 => x"08001b04",
			677 => x"ff220aa1",
			678 => x"008b0aa1",
			679 => x"ff040aa1",
			680 => x"00009e2c",
			681 => x"08001604",
			682 => x"ffa70b75",
			683 => x"06005524",
			684 => x"00008318",
			685 => x"0c001910",
			686 => x"05001208",
			687 => x"0a000a04",
			688 => x"000e0b75",
			689 => x"ffcc0b75",
			690 => x"01000704",
			691 => x"00040b75",
			692 => x"00a50b75",
			693 => x"01001604",
			694 => x"ffc00b75",
			695 => x"00000b75",
			696 => x"01000b08",
			697 => x"00009304",
			698 => x"ff850b75",
			699 => x"fffc0b75",
			700 => x"00120b75",
			701 => x"00920b75",
			702 => x"04003e2c",
			703 => x"0e006510",
			704 => x"0d001704",
			705 => x"ff4d0b75",
			706 => x"0d001a08",
			707 => x"0000c204",
			708 => x"003e0b75",
			709 => x"ffe20b75",
			710 => x"ffc10b75",
			711 => x"0300240c",
			712 => x"03002304",
			713 => x"ffd50b75",
			714 => x"0000f404",
			715 => x"00680b75",
			716 => x"fff50b75",
			717 => x"0d001208",
			718 => x"06009a04",
			719 => x"00400b75",
			720 => x"fff60b75",
			721 => x"04003b04",
			722 => x"ff6a0b75",
			723 => x"00070b75",
			724 => x"0a004808",
			725 => x"03003e04",
			726 => x"fff00b75",
			727 => x"00690b75",
			728 => x"04004d04",
			729 => x"ff9e0b75",
			730 => x"04005a04",
			731 => x"00050b75",
			732 => x"fffa0b75",
			733 => x"0000be48",
			734 => x"0e005738",
			735 => x"00009e24",
			736 => x"0e004818",
			737 => x"0b001208",
			738 => x"00004804",
			739 => x"00870c59",
			740 => x"ffed0c59",
			741 => x"01000a08",
			742 => x"08001f04",
			743 => x"ff370c59",
			744 => x"00150c59",
			745 => x"04001904",
			746 => x"ffca0c59",
			747 => x"00670c59",
			748 => x"0c001808",
			749 => x"0a002d04",
			750 => x"00720c59",
			751 => x"ffa20c59",
			752 => x"00bc0c59",
			753 => x"08001b08",
			754 => x"0e005204",
			755 => x"ffc60c59",
			756 => x"00310c59",
			757 => x"08001d04",
			758 => x"ff2e0c59",
			759 => x"08002204",
			760 => x"00070c59",
			761 => x"ffe80c59",
			762 => x"01000908",
			763 => x"0a003d04",
			764 => x"ff720c59",
			765 => x"00650c59",
			766 => x"0d001804",
			767 => x"00b60c59",
			768 => x"ffb10c59",
			769 => x"0e006304",
			770 => x"ff130c59",
			771 => x"06007914",
			772 => x"0600750c",
			773 => x"0e006808",
			774 => x"0f007904",
			775 => x"00270c59",
			776 => x"ff6c0c59",
			777 => x"00550c59",
			778 => x"0000e304",
			779 => x"00ab0c59",
			780 => x"ffe60c59",
			781 => x"07002c10",
			782 => x"01000908",
			783 => x"00010e04",
			784 => x"007d0c59",
			785 => x"ffd20c59",
			786 => x"07002b04",
			787 => x"ff530c59",
			788 => x"006d0c59",
			789 => x"ff530c59",
			790 => x"0200ac38",
			791 => x"0e005228",
			792 => x"00008118",
			793 => x"0c001910",
			794 => x"08001604",
			795 => x"ffe90d35",
			796 => x"05000c04",
			797 => x"fff30d35",
			798 => x"01000704",
			799 => x"ffff0d35",
			800 => x"00610d35",
			801 => x"01001604",
			802 => x"ffdf0d35",
			803 => x"00010d35",
			804 => x"01000b08",
			805 => x"0e004d04",
			806 => x"ff990d35",
			807 => x"fff60d35",
			808 => x"0e004804",
			809 => x"fffd0d35",
			810 => x"00240d35",
			811 => x"0d00190c",
			812 => x"08001b08",
			813 => x"06006204",
			814 => x"ffdf0d35",
			815 => x"00180d35",
			816 => x"00960d35",
			817 => x"ffd50d35",
			818 => x"06006b04",
			819 => x"ff9d0d35",
			820 => x"04002518",
			821 => x"0300240c",
			822 => x"03002304",
			823 => x"ffda0d35",
			824 => x"07002b04",
			825 => x"fffc0d35",
			826 => x"00360d35",
			827 => x"0c001508",
			828 => x"0c001404",
			829 => x"ffef0d35",
			830 => x"000f0d35",
			831 => x"ff9d0d35",
			832 => x"0000cb04",
			833 => x"00710d35",
			834 => x"07002c0c",
			835 => x"0000dd04",
			836 => x"ffdd0d35",
			837 => x"00011204",
			838 => x"00530d35",
			839 => x"fff20d35",
			840 => x"04004704",
			841 => x"ff9f0d35",
			842 => x"0e006904",
			843 => x"ffe60d35",
			844 => x"002b0d35",
			845 => x"0200bb48",
			846 => x"05002110",
			847 => x"0c00140c",
			848 => x"08001604",
			849 => x"fe2a0df9",
			850 => x"01000a04",
			851 => x"02240df9",
			852 => x"03070df9",
			853 => x"fe570df9",
			854 => x"01000918",
			855 => x"0d001514",
			856 => x"0000a60c",
			857 => x"0e004d08",
			858 => x"00008304",
			859 => x"00990df9",
			860 => x"fe340df9",
			861 => x"02900df9",
			862 => x"0e005b04",
			863 => x"fe3a0df9",
			864 => x"00480df9",
			865 => x"02280df9",
			866 => x"0c001e1c",
			867 => x"0c00160c",
			868 => x"0a002a08",
			869 => x"01000e04",
			870 => x"04070df9",
			871 => x"02de0df9",
			872 => x"027c0df9",
			873 => x"05003708",
			874 => x"0b001704",
			875 => x"01e80df9",
			876 => x"fe9f0df9",
			877 => x"0e005a04",
			878 => x"01ef0df9",
			879 => x"03740df9",
			880 => x"fe5b0df9",
			881 => x"0e007218",
			882 => x"0f007d08",
			883 => x"0000c704",
			884 => x"ffbd0df9",
			885 => x"fe550df9",
			886 => x"07002f0c",
			887 => x"08001b08",
			888 => x"0c001804",
			889 => x"fe4f0df9",
			890 => x"01d30df9",
			891 => x"02c20df9",
			892 => x"fe5a0df9",
			893 => x"fe550df9",
			894 => x"07003030",
			895 => x"06008d2c",
			896 => x"00002504",
			897 => x"fe640e5d",
			898 => x"08001810",
			899 => x"08001604",
			900 => x"fe520e5d",
			901 => x"0000a608",
			902 => x"0c001604",
			903 => x"00260e5d",
			904 => x"015b0e5d",
			905 => x"fe520e5d",
			906 => x"0c00150c",
			907 => x"08001b04",
			908 => x"014b0e5d",
			909 => x"0d001304",
			910 => x"01d40e5d",
			911 => x"02450e5d",
			912 => x"05002504",
			913 => x"fe5d0e5d",
			914 => x"0e006b04",
			915 => x"00c10e5d",
			916 => x"02110e5d",
			917 => x"fe610e5d",
			918 => x"fe600e5d",
			919 => x"06008d34",
			920 => x"08001604",
			921 => x"fe7b0ec9",
			922 => x"04000a08",
			923 => x"02002504",
			924 => x"00c40ec9",
			925 => x"fdfc0ec9",
			926 => x"0c001508",
			927 => x"08001b04",
			928 => x"00270ec9",
			929 => x"01850ec9",
			930 => x"05003710",
			931 => x"09001e08",
			932 => x"01000a04",
			933 => x"febb0ec9",
			934 => x"00de0ec9",
			935 => x"07002904",
			936 => x"ff3f0ec9",
			937 => x"fe4f0ec9",
			938 => x"01000808",
			939 => x"07002b04",
			940 => x"01280ec9",
			941 => x"ffc70ec9",
			942 => x"0d001404",
			943 => x"ff0f0ec9",
			944 => x"00550ec9",
			945 => x"fe7d0ec9",
			946 => x"0200a844",
			947 => x"0e005538",
			948 => x"09002020",
			949 => x"0f005d1c",
			950 => x"00008310",
			951 => x"05001208",
			952 => x"07001704",
			953 => x"001f0fd5",
			954 => x"ffb00fd5",
			955 => x"09001e04",
			956 => x"007c0fd5",
			957 => x"ffdc0fd5",
			958 => x"0d001508",
			959 => x"01000604",
			960 => x"00060fd5",
			961 => x"ff620fd5",
			962 => x"00280fd5",
			963 => x"00790fd5",
			964 => x"08001d08",
			965 => x"09002304",
			966 => x"ff6c0fd5",
			967 => x"00110fd5",
			968 => x"07002908",
			969 => x"00006e04",
			970 => x"fff90fd5",
			971 => x"00410fd5",
			972 => x"08002004",
			973 => x"00010fd5",
			974 => x"ffd10fd5",
			975 => x"0d001808",
			976 => x"09001e04",
			977 => x"00000fd5",
			978 => x"00ca0fd5",
			979 => x"ffd30fd5",
			980 => x"0e006518",
			981 => x"0d001508",
			982 => x"09002104",
			983 => x"ff4d0fd5",
			984 => x"000e0fd5",
			985 => x"04002504",
			986 => x"ffa20fd5",
			987 => x"0d001804",
			988 => x"00630fd5",
			989 => x"0e005c04",
			990 => x"00030fd5",
			991 => x"ffb70fd5",
			992 => x"06007910",
			993 => x"0f007b08",
			994 => x"0f007704",
			995 => x"00230fd5",
			996 => x"ffb90fd5",
			997 => x"0c001b04",
			998 => x"00830fd5",
			999 => x"ffe50fd5",
			1000 => x"07002c10",
			1001 => x"05002904",
			1002 => x"ff980fd5",
			1003 => x"0d001308",
			1004 => x"0d001204",
			1005 => x"00310fd5",
			1006 => x"ffba0fd5",
			1007 => x"006f0fd5",
			1008 => x"0c001408",
			1009 => x"04001904",
			1010 => x"fffa0fd5",
			1011 => x"00210fd5",
			1012 => x"ff730fd5",
			1013 => x"06008d44",
			1014 => x"0d001938",
			1015 => x"04004730",
			1016 => x"01000b18",
			1017 => x"0400290c",
			1018 => x"0c001104",
			1019 => x"01611061",
			1020 => x"0a002a04",
			1021 => x"ff5b1061",
			1022 => x"fe1b1061",
			1023 => x"07002504",
			1024 => x"fe701061",
			1025 => x"03003804",
			1026 => x"00cc1061",
			1027 => x"ffb91061",
			1028 => x"0000be10",
			1029 => x"0c001908",
			1030 => x"0a001404",
			1031 => x"00311061",
			1032 => x"01791061",
			1033 => x"0d001704",
			1034 => x"ff621061",
			1035 => x"00f51061",
			1036 => x"06007804",
			1037 => x"fed91061",
			1038 => x"008d1061",
			1039 => x"07002f04",
			1040 => x"01991061",
			1041 => x"fee51061",
			1042 => x"07002808",
			1043 => x"06004304",
			1044 => x"ff381061",
			1045 => x"01051061",
			1046 => x"fe551061",
			1047 => x"fe771061",
			1048 => x"08001810",
			1049 => x"0700260c",
			1050 => x"08001604",
			1051 => x"ff271115",
			1052 => x"0c001604",
			1053 => x"000d1115",
			1054 => x"009d1115",
			1055 => x"feb81115",
			1056 => x"04004744",
			1057 => x"03003e34",
			1058 => x"04003420",
			1059 => x"0b001710",
			1060 => x"01000b08",
			1061 => x"00010104",
			1062 => x"ff9d1115",
			1063 => x"00c21115",
			1064 => x"04002104",
			1065 => x"00191115",
			1066 => x"01581115",
			1067 => x"04003108",
			1068 => x"08001904",
			1069 => x"00211115",
			1070 => x"fee01115",
			1071 => x"03003504",
			1072 => x"008a1115",
			1073 => x"ff951115",
			1074 => x"09001e04",
			1075 => x"ff881115",
			1076 => x"05004c08",
			1077 => x"0000ae04",
			1078 => x"01501115",
			1079 => x"00291115",
			1080 => x"03003a04",
			1081 => x"ff3f1115",
			1082 => x"00691115",
			1083 => x"04003e08",
			1084 => x"0c001b04",
			1085 => x"feaf1115",
			1086 => x"ffd51115",
			1087 => x"0000c004",
			1088 => x"008e1115",
			1089 => x"ff231115",
			1090 => x"07002f04",
			1091 => x"01191115",
			1092 => x"ff461115",
			1093 => x"00008318",
			1094 => x"05001208",
			1095 => x"07001804",
			1096 => x"002311e1",
			1097 => x"ff6e11e1",
			1098 => x"0c001908",
			1099 => x"08001804",
			1100 => x"000011e1",
			1101 => x"00e911e1",
			1102 => x"01001604",
			1103 => x"ff9211e1",
			1104 => x"001c11e1",
			1105 => x"0e004d08",
			1106 => x"08001f04",
			1107 => x"ff0c11e1",
			1108 => x"001611e1",
			1109 => x"05003828",
			1110 => x"01000b0c",
			1111 => x"05002208",
			1112 => x"05002104",
			1113 => x"ffc711e1",
			1114 => x"001f11e1",
			1115 => x"fef111e1",
			1116 => x"0d00160c",
			1117 => x"05002204",
			1118 => x"ff9311e1",
			1119 => x"0a002d04",
			1120 => x"00ff11e1",
			1121 => x"ffac11e1",
			1122 => x"0000eb08",
			1123 => x"0f006504",
			1124 => x"003f11e1",
			1125 => x"ff0a11e1",
			1126 => x"02010204",
			1127 => x"006d11e1",
			1128 => x"ffdc11e1",
			1129 => x"00009e04",
			1130 => x"00d611e1",
			1131 => x"06007510",
			1132 => x"0000b908",
			1133 => x"06006404",
			1134 => x"ffcd11e1",
			1135 => x"00e511e1",
			1136 => x"08001f04",
			1137 => x"ff2d11e1",
			1138 => x"002211e1",
			1139 => x"08001f08",
			1140 => x"0c001b04",
			1141 => x"009811e1",
			1142 => x"ffc511e1",
			1143 => x"ff8c11e1",
			1144 => x"0000ca3c",
			1145 => x"00002504",
			1146 => x"fe5b127d",
			1147 => x"01000504",
			1148 => x"fe46127d",
			1149 => x"0b00191c",
			1150 => x"01000b10",
			1151 => x"0e004e08",
			1152 => x"0c001404",
			1153 => x"0249127d",
			1154 => x"ff06127d",
			1155 => x"0d001404",
			1156 => x"00aa127d",
			1157 => x"029f127d",
			1158 => x"0000a208",
			1159 => x"0a001404",
			1160 => x"0187127d",
			1161 => x"02b7127d",
			1162 => x"012a127d",
			1163 => x"0400310c",
			1164 => x"01001608",
			1165 => x"04002004",
			1166 => x"fe5e127d",
			1167 => x"fe07127d",
			1168 => x"ffbd127d",
			1169 => x"0a004c08",
			1170 => x"03003d04",
			1171 => x"0126127d",
			1172 => x"0216127d",
			1173 => x"fe54127d",
			1174 => x"0e007210",
			1175 => x"06007504",
			1176 => x"fe58127d",
			1177 => x"01000904",
			1178 => x"024a127d",
			1179 => x"0f008704",
			1180 => x"00b5127d",
			1181 => x"fe1a127d",
			1182 => x"fe5a127d",
			1183 => x"06008d3c",
			1184 => x"08001604",
			1185 => x"fe7512f9",
			1186 => x"0d00192c",
			1187 => x"08001d14",
			1188 => x"0a004510",
			1189 => x"0a004208",
			1190 => x"09002004",
			1191 => x"003a12f9",
			1192 => x"ff1712f9",
			1193 => x"05005204",
			1194 => x"018712f9",
			1195 => x"00aa12f9",
			1196 => x"fe7e12f9",
			1197 => x"01000a0c",
			1198 => x"07002704",
			1199 => x"003312f9",
			1200 => x"09002304",
			1201 => x"01ee12f9",
			1202 => x"ff8812f9",
			1203 => x"06007008",
			1204 => x"0d001504",
			1205 => x"ffb212f9",
			1206 => x"014512f9",
			1207 => x"ff8b12f9",
			1208 => x"07002908",
			1209 => x"0c001c04",
			1210 => x"012412f9",
			1211 => x"ff3912f9",
			1212 => x"fe5c12f9",
			1213 => x"fe7a12f9",
			1214 => x"06008664",
			1215 => x"0d00142c",
			1216 => x"0300351c",
			1217 => x"03003218",
			1218 => x"08001b0c",
			1219 => x"0c001104",
			1220 => x"00a513dd",
			1221 => x"09001c04",
			1222 => x"fecc13dd",
			1223 => x"ffd113dd",
			1224 => x"0c001604",
			1225 => x"010413dd",
			1226 => x"07002704",
			1227 => x"ff4613dd",
			1228 => x"005813dd",
			1229 => x"011113dd",
			1230 => x"0900210c",
			1231 => x"04003c04",
			1232 => x"fe9d13dd",
			1233 => x"04004004",
			1234 => x"ffbd13dd",
			1235 => x"ff2813dd",
			1236 => x"001413dd",
			1237 => x"0b001918",
			1238 => x"04003c14",
			1239 => x"0200aa0c",
			1240 => x"04002c08",
			1241 => x"0c001604",
			1242 => x"010c13dd",
			1243 => x"ffb313dd",
			1244 => x"012513dd",
			1245 => x"0000c804",
			1246 => x"ff3213dd",
			1247 => x"008a13dd",
			1248 => x"010d13dd",
			1249 => x"03003b14",
			1250 => x"08001d04",
			1251 => x"feae13dd",
			1252 => x"08001f08",
			1253 => x"0d001704",
			1254 => x"fff913dd",
			1255 => x"006013dd",
			1256 => x"01001604",
			1257 => x"ff7a13dd",
			1258 => x"002313dd",
			1259 => x"0a004704",
			1260 => x"00f913dd",
			1261 => x"0000c004",
			1262 => x"005113dd",
			1263 => x"ff1713dd",
			1264 => x"0100080c",
			1265 => x"0a003604",
			1266 => x"ff6e13dd",
			1267 => x"0a003b04",
			1268 => x"003713dd",
			1269 => x"ffee13dd",
			1270 => x"fee413dd",
			1271 => x"06008d54",
			1272 => x"0d001948",
			1273 => x"01000b2c",
			1274 => x"0e005a18",
			1275 => x"0200970c",
			1276 => x"0f005d08",
			1277 => x"0b001204",
			1278 => x"015c1489",
			1279 => x"ff631489",
			1280 => x"01671489",
			1281 => x"01000a08",
			1282 => x"06006204",
			1283 => x"ffc91489",
			1284 => x"fda71489",
			1285 => x"fe001489",
			1286 => x"05003808",
			1287 => x"0000af04",
			1288 => x"fff31489",
			1289 => x"fe171489",
			1290 => x"0000be04",
			1291 => x"018e1489",
			1292 => x"0e006304",
			1293 => x"fe5f1489",
			1294 => x"00da1489",
			1295 => x"0200a110",
			1296 => x"0c001a08",
			1297 => x"0a001404",
			1298 => x"00611489",
			1299 => x"019c1489",
			1300 => x"05001904",
			1301 => x"feef1489",
			1302 => x"00191489",
			1303 => x"0e005b04",
			1304 => x"fe591489",
			1305 => x"0d001604",
			1306 => x"012e1489",
			1307 => x"ffdd1489",
			1308 => x"07002908",
			1309 => x"0c001c04",
			1310 => x"01501489",
			1311 => x"feee1489",
			1312 => x"fe431489",
			1313 => x"fe6c1489",
			1314 => x"08001810",
			1315 => x"00003d04",
			1316 => x"0040156d",
			1317 => x"03003408",
			1318 => x"03003104",
			1319 => x"ff78156d",
			1320 => x"0043156d",
			1321 => x"ff3b156d",
			1322 => x"0b001944",
			1323 => x"0f008930",
			1324 => x"07002718",
			1325 => x"0000890c",
			1326 => x"04000a04",
			1327 => x"ff94156d",
			1328 => x"09001e04",
			1329 => x"00c3156d",
			1330 => x"ffb8156d",
			1331 => x"0d001508",
			1332 => x"02009704",
			1333 => x"fffb156d",
			1334 => x"ff30156d",
			1335 => x"002d156d",
			1336 => x"08001b0c",
			1337 => x"0e005f08",
			1338 => x"0000a404",
			1339 => x"0008156d",
			1340 => x"ff7d156d",
			1341 => x"0032156d",
			1342 => x"01000c08",
			1343 => x"06005304",
			1344 => x"fff5156d",
			1345 => x"00da156d",
			1346 => x"0036156d",
			1347 => x"0500380c",
			1348 => x"0c001408",
			1349 => x"00011504",
			1350 => x"002c156d",
			1351 => x"fff2156d",
			1352 => x"ff28156d",
			1353 => x"0c001804",
			1354 => x"0086156d",
			1355 => x"ffc8156d",
			1356 => x"0c001a08",
			1357 => x"06004d04",
			1358 => x"ffec156d",
			1359 => x"004e156d",
			1360 => x"09001f04",
			1361 => x"005b156d",
			1362 => x"07002904",
			1363 => x"ff10156d",
			1364 => x"07002b08",
			1365 => x"0e004a04",
			1366 => x"fff9156d",
			1367 => x"0067156d",
			1368 => x"04004c04",
			1369 => x"ff71156d",
			1370 => x"0044156d",
			1371 => x"00009e30",
			1372 => x"08001604",
			1373 => x"ff521661",
			1374 => x"04003628",
			1375 => x"0c00160c",
			1376 => x"01000908",
			1377 => x"00006504",
			1378 => x"006c1661",
			1379 => x"ff601661",
			1380 => x"00eb1661",
			1381 => x"01000b0c",
			1382 => x"00009408",
			1383 => x"07002704",
			1384 => x"ff1c1661",
			1385 => x"001c1661",
			1386 => x"00211661",
			1387 => x"07002908",
			1388 => x"0e003704",
			1389 => x"ffd01661",
			1390 => x"00c71661",
			1391 => x"08001f04",
			1392 => x"00061661",
			1393 => x"ff831661",
			1394 => x"00e51661",
			1395 => x"0e005718",
			1396 => x"0100080c",
			1397 => x"04003308",
			1398 => x"04002104",
			1399 => x"fff21661",
			1400 => x"00671661",
			1401 => x"ff8e1661",
			1402 => x"0d001704",
			1403 => x"fef01661",
			1404 => x"0d001a04",
			1405 => x"002f1661",
			1406 => x"ffa91661",
			1407 => x"0000b20c",
			1408 => x"01000904",
			1409 => x"ffd41661",
			1410 => x"03003a04",
			1411 => x"01061661",
			1412 => x"002b1661",
			1413 => x"0400441c",
			1414 => x"01000b0c",
			1415 => x"0d001708",
			1416 => x"06008a04",
			1417 => x"ff211661",
			1418 => x"002c1661",
			1419 => x"00661661",
			1420 => x"0a002c08",
			1421 => x"05002804",
			1422 => x"ff4a1661",
			1423 => x"00ff1661",
			1424 => x"06007004",
			1425 => x"00591661",
			1426 => x"ff071661",
			1427 => x"03004908",
			1428 => x"0b001a04",
			1429 => x"00b81661",
			1430 => x"ffff1661",
			1431 => x"ff9d1661",
			1432 => x"06008d44",
			1433 => x"09002440",
			1434 => x"0e006524",
			1435 => x"0200b714",
			1436 => x"01000504",
			1437 => x"fe6416ed",
			1438 => x"0c001408",
			1439 => x"0d001104",
			1440 => x"008416ed",
			1441 => x"01b116ed",
			1442 => x"05002504",
			1443 => x"fe9516ed",
			1444 => x"004516ed",
			1445 => x"08001f0c",
			1446 => x"07002c08",
			1447 => x"0a002f04",
			1448 => x"fd7f16ed",
			1449 => x"fe5416ed",
			1450 => x"ff2616ed",
			1451 => x"fff716ed",
			1452 => x"06007908",
			1453 => x"0a004304",
			1454 => x"021116ed",
			1455 => x"007516ed",
			1456 => x"0f008e08",
			1457 => x"04001d04",
			1458 => x"001e16ed",
			1459 => x"fe5016ed",
			1460 => x"09001b04",
			1461 => x"fe5b16ed",
			1462 => x"01000904",
			1463 => x"01ff16ed",
			1464 => x"003d16ed",
			1465 => x"fe6e16ed",
			1466 => x"fe6a16ed",
			1467 => x"08001808",
			1468 => x"00003d04",
			1469 => x"004217c1",
			1470 => x"ff5017c1",
			1471 => x"0b001944",
			1472 => x"0f008930",
			1473 => x"07002718",
			1474 => x"0000890c",
			1475 => x"04000a04",
			1476 => x"ff9117c1",
			1477 => x"09001e04",
			1478 => x"00cd17c1",
			1479 => x"ffb317c1",
			1480 => x"0d001508",
			1481 => x"02009704",
			1482 => x"fffa17c1",
			1483 => x"ff2617c1",
			1484 => x"003317c1",
			1485 => x"08001b0c",
			1486 => x"0e005f08",
			1487 => x"0000af04",
			1488 => x"000617c1",
			1489 => x"ff7317c1",
			1490 => x"003617c1",
			1491 => x"01000c08",
			1492 => x"06005304",
			1493 => x"fff517c1",
			1494 => x"00e617c1",
			1495 => x"003c17c1",
			1496 => x"0500380c",
			1497 => x"0c001408",
			1498 => x"00011504",
			1499 => x"002d17c1",
			1500 => x"fff117c1",
			1501 => x"ff2017c1",
			1502 => x"0c001804",
			1503 => x"008b17c1",
			1504 => x"ffc217c1",
			1505 => x"0c001a08",
			1506 => x"06004d04",
			1507 => x"ffed17c1",
			1508 => x"005217c1",
			1509 => x"09001f04",
			1510 => x"006117c1",
			1511 => x"07002904",
			1512 => x"ff0517c1",
			1513 => x"07002b08",
			1514 => x"0e004a04",
			1515 => x"fff817c1",
			1516 => x"006c17c1",
			1517 => x"04004c04",
			1518 => x"ff6717c1",
			1519 => x"004817c1",
			1520 => x"0e007248",
			1521 => x"0c001e44",
			1522 => x"08001810",
			1523 => x"09001e08",
			1524 => x"04000a04",
			1525 => x"ff971855",
			1526 => x"fe561855",
			1527 => x"0b001704",
			1528 => x"01cc1855",
			1529 => x"fe551855",
			1530 => x"0c001614",
			1531 => x"0000890c",
			1532 => x"05001304",
			1533 => x"00421855",
			1534 => x"00005c04",
			1535 => x"01bc1855",
			1536 => x"02131855",
			1537 => x"01000904",
			1538 => x"fef71855",
			1539 => x"00b81855",
			1540 => x"05003710",
			1541 => x"0b001608",
			1542 => x"01000b04",
			1543 => x"fe2e1855",
			1544 => x"01171855",
			1545 => x"09001d04",
			1546 => x"000d1855",
			1547 => x"fe601855",
			1548 => x"0e005a08",
			1549 => x"00009f04",
			1550 => x"01291855",
			1551 => x"ff401855",
			1552 => x"0000ba04",
			1553 => x"02281855",
			1554 => x"00b41855",
			1555 => x"fe661855",
			1556 => x"fe621855",
			1557 => x"06008d60",
			1558 => x"07002724",
			1559 => x"03003820",
			1560 => x"0c001a1c",
			1561 => x"0c001810",
			1562 => x"03002c08",
			1563 => x"05002b04",
			1564 => x"ffc51919",
			1565 => x"01691919",
			1566 => x"03003304",
			1567 => x"fe9d1919",
			1568 => x"ffd21919",
			1569 => x"0e004808",
			1570 => x"0d001504",
			1571 => x"ff0a1919",
			1572 => x"00581919",
			1573 => x"017e1919",
			1574 => x"fea71919",
			1575 => x"fe711919",
			1576 => x"05004820",
			1577 => x"09001e0c",
			1578 => x"07002b08",
			1579 => x"07002904",
			1580 => x"00be1919",
			1581 => x"ff501919",
			1582 => x"01641919",
			1583 => x"0000b20c",
			1584 => x"04002608",
			1585 => x"07002d04",
			1586 => x"fe9e1919",
			1587 => x"001e1919",
			1588 => x"00f31919",
			1589 => x"07002a04",
			1590 => x"ff581919",
			1591 => x"fe5c1919",
			1592 => x"09002008",
			1593 => x"01000504",
			1594 => x"fee51919",
			1595 => x"01811919",
			1596 => x"09002108",
			1597 => x"0c001a04",
			1598 => x"000d1919",
			1599 => x"fe8d1919",
			1600 => x"0200cc08",
			1601 => x"0a004804",
			1602 => x"01201919",
			1603 => x"ff8d1919",
			1604 => x"fecb1919",
			1605 => x"fe901919",
			1606 => x"0e007750",
			1607 => x"0900244c",
			1608 => x"0e006530",
			1609 => x"0200b720",
			1610 => x"01000b10",
			1611 => x"0e005a08",
			1612 => x"0000ae04",
			1613 => x"ffe319bd",
			1614 => x"fe7019bd",
			1615 => x"01000904",
			1616 => x"002319bd",
			1617 => x"01af19bd",
			1618 => x"02008f08",
			1619 => x"05001304",
			1620 => x"ff6819bd",
			1621 => x"019719bd",
			1622 => x"04002304",
			1623 => x"fe2a19bd",
			1624 => x"00d419bd",
			1625 => x"08001f0c",
			1626 => x"07002c08",
			1627 => x"0a002f04",
			1628 => x"fd5119bd",
			1629 => x"fe4c19bd",
			1630 => x"ff1b19bd",
			1631 => x"ffec19bd",
			1632 => x"06007908",
			1633 => x"0a004304",
			1634 => x"024619bd",
			1635 => x"007f19bd",
			1636 => x"0000fa0c",
			1637 => x"09001b04",
			1638 => x"fe5219bd",
			1639 => x"0f008e04",
			1640 => x"feef19bd",
			1641 => x"00e219bd",
			1642 => x"03002904",
			1643 => x"feec19bd",
			1644 => x"01d619bd",
			1645 => x"fe6c19bd",
			1646 => x"fe6919bd",
			1647 => x"04004780",
			1648 => x"00009e30",
			1649 => x"06005524",
			1650 => x"0000831c",
			1651 => x"04000a0c",
			1652 => x"02002508",
			1653 => x"0a000d04",
			1654 => x"00b81ac9",
			1655 => x"ffea1ac9",
			1656 => x"fe831ac9",
			1657 => x"09001e08",
			1658 => x"01000704",
			1659 => x"ff9d1ac9",
			1660 => x"011d1ac9",
			1661 => x"01001404",
			1662 => x"fed41ac9",
			1663 => x"008e1ac9",
			1664 => x"0c001804",
			1665 => x"fe8c1ac9",
			1666 => x"00191ac9",
			1667 => x"03002404",
			1668 => x"ffef1ac9",
			1669 => x"06005a04",
			1670 => x"00bd1ac9",
			1671 => x"01811ac9",
			1672 => x"0e005a20",
			1673 => x"08001d14",
			1674 => x"0a00370c",
			1675 => x"06005d08",
			1676 => x"09001e04",
			1677 => x"ff7a1ac9",
			1678 => x"01301ac9",
			1679 => x"feb51ac9",
			1680 => x"0e005604",
			1681 => x"fe2a1ac9",
			1682 => x"fef61ac9",
			1683 => x"07002804",
			1684 => x"ff241ac9",
			1685 => x"08002004",
			1686 => x"01451ac9",
			1687 => x"ffc51ac9",
			1688 => x"05003718",
			1689 => x"0300240c",
			1690 => x"09001c08",
			1691 => x"0000b104",
			1692 => x"007a1ac9",
			1693 => x"fe8f1ac9",
			1694 => x"01501ac9",
			1695 => x"04001b08",
			1696 => x"0f00ad04",
			1697 => x"00bd1ac9",
			1698 => x"ff1b1ac9",
			1699 => x"fe4a1ac9",
			1700 => x"0200bb0c",
			1701 => x"08001b04",
			1702 => x"00341ac9",
			1703 => x"0200af04",
			1704 => x"01931ac9",
			1705 => x"00f71ac9",
			1706 => x"0f008804",
			1707 => x"fe671ac9",
			1708 => x"01000904",
			1709 => x"01321ac9",
			1710 => x"ff171ac9",
			1711 => x"07002f04",
			1712 => x"01421ac9",
			1713 => x"fef01ac9",
			1714 => x"06008d54",
			1715 => x"0c001e50",
			1716 => x"0b001414",
			1717 => x"08001604",
			1718 => x"fe711b77",
			1719 => x"0500280c",
			1720 => x"0c001408",
			1721 => x"08001b04",
			1722 => x"01221b77",
			1723 => x"01d61b77",
			1724 => x"ffc91b77",
			1725 => x"02201b77",
			1726 => x"0400211c",
			1727 => x"0b001610",
			1728 => x"09001c08",
			1729 => x"02007a04",
			1730 => x"00431b77",
			1731 => x"fe181b77",
			1732 => x"0d001304",
			1733 => x"fefc1b77",
			1734 => x"01131b77",
			1735 => x"0c001704",
			1736 => x"ffd11b77",
			1737 => x"0d001904",
			1738 => x"fe621b77",
			1739 => x"fd9d1b77",
			1740 => x"0d001510",
			1741 => x"03003e08",
			1742 => x"04003404",
			1743 => x"ffb11b77",
			1744 => x"00e91b77",
			1745 => x"0c001904",
			1746 => x"fe361b77",
			1747 => x"ffa11b77",
			1748 => x"0b001908",
			1749 => x"04002b04",
			1750 => x"00801b77",
			1751 => x"01d81b77",
			1752 => x"01000a04",
			1753 => x"fede1b77",
			1754 => x"00d51b77",
			1755 => x"fe6c1b77",
			1756 => x"fe671b77",
			1757 => x"06008624",
			1758 => x"0000dd1c",
			1759 => x"0f008918",
			1760 => x"06007510",
			1761 => x"0000ca0c",
			1762 => x"01000504",
			1763 => x"ff041bd1",
			1764 => x"0a004504",
			1765 => x"00271bd1",
			1766 => x"ff6c1bd1",
			1767 => x"fed41bd1",
			1768 => x"0000d504",
			1769 => x"010a1bd1",
			1770 => x"00491bd1",
			1771 => x"feff1bd1",
			1772 => x"07002d04",
			1773 => x"01071bd1",
			1774 => x"ff6e1bd1",
			1775 => x"01000808",
			1776 => x"0b001604",
			1777 => x"ff421bd1",
			1778 => x"00991bd1",
			1779 => x"fec61bd1",
			1780 => x"0400472c",
			1781 => x"02010220",
			1782 => x"0000fa18",
			1783 => x"01000504",
			1784 => x"fe9a1c35",
			1785 => x"04004310",
			1786 => x"0000ae08",
			1787 => x"0f005d04",
			1788 => x"ffca1c35",
			1789 => x"00b31c35",
			1790 => x"06006404",
			1791 => x"fe681c35",
			1792 => x"fff81c35",
			1793 => x"feda1c35",
			1794 => x"06008f04",
			1795 => x"013e1c35",
			1796 => x"ffa91c35",
			1797 => x"01000608",
			1798 => x"0b001504",
			1799 => x"ff621c35",
			1800 => x"007d1c35",
			1801 => x"fe961c35",
			1802 => x"03004904",
			1803 => x"01381c35",
			1804 => x"ff211c35",
			1805 => x"0000be38",
			1806 => x"0b001924",
			1807 => x"0800180c",
			1808 => x"0000af08",
			1809 => x"00003d04",
			1810 => x"00031ce1",
			1811 => x"ffb11ce1",
			1812 => x"00111ce1",
			1813 => x"04000a04",
			1814 => x"ffce1ce1",
			1815 => x"01000504",
			1816 => x"ffdf1ce1",
			1817 => x"0200aa08",
			1818 => x"06005804",
			1819 => x"001f1ce1",
			1820 => x"007f1ce1",
			1821 => x"0e005c04",
			1822 => x"ffc81ce1",
			1823 => x"00271ce1",
			1824 => x"0e005a10",
			1825 => x"09001f04",
			1826 => x"001c1ce1",
			1827 => x"08001d04",
			1828 => x"ff7a1ce1",
			1829 => x"08001f04",
			1830 => x"00201ce1",
			1831 => x"ffeb1ce1",
			1832 => x"00291ce1",
			1833 => x"04004418",
			1834 => x"0700280c",
			1835 => x"04002508",
			1836 => x"04001904",
			1837 => x"000f1ce1",
			1838 => x"ffc11ce1",
			1839 => x"00391ce1",
			1840 => x"06007804",
			1841 => x"ff801ce1",
			1842 => x"06008604",
			1843 => x"00181ce1",
			1844 => x"ffb11ce1",
			1845 => x"05005d04",
			1846 => x"00491ce1",
			1847 => x"ffcf1ce1",
			1848 => x"0b001934",
			1849 => x"08001808",
			1850 => x"00004304",
			1851 => x"00051d85",
			1852 => x"ffac1d85",
			1853 => x"02010224",
			1854 => x"0500120c",
			1855 => x"04000d08",
			1856 => x"06001d04",
			1857 => x"00041d85",
			1858 => x"ffe31d85",
			1859 => x"00061d85",
			1860 => x"0a004510",
			1861 => x"01000508",
			1862 => x"07002904",
			1863 => x"00101d85",
			1864 => x"ffdb1d85",
			1865 => x"06008c04",
			1866 => x"00581d85",
			1867 => x"fff91d85",
			1868 => x"01000704",
			1869 => x"000a1d85",
			1870 => x"ffed1d85",
			1871 => x"01000604",
			1872 => x"00091d85",
			1873 => x"ffd61d85",
			1874 => x"0c001a08",
			1875 => x"03002e04",
			1876 => x"ffec1d85",
			1877 => x"00301d85",
			1878 => x"04004c10",
			1879 => x"09001f04",
			1880 => x"00161d85",
			1881 => x"0200ef04",
			1882 => x"ff6a1d85",
			1883 => x"0e007e04",
			1884 => x"00101d85",
			1885 => x"fff91d85",
			1886 => x"0200c904",
			1887 => x"00221d85",
			1888 => x"fff41d85",
			1889 => x"00009f1c",
			1890 => x"05002d0c",
			1891 => x"0c001408",
			1892 => x"08001604",
			1893 => x"ffe11e49",
			1894 => x"004a1e49",
			1895 => x"ffb21e49",
			1896 => x"0d001304",
			1897 => x"00001e49",
			1898 => x"0e004908",
			1899 => x"06004404",
			1900 => x"001b1e49",
			1901 => x"ffee1e49",
			1902 => x"00871e49",
			1903 => x"0e005a14",
			1904 => x"03003d0c",
			1905 => x"0e005308",
			1906 => x"06005804",
			1907 => x"fff01e49",
			1908 => x"00311e49",
			1909 => x"ff701e49",
			1910 => x"08001b04",
			1911 => x"fffa1e49",
			1912 => x"000c1e49",
			1913 => x"0200bb10",
			1914 => x"08001908",
			1915 => x"0b001604",
			1916 => x"000e1e49",
			1917 => x"ffe51e49",
			1918 => x"03002f04",
			1919 => x"00081e49",
			1920 => x"007d1e49",
			1921 => x"07002c18",
			1922 => x"04001f08",
			1923 => x"04001804",
			1924 => x"000d1e49",
			1925 => x"ffc01e49",
			1926 => x"05003f08",
			1927 => x"0c001404",
			1928 => x"fff51e49",
			1929 => x"005c1e49",
			1930 => x"0c001904",
			1931 => x"ffdc1e49",
			1932 => x"00101e49",
			1933 => x"04004704",
			1934 => x"ff851e49",
			1935 => x"03004904",
			1936 => x"002c1e49",
			1937 => x"ffe81e49",
			1938 => x"0600863c",
			1939 => x"0e006b30",
			1940 => x"0000d224",
			1941 => x"0c001104",
			1942 => x"00f71ed5",
			1943 => x"0e004d10",
			1944 => x"08001d08",
			1945 => x"01000b04",
			1946 => x"fef41ed5",
			1947 => x"003a1ed5",
			1948 => x"0c001a04",
			1949 => x"01071ed5",
			1950 => x"ff821ed5",
			1951 => x"0000b208",
			1952 => x"04002604",
			1953 => x"ff991ed5",
			1954 => x"00831ed5",
			1955 => x"06006604",
			1956 => x"feb31ed5",
			1957 => x"00101ed5",
			1958 => x"0e006904",
			1959 => x"febc1ed5",
			1960 => x"0200d704",
			1961 => x"ff701ed5",
			1962 => x"002f1ed5",
			1963 => x"05002204",
			1964 => x"ff121ed5",
			1965 => x"07003104",
			1966 => x"013b1ed5",
			1967 => x"ffbe1ed5",
			1968 => x"01000808",
			1969 => x"0b001604",
			1970 => x"ff221ed5",
			1971 => x"009c1ed5",
			1972 => x"febd1ed5",
			1973 => x"04004738",
			1974 => x"0201022c",
			1975 => x"0000fa24",
			1976 => x"01000504",
			1977 => x"fe931f51",
			1978 => x"0c001510",
			1979 => x"08001b08",
			1980 => x"0c001104",
			1981 => x"01001f51",
			1982 => x"fec51f51",
			1983 => x"0d001304",
			1984 => x"00a31f51",
			1985 => x"01601f51",
			1986 => x"05002908",
			1987 => x"00009304",
			1988 => x"ff8d1f51",
			1989 => x"fe7f1f51",
			1990 => x"03003504",
			1991 => x"003b1f51",
			1992 => x"ff9c1f51",
			1993 => x"06008f04",
			1994 => x"014c1f51",
			1995 => x"ffa41f51",
			1996 => x"01000608",
			1997 => x"0b001504",
			1998 => x"ff591f51",
			1999 => x"007b1f51",
			2000 => x"fe8c1f51",
			2001 => x"03004904",
			2002 => x"01491f51",
			2003 => x"ff141f51",
			2004 => x"06008d38",
			2005 => x"0c001b28",
			2006 => x"01000508",
			2007 => x"0e006804",
			2008 => x"fe581fc5",
			2009 => x"01581fc5",
			2010 => x"0a00451c",
			2011 => x"0c00150c",
			2012 => x"08001804",
			2013 => x"00101fc5",
			2014 => x"08001b04",
			2015 => x"01131fc5",
			2016 => x"01cb1fc5",
			2017 => x"04001f08",
			2018 => x"01000c04",
			2019 => x"fe471fc5",
			2020 => x"00521fc5",
			2021 => x"01000804",
			2022 => x"016e1fc5",
			2023 => x"00a41fc5",
			2024 => x"fe6c1fc5",
			2025 => x"05004704",
			2026 => x"fe511fc5",
			2027 => x"0000c808",
			2028 => x"0e005f04",
			2029 => x"00271fc5",
			2030 => x"01ad1fc5",
			2031 => x"fe6e1fc5",
			2032 => x"fe661fc5",
			2033 => x"0700302c",
			2034 => x"06008d28",
			2035 => x"00002504",
			2036 => x"fe622021",
			2037 => x"0800180c",
			2038 => x"06002604",
			2039 => x"00822021",
			2040 => x"0d001304",
			2041 => x"fe522021",
			2042 => x"ffe62021",
			2043 => x"0c00150c",
			2044 => x"01000904",
			2045 => x"015c2021",
			2046 => x"03001f04",
			2047 => x"01e62021",
			2048 => x"02882021",
			2049 => x"05002504",
			2050 => x"fe5b2021",
			2051 => x"0e006904",
			2052 => x"00da2021",
			2053 => x"02562021",
			2054 => x"fe602021",
			2055 => x"fe5f2021",
			2056 => x"0200a840",
			2057 => x"06005a30",
			2058 => x"0d001518",
			2059 => x"0b001208",
			2060 => x"00005204",
			2061 => x"00462105",
			2062 => x"ffed2105",
			2063 => x"0b001808",
			2064 => x"01000d04",
			2065 => x"ff922105",
			2066 => x"00152105",
			2067 => x"0b001904",
			2068 => x"002c2105",
			2069 => x"ffe82105",
			2070 => x"08001b08",
			2071 => x"07002604",
			2072 => x"ffe62105",
			2073 => x"00012105",
			2074 => x"0b001a0c",
			2075 => x"04001a08",
			2076 => x"00003504",
			2077 => x"00022105",
			2078 => x"fff92105",
			2079 => x"00652105",
			2080 => x"fff12105",
			2081 => x"0f006c0c",
			2082 => x"0c001b08",
			2083 => x"04002604",
			2084 => x"fff32105",
			2085 => x"009f2105",
			2086 => x"ffe82105",
			2087 => x"ffeb2105",
			2088 => x"0400250c",
			2089 => x"04001808",
			2090 => x"0f008a04",
			2091 => x"00182105",
			2092 => x"fff32105",
			2093 => x"ff922105",
			2094 => x"06006b10",
			2095 => x"0e005f08",
			2096 => x"0d001704",
			2097 => x"ff912105",
			2098 => x"00022105",
			2099 => x"0e006104",
			2100 => x"00042105",
			2101 => x"fffe2105",
			2102 => x"0000d004",
			2103 => x"00702105",
			2104 => x"07002c08",
			2105 => x"02010204",
			2106 => x"004b2105",
			2107 => x"ffeb2105",
			2108 => x"05005c04",
			2109 => x"ff972105",
			2110 => x"03004904",
			2111 => x"00192105",
			2112 => x"ffe82105",
			2113 => x"0000be4c",
			2114 => x"0e004e30",
			2115 => x"00008320",
			2116 => x"09001e14",
			2117 => x"0500120c",
			2118 => x"04000604",
			2119 => x"001821f9",
			2120 => x"04000b04",
			2121 => x"ffd021f9",
			2122 => x"ffff21f9",
			2123 => x"08001804",
			2124 => x"fffe21f9",
			2125 => x"006f21f9",
			2126 => x"01001408",
			2127 => x"0d001304",
			2128 => x"000221f9",
			2129 => x"ffce21f9",
			2130 => x"000521f9",
			2131 => x"01000b08",
			2132 => x"08001904",
			2133 => x"000121f9",
			2134 => x"ff8121f9",
			2135 => x"08002004",
			2136 => x"fffe21f9",
			2137 => x"001421f9",
			2138 => x"08002318",
			2139 => x"01000708",
			2140 => x"0000a604",
			2141 => x"004521f9",
			2142 => x"ff9d21f9",
			2143 => x"08001904",
			2144 => x"ffe921f9",
			2145 => x"0a002a04",
			2146 => x"000721f9",
			2147 => x"0b001904",
			2148 => x"00a521f9",
			2149 => x"001e21f9",
			2150 => x"ffcc21f9",
			2151 => x"06007514",
			2152 => x"08001f08",
			2153 => x"04004904",
			2154 => x"ff7321f9",
			2155 => x"000121f9",
			2156 => x"06007008",
			2157 => x"06006e04",
			2158 => x"fff921f9",
			2159 => x"003e21f9",
			2160 => x"ffe721f9",
			2161 => x"06008610",
			2162 => x"07002c04",
			2163 => x"005721f9",
			2164 => x"04004704",
			2165 => x"ffa721f9",
			2166 => x"0f008104",
			2167 => x"004121f9",
			2168 => x"fffb21f9",
			2169 => x"01000808",
			2170 => x"01000504",
			2171 => x"ffe721f9",
			2172 => x"001421f9",
			2173 => x"ff9e21f9",
			2174 => x"0200a834",
			2175 => x"0e005224",
			2176 => x"00009e20",
			2177 => x"05001210",
			2178 => x"04000504",
			2179 => x"001422dd",
			2180 => x"04000d04",
			2181 => x"ffc122dd",
			2182 => x"01000904",
			2183 => x"fff922dd",
			2184 => x"000722dd",
			2185 => x"0c001b0c",
			2186 => x"08001604",
			2187 => x"ffde22dd",
			2188 => x"0b001704",
			2189 => x"005f22dd",
			2190 => x"000722dd",
			2191 => x"ffd922dd",
			2192 => x"ffb022dd",
			2193 => x"0f006c0c",
			2194 => x"07002b08",
			2195 => x"09001e04",
			2196 => x"fff922dd",
			2197 => x"008b22dd",
			2198 => x"ffe922dd",
			2199 => x"ffed22dd",
			2200 => x"0e006518",
			2201 => x"0d001508",
			2202 => x"0e006104",
			2203 => x"ff8322dd",
			2204 => x"fffc22dd",
			2205 => x"04002504",
			2206 => x"ffca22dd",
			2207 => x"0d001804",
			2208 => x"004322dd",
			2209 => x"0e005c04",
			2210 => x"000322dd",
			2211 => x"ffd722dd",
			2212 => x"0f008910",
			2213 => x"0a004304",
			2214 => x"005922dd",
			2215 => x"04004704",
			2216 => x"ffd622dd",
			2217 => x"0f007804",
			2218 => x"fff722dd",
			2219 => x"002122dd",
			2220 => x"0100080c",
			2221 => x"03003508",
			2222 => x"05003604",
			2223 => x"ffea22dd",
			2224 => x"005b22dd",
			2225 => x"ffd822dd",
			2226 => x"05004a04",
			2227 => x"ff8822dd",
			2228 => x"04003804",
			2229 => x"001522dd",
			2230 => x"fff822dd",
			2231 => x"0d001320",
			2232 => x"00008814",
			2233 => x"05001208",
			2234 => x"02002904",
			2235 => x"001223c1",
			2236 => x"ffc823c1",
			2237 => x"01000c08",
			2238 => x"0b001404",
			2239 => x"005123c1",
			2240 => x"000623c1",
			2241 => x"000023c1",
			2242 => x"06008c04",
			2243 => x"ff7623c1",
			2244 => x"00010e04",
			2245 => x"002d23c1",
			2246 => x"ffec23c1",
			2247 => x"04003e40",
			2248 => x"0000ae20",
			2249 => x"0e005118",
			2250 => x"0b001608",
			2251 => x"01000904",
			2252 => x"ffff23c1",
			2253 => x"004323c1",
			2254 => x"01001008",
			2255 => x"07002004",
			2256 => x"000823c1",
			2257 => x"ff9f23c1",
			2258 => x"0d001b04",
			2259 => x"001623c1",
			2260 => x"fff723c1",
			2261 => x"05003504",
			2262 => x"ffd023c1",
			2263 => x"008623c1",
			2264 => x"0a002c0c",
			2265 => x"05002808",
			2266 => x"0d001504",
			2267 => x"001723c1",
			2268 => x"ffc223c1",
			2269 => x"005323c1",
			2270 => x"0e006804",
			2271 => x"ff8023c1",
			2272 => x"01000908",
			2273 => x"05003804",
			2274 => x"fff623c1",
			2275 => x"004e23c1",
			2276 => x"05004a04",
			2277 => x"ffc423c1",
			2278 => x"000c23c1",
			2279 => x"0a004808",
			2280 => x"0d001504",
			2281 => x"000d23c1",
			2282 => x"008f23c1",
			2283 => x"04004d04",
			2284 => x"ffd623c1",
			2285 => x"08001f04",
			2286 => x"000723c1",
			2287 => x"fffb23c1",
			2288 => x"0200aa40",
			2289 => x"0e00522c",
			2290 => x"0b00171c",
			2291 => x"01000910",
			2292 => x"09001e0c",
			2293 => x"00006508",
			2294 => x"0c001404",
			2295 => x"004e24ad",
			2296 => x"ffd524ad",
			2297 => x"ff0d24ad",
			2298 => x"001424ad",
			2299 => x"00008608",
			2300 => x"04001204",
			2301 => x"003324ad",
			2302 => x"010224ad",
			2303 => x"ffdb24ad",
			2304 => x"01001004",
			2305 => x"ff0024ad",
			2306 => x"08002408",
			2307 => x"08002004",
			2308 => x"fffc24ad",
			2309 => x"005d24ad",
			2310 => x"ffe024ad",
			2311 => x"0500470c",
			2312 => x"0f006604",
			2313 => x"00d924ad",
			2314 => x"01000904",
			2315 => x"ff3124ad",
			2316 => x"005924ad",
			2317 => x"0a004304",
			2318 => x"010d24ad",
			2319 => x"ffe324ad",
			2320 => x"0600660c",
			2321 => x"09002304",
			2322 => x"fef224ad",
			2323 => x"0c002104",
			2324 => x"002624ad",
			2325 => x"fffb24ad",
			2326 => x"04002510",
			2327 => x"09001c04",
			2328 => x"fee324ad",
			2329 => x"03002404",
			2330 => x"00d224ad",
			2331 => x"04001b04",
			2332 => x"004724ad",
			2333 => x"ff1b24ad",
			2334 => x"0000c004",
			2335 => x"00c824ad",
			2336 => x"09001d08",
			2337 => x"0a003704",
			2338 => x"00f224ad",
			2339 => x"ffaf24ad",
			2340 => x"08001908",
			2341 => x"0e006304",
			2342 => x"ffa324ad",
			2343 => x"00a424ad",
			2344 => x"0e006804",
			2345 => x"ff1c24ad",
			2346 => x"000124ad",
			2347 => x"06008d3c",
			2348 => x"0d00192c",
			2349 => x"0000fa28",
			2350 => x"01000508",
			2351 => x"0a004504",
			2352 => x"fe542529",
			2353 => x"00fb2529",
			2354 => x"0000c710",
			2355 => x"0e005a08",
			2356 => x"0000ae04",
			2357 => x"00a02529",
			2358 => x"fdd92529",
			2359 => x"05002204",
			2360 => x"ff0c2529",
			2361 => x"01852529",
			2362 => x"09001f08",
			2363 => x"09001c04",
			2364 => x"fee32529",
			2365 => x"01782529",
			2366 => x"04004c04",
			2367 => x"fe982529",
			2368 => x"01ad2529",
			2369 => x"01ed2529",
			2370 => x"07002908",
			2371 => x"06004504",
			2372 => x"feb52529",
			2373 => x"018d2529",
			2374 => x"07002b04",
			2375 => x"fda02529",
			2376 => x"fe6c2529",
			2377 => x"fe682529",
			2378 => x"0d00153c",
			2379 => x"0300352c",
			2380 => x"04003428",
			2381 => x"0b001410",
			2382 => x"04000c04",
			2383 => x"ffcc261d",
			2384 => x"08001604",
			2385 => x"ffc6261d",
			2386 => x"0e007104",
			2387 => x"009b261d",
			2388 => x"ffe0261d",
			2389 => x"0c001508",
			2390 => x"0000d304",
			2391 => x"003e261d",
			2392 => x"ffe2261d",
			2393 => x"05003808",
			2394 => x"01000e04",
			2395 => x"ff38261d",
			2396 => x"000f261d",
			2397 => x"04002d04",
			2398 => x"006d261d",
			2399 => x"ff9a261d",
			2400 => x"008d261d",
			2401 => x"09002108",
			2402 => x"0b001804",
			2403 => x"ff12261d",
			2404 => x"000c261d",
			2405 => x"0c001b04",
			2406 => x"0063261d",
			2407 => x"ffba261d",
			2408 => x"0700291c",
			2409 => x"0c001a0c",
			2410 => x"05002808",
			2411 => x"07002204",
			2412 => x"0014261d",
			2413 => x"ffd9261d",
			2414 => x"00e2261d",
			2415 => x"0000a90c",
			2416 => x"09002104",
			2417 => x"ff78261d",
			2418 => x"09002204",
			2419 => x"0006261d",
			2420 => x"fff7261d",
			2421 => x"004c261d",
			2422 => x"04003e14",
			2423 => x"0f008e0c",
			2424 => x"0f006c08",
			2425 => x"0e005604",
			2426 => x"ffc5261d",
			2427 => x"0039261d",
			2428 => x"ff55261d",
			2429 => x"07002e04",
			2430 => x"0069261d",
			2431 => x"ffc9261d",
			2432 => x"0a004804",
			2433 => x"008b261d",
			2434 => x"04004d04",
			2435 => x"ffbb261d",
			2436 => x"04005a04",
			2437 => x"0008261d",
			2438 => x"fff8261d",
			2439 => x"06008d54",
			2440 => x"0e00652c",
			2441 => x"0200b720",
			2442 => x"0e005a14",
			2443 => x"0000ae0c",
			2444 => x"0a003e08",
			2445 => x"05001204",
			2446 => x"feb826c9",
			2447 => x"005926c9",
			2448 => x"ff2426c9",
			2449 => x"0a003e04",
			2450 => x"fe1926c9",
			2451 => x"002f26c9",
			2452 => x"04003604",
			2453 => x"ffcc26c9",
			2454 => x"01000904",
			2455 => x"008926c9",
			2456 => x"01cd26c9",
			2457 => x"07002c04",
			2458 => x"fe3526c9",
			2459 => x"0a004504",
			2460 => x"004e26c9",
			2461 => x"fea926c9",
			2462 => x"08001f18",
			2463 => x"08001c10",
			2464 => x"04002108",
			2465 => x"0200a904",
			2466 => x"000526c9",
			2467 => x"fe6d26c9",
			2468 => x"09002004",
			2469 => x"016f26c9",
			2470 => x"ffe826c9",
			2471 => x"07003404",
			2472 => x"01d726c9",
			2473 => x"ff8d26c9",
			2474 => x"0f00890c",
			2475 => x"08002208",
			2476 => x"0200d504",
			2477 => x"018526c9",
			2478 => x"ffa126c9",
			2479 => x"feed26c9",
			2480 => x"fe3c26c9",
			2481 => x"fe7526c9",
			2482 => x"0000ae3c",
			2483 => x"0e00522c",
			2484 => x"0b001208",
			2485 => x"00004904",
			2486 => x"007027ad",
			2487 => x"fff327ad",
			2488 => x"01000b10",
			2489 => x"0400340c",
			2490 => x"08001d04",
			2491 => x"ff5627ad",
			2492 => x"08001f04",
			2493 => x"ffed27ad",
			2494 => x"001127ad",
			2495 => x"ffee27ad",
			2496 => x"0400170c",
			2497 => x"05001804",
			2498 => x"ffd727ad",
			2499 => x"05001b04",
			2500 => x"000627ad",
			2501 => x"fffb27ad",
			2502 => x"0c001b04",
			2503 => x"008427ad",
			2504 => x"ffe727ad",
			2505 => x"0f006c0c",
			2506 => x"0a004008",
			2507 => x"07002704",
			2508 => x"002627ad",
			2509 => x"00cb27ad",
			2510 => x"000327ad",
			2511 => x"ffd927ad",
			2512 => x"0e00651c",
			2513 => x"04004414",
			2514 => x"01001210",
			2515 => x"08001604",
			2516 => x"002327ad",
			2517 => x"07002d08",
			2518 => x"0c001b04",
			2519 => x"ff3a27ad",
			2520 => x"ffe527ad",
			2521 => x"001327ad",
			2522 => x"002d27ad",
			2523 => x"07002f04",
			2524 => x"004027ad",
			2525 => x"ffe227ad",
			2526 => x"02010218",
			2527 => x"07002c08",
			2528 => x"05002804",
			2529 => x"ffd327ad",
			2530 => x"009d27ad",
			2531 => x"0200cc0c",
			2532 => x"05005008",
			2533 => x"0f009204",
			2534 => x"ffb527ad",
			2535 => x"002227ad",
			2536 => x"008827ad",
			2537 => x"ff6f27ad",
			2538 => x"ff8927ad",
			2539 => x"02009730",
			2540 => x"0e004820",
			2541 => x"07001704",
			2542 => x"004b2899",
			2543 => x"08001d10",
			2544 => x"01000a04",
			2545 => x"ff7e2899",
			2546 => x"01000c08",
			2547 => x"01000b04",
			2548 => x"00012899",
			2549 => x"00112899",
			2550 => x"ffe12899",
			2551 => x"05001e04",
			2552 => x"ffe42899",
			2553 => x"0c001a04",
			2554 => x"00462899",
			2555 => x"fffa2899",
			2556 => x"0100120c",
			2557 => x"08001904",
			2558 => x"000e2899",
			2559 => x"07002504",
			2560 => x"00002899",
			2561 => x"00a52899",
			2562 => x"fff12899",
			2563 => x"0e005a14",
			2564 => x"0d00150c",
			2565 => x"03003508",
			2566 => x"01000704",
			2567 => x"00162899",
			2568 => x"ffdf2899",
			2569 => x"ff762899",
			2570 => x"03003a04",
			2571 => x"ffc42899",
			2572 => x"00372899",
			2573 => x"0200b70c",
			2574 => x"08001904",
			2575 => x"ffe82899",
			2576 => x"0f007504",
			2577 => x"00912899",
			2578 => x"000b2899",
			2579 => x"0700290c",
			2580 => x"0a002804",
			2581 => x"ffba2899",
			2582 => x"0a003404",
			2583 => x"00742899",
			2584 => x"00032899",
			2585 => x"01000610",
			2586 => x"0200d908",
			2587 => x"06007104",
			2588 => x"ffde2899",
			2589 => x"005c2899",
			2590 => x"03003304",
			2591 => x"00162899",
			2592 => x"ffae2899",
			2593 => x"0e006904",
			2594 => x"ff582899",
			2595 => x"06008604",
			2596 => x"00652899",
			2597 => x"ff892899",
			2598 => x"00008320",
			2599 => x"05001208",
			2600 => x"07001704",
			2601 => x"002f298d",
			2602 => x"ff75298d",
			2603 => x"09001e0c",
			2604 => x"0c001908",
			2605 => x"08001904",
			2606 => x"0021298d",
			2607 => x"00dd298d",
			2608 => x"ffe7298d",
			2609 => x"01001404",
			2610 => x"ff92298d",
			2611 => x"08002604",
			2612 => x"002e298d",
			2613 => x"fff7298d",
			2614 => x"0400251c",
			2615 => x"0e00650c",
			2616 => x"00009608",
			2617 => x"06004f04",
			2618 => x"ffcb298d",
			2619 => x"0036298d",
			2620 => x"fefc298d",
			2621 => x"0f008b04",
			2622 => x"00a2298d",
			2623 => x"0c001704",
			2624 => x"ff22298d",
			2625 => x"03002404",
			2626 => x"0066298d",
			2627 => x"ffca298d",
			2628 => x"0d001524",
			2629 => x"03003510",
			2630 => x"01000a0c",
			2631 => x"07002504",
			2632 => x"ffdf298d",
			2633 => x"0e007204",
			2634 => x"00b6298d",
			2635 => x"fff6298d",
			2636 => x"ff70298d",
			2637 => x"0b001808",
			2638 => x"07002b04",
			2639 => x"fef9298d",
			2640 => x"ffef298d",
			2641 => x"01000704",
			2642 => x"ff63298d",
			2643 => x"04004004",
			2644 => x"00b7298d",
			2645 => x"ffdb298d",
			2646 => x"0c001a08",
			2647 => x"06007104",
			2648 => x"010d298d",
			2649 => x"fffe298d",
			2650 => x"0b001904",
			2651 => x"0078298d",
			2652 => x"0a003b08",
			2653 => x"0a003704",
			2654 => x"ffbb298d",
			2655 => x"007c298d",
			2656 => x"08001d04",
			2657 => x"fefc298d",
			2658 => x"000c298d",
			2659 => x"07002c58",
			2660 => x"04001714",
			2661 => x"0c00130c",
			2662 => x"00009408",
			2663 => x"08001904",
			2664 => x"031d2a69",
			2665 => x"05122a69",
			2666 => x"fe5d2a69",
			2667 => x"0c001404",
			2668 => x"ff7a2a69",
			2669 => x"fe4c2a69",
			2670 => x"08001b18",
			2671 => x"05003808",
			2672 => x"07001f04",
			2673 => x"ff692a69",
			2674 => x"fe4b2a69",
			2675 => x"03003508",
			2676 => x"07002504",
			2677 => x"ff5d2a69",
			2678 => x"06f82a69",
			2679 => x"0d001404",
			2680 => x"fe482a69",
			2681 => x"00ff2a69",
			2682 => x"0000b51c",
			2683 => x"0b00160c",
			2684 => x"04002b08",
			2685 => x"0e004204",
			2686 => x"05162a69",
			2687 => x"07442a69",
			2688 => x"02672a69",
			2689 => x"05003808",
			2690 => x"09002004",
			2691 => x"00a82a69",
			2692 => x"fe342a69",
			2693 => x"0e005a04",
			2694 => x"03cf2a69",
			2695 => x"06642a69",
			2696 => x"0e005b04",
			2697 => x"fe412a69",
			2698 => x"0d001304",
			2699 => x"ff222a69",
			2700 => x"0a003604",
			2701 => x"02b02a69",
			2702 => x"06272a69",
			2703 => x"07002f14",
			2704 => x"05004e0c",
			2705 => x"04002204",
			2706 => x"fe4e2a69",
			2707 => x"0b001604",
			2708 => x"ffb82a69",
			2709 => x"fe4d2a69",
			2710 => x"03004504",
			2711 => x"064d2a69",
			2712 => x"ffe92a69",
			2713 => x"fe4c2a69",
			2714 => x"0c00140c",
			2715 => x"08001604",
			2716 => x"ffdc2b35",
			2717 => x"0000c504",
			2718 => x"00872b35",
			2719 => x"ffdf2b35",
			2720 => x"04003434",
			2721 => x"01000b14",
			2722 => x"08001c04",
			2723 => x"ff742b35",
			2724 => x"00006e04",
			2725 => x"00152b35",
			2726 => x"00010c08",
			2727 => x"0e006604",
			2728 => x"ffc92b35",
			2729 => x"fffd2b35",
			2730 => x"00102b35",
			2731 => x"0b001614",
			2732 => x"05002808",
			2733 => x"03002604",
			2734 => x"ffca2b35",
			2735 => x"00052b35",
			2736 => x"0a002c04",
			2737 => x"00872b35",
			2738 => x"03002a04",
			2739 => x"ffe82b35",
			2740 => x"00092b35",
			2741 => x"05003504",
			2742 => x"ffa12b35",
			2743 => x"0e005b04",
			2744 => x"00312b35",
			2745 => x"ffe62b35",
			2746 => x"0a00451c",
			2747 => x"01000708",
			2748 => x"05004b04",
			2749 => x"001b2b35",
			2750 => x"ffc72b35",
			2751 => x"01000804",
			2752 => x"007f2b35",
			2753 => x"09002108",
			2754 => x"04003b04",
			2755 => x"00152b35",
			2756 => x"ff9a2b35",
			2757 => x"0000d004",
			2758 => x"00862b35",
			2759 => x"ffdf2b35",
			2760 => x"07002e04",
			2761 => x"ffaf2b35",
			2762 => x"09002504",
			2763 => x"002f2b35",
			2764 => x"ffe42b35",
			2765 => x"04003454",
			2766 => x"0b00173c",
			2767 => x"0000941c",
			2768 => x"01000910",
			2769 => x"05001204",
			2770 => x"fe492c19",
			2771 => x"03001804",
			2772 => x"01432c19",
			2773 => x"08001804",
			2774 => x"fec22c19",
			2775 => x"000d2c19",
			2776 => x"05001804",
			2777 => x"00d02c19",
			2778 => x"03002904",
			2779 => x"01882c19",
			2780 => x"00c32c19",
			2781 => x"0d001618",
			2782 => x"01000c10",
			2783 => x"05003808",
			2784 => x"0c001504",
			2785 => x"ffc12c19",
			2786 => x"fe5b2c19",
			2787 => x"05003f04",
			2788 => x"01202c19",
			2789 => x"ff1d2c19",
			2790 => x"0a002c04",
			2791 => x"019f2c19",
			2792 => x"fef72c19",
			2793 => x"03002c04",
			2794 => x"fe542c19",
			2795 => x"00be2c19",
			2796 => x"0100080c",
			2797 => x"09002008",
			2798 => x"06005504",
			2799 => x"fefa2c19",
			2800 => x"01202c19",
			2801 => x"fe982c19",
			2802 => x"01001404",
			2803 => x"fe4d2c19",
			2804 => x"08002404",
			2805 => x"00c92c19",
			2806 => x"fea32c19",
			2807 => x"03003504",
			2808 => x"00fb2c19",
			2809 => x"0d001304",
			2810 => x"fe662c19",
			2811 => x"0e005604",
			2812 => x"ff9b2c19",
			2813 => x"08001b08",
			2814 => x"01000704",
			2815 => x"fe6f2c19",
			2816 => x"00962c19",
			2817 => x"07002f08",
			2818 => x"0000b504",
			2819 => x"01b52c19",
			2820 => x"00ab2c19",
			2821 => x"febd2c19",
			2822 => x"08001808",
			2823 => x"00003504",
			2824 => x"00382cdd",
			2825 => x"ff6b2cdd",
			2826 => x"00009e28",
			2827 => x"0e00481c",
			2828 => x"0c001608",
			2829 => x"05001204",
			2830 => x"ffb82cdd",
			2831 => x"008f2cdd",
			2832 => x"08001d08",
			2833 => x"01000b04",
			2834 => x"ff582cdd",
			2835 => x"00012cdd",
			2836 => x"07002408",
			2837 => x"07001f04",
			2838 => x"fff92cdd",
			2839 => x"00272cdd",
			2840 => x"ffe32cdd",
			2841 => x"0c001808",
			2842 => x"04002004",
			2843 => x"006e2cdd",
			2844 => x"ffad2cdd",
			2845 => x"00e62cdd",
			2846 => x"0e005710",
			2847 => x"08001b04",
			2848 => x"002b2cdd",
			2849 => x"08001d04",
			2850 => x"ff372cdd",
			2851 => x"08001f04",
			2852 => x"002a2cdd",
			2853 => x"ffc72cdd",
			2854 => x"0000b208",
			2855 => x"0f006c04",
			2856 => x"00d22cdd",
			2857 => x"000b2cdd",
			2858 => x"0e00610c",
			2859 => x"0d001504",
			2860 => x"ff312cdd",
			2861 => x"04003f04",
			2862 => x"003c2cdd",
			2863 => x"ffb32cdd",
			2864 => x"04003c08",
			2865 => x"09001f04",
			2866 => x"00262cdd",
			2867 => x"ff722cdd",
			2868 => x"0000d004",
			2869 => x"00bb2cdd",
			2870 => x"ffdb2cdd",
			2871 => x"0c00140c",
			2872 => x"08001604",
			2873 => x"ffdb2db9",
			2874 => x"0000c504",
			2875 => x"008c2db9",
			2876 => x"ffdf2db9",
			2877 => x"04003438",
			2878 => x"01000b18",
			2879 => x"08002014",
			2880 => x"0e007008",
			2881 => x"0d001704",
			2882 => x"ff712db9",
			2883 => x"00052db9",
			2884 => x"0d001304",
			2885 => x"ffdc2db9",
			2886 => x"0f00a704",
			2887 => x"00242db9",
			2888 => x"fff32db9",
			2889 => x"00082db9",
			2890 => x"0b001614",
			2891 => x"05002808",
			2892 => x"03002604",
			2893 => x"ffc72db9",
			2894 => x"00052db9",
			2895 => x"0a002c04",
			2896 => x"008b2db9",
			2897 => x"03002a04",
			2898 => x"ffe72db9",
			2899 => x"00092db9",
			2900 => x"05003504",
			2901 => x"ff9e2db9",
			2902 => x"0e005b04",
			2903 => x"00322db9",
			2904 => x"ffe52db9",
			2905 => x"0a004520",
			2906 => x"0d00140c",
			2907 => x"05004904",
			2908 => x"004d2db9",
			2909 => x"08001b04",
			2910 => x"ff9d2db9",
			2911 => x"fff62db9",
			2912 => x"0000d00c",
			2913 => x"03003b08",
			2914 => x"0a003b04",
			2915 => x"00342db9",
			2916 => x"ffd32db9",
			2917 => x"00972db9",
			2918 => x"03003a04",
			2919 => x"000a2db9",
			2920 => x"ffd62db9",
			2921 => x"07002e04",
			2922 => x"ffad2db9",
			2923 => x"09002504",
			2924 => x"00312db9",
			2925 => x"ffe32db9",
			2926 => x"0000be4c",
			2927 => x"08001814",
			2928 => x"03003410",
			2929 => x"08001608",
			2930 => x"00008f04",
			2931 => x"ffb72e9d",
			2932 => x"000f2e9d",
			2933 => x"01000504",
			2934 => x"ffe62e9d",
			2935 => x"005f2e9d",
			2936 => x"ff672e9d",
			2937 => x"0e005a30",
			2938 => x"00009e20",
			2939 => x"0e004810",
			2940 => x"0c001608",
			2941 => x"04000e04",
			2942 => x"ffcf2e9d",
			2943 => x"00952e9d",
			2944 => x"08001d04",
			2945 => x"ff5c2e9d",
			2946 => x"000f2e9d",
			2947 => x"04002608",
			2948 => x"0c001604",
			2949 => x"00722e9d",
			2950 => x"ffbd2e9d",
			2951 => x"0c001804",
			2952 => x"00132e9d",
			2953 => x"00ef2e9d",
			2954 => x"03003b0c",
			2955 => x"07002808",
			2956 => x"09001e04",
			2957 => x"ff5f2e9d",
			2958 => x"00912e9d",
			2959 => x"ff172e9d",
			2960 => x"005b2e9d",
			2961 => x"04002104",
			2962 => x"ffec2e9d",
			2963 => x"00d52e9d",
			2964 => x"0e006308",
			2965 => x"01001204",
			2966 => x"ff142e9d",
			2967 => x"00322e9d",
			2968 => x"04003c18",
			2969 => x"07002c14",
			2970 => x"0100080c",
			2971 => x"03003108",
			2972 => x"07002b04",
			2973 => x"ffbf2e9d",
			2974 => x"001e2e9d",
			2975 => x"009a2e9d",
			2976 => x"07002b04",
			2977 => x"ff362e9d",
			2978 => x"007b2e9d",
			2979 => x"ff292e9d",
			2980 => x"0a004804",
			2981 => x"009a2e9d",
			2982 => x"ffc22e9d",
			2983 => x"04003460",
			2984 => x"0b00173c",
			2985 => x"0000941c",
			2986 => x"01000910",
			2987 => x"05001204",
			2988 => x"fe5c2fa1",
			2989 => x"03001804",
			2990 => x"01352fa1",
			2991 => x"08001804",
			2992 => x"fecc2fa1",
			2993 => x"000e2fa1",
			2994 => x"05001804",
			2995 => x"00bf2fa1",
			2996 => x"03002904",
			2997 => x"01812fa1",
			2998 => x"00b82fa1",
			2999 => x"0d001618",
			3000 => x"01000c10",
			3001 => x"05003808",
			3002 => x"0c001504",
			3003 => x"ffbe2fa1",
			3004 => x"fe612fa1",
			3005 => x"0000ed04",
			3006 => x"ff632fa1",
			3007 => x"01632fa1",
			3008 => x"0a002c04",
			3009 => x"01902fa1",
			3010 => x"ff042fa1",
			3011 => x"03002c04",
			3012 => x"fe612fa1",
			3013 => x"00ad2fa1",
			3014 => x"0100080c",
			3015 => x"09002008",
			3016 => x"06005504",
			3017 => x"ff052fa1",
			3018 => x"010b2fa1",
			3019 => x"fea52fa1",
			3020 => x"0100140c",
			3021 => x"07002608",
			3022 => x"07002404",
			3023 => x"feb42fa1",
			3024 => x"ffd52fa1",
			3025 => x"fe352fa1",
			3026 => x"0e005408",
			3027 => x"0d002004",
			3028 => x"00fb2fa1",
			3029 => x"ffb02fa1",
			3030 => x"feaf2fa1",
			3031 => x"04003504",
			3032 => x"013c2fa1",
			3033 => x"08001d18",
			3034 => x"01000708",
			3035 => x"0200bb04",
			3036 => x"ffb52fa1",
			3037 => x"fe722fa1",
			3038 => x"0e005604",
			3039 => x"ff532fa1",
			3040 => x"0a004508",
			3041 => x"04003e04",
			3042 => x"00842fa1",
			3043 => x"01962fa1",
			3044 => x"fea72fa1",
			3045 => x"07002f04",
			3046 => x"01472fa1",
			3047 => x"fed52fa1",
			3048 => x"09002154",
			3049 => x"05004b44",
			3050 => x"03003330",
			3051 => x"01000a10",
			3052 => x"0c001104",
			3053 => x"00ab30a5",
			3054 => x"08001d08",
			3055 => x"06008104",
			3056 => x"fed430a5",
			3057 => x"ffd930a5",
			3058 => x"007230a5",
			3059 => x"0f008010",
			3060 => x"0b001608",
			3061 => x"0d001204",
			3062 => x"ffcd30a5",
			3063 => x"00f530a5",
			3064 => x"00009e04",
			3065 => x"ff7730a5",
			3066 => x"008730a5",
			3067 => x"05002908",
			3068 => x"07002f04",
			3069 => x"fee830a5",
			3070 => x"003230a5",
			3071 => x"09001e04",
			3072 => x"007430a5",
			3073 => x"ff5230a5",
			3074 => x"0e004d04",
			3075 => x"ff1e30a5",
			3076 => x"0300390c",
			3077 => x"02010208",
			3078 => x"05004504",
			3079 => x"008230a5",
			3080 => x"014130a5",
			3081 => x"ff6730a5",
			3082 => x"ff7030a5",
			3083 => x"03004008",
			3084 => x"0e005c04",
			3085 => x"fef830a5",
			3086 => x"ffaf30a5",
			3087 => x"03004504",
			3088 => x"006b30a5",
			3089 => x"ffc930a5",
			3090 => x"05004b14",
			3091 => x"0b001804",
			3092 => x"004d30a5",
			3093 => x"07002808",
			3094 => x"00008104",
			3095 => x"ffd530a5",
			3096 => x"003d30a5",
			3097 => x"05004704",
			3098 => x"fefb30a5",
			3099 => x"ffd430a5",
			3100 => x"0200b904",
			3101 => x"012030a5",
			3102 => x"0e00680c",
			3103 => x"08001f04",
			3104 => x"ff2030a5",
			3105 => x"01000e04",
			3106 => x"fff230a5",
			3107 => x"003a30a5",
			3108 => x"0f008108",
			3109 => x"08002004",
			3110 => x"010830a5",
			3111 => x"fff930a5",
			3112 => x"ff9b30a5",
			3113 => x"0e007240",
			3114 => x"0c001e3c",
			3115 => x"05001308",
			3116 => x"07001704",
			3117 => x"00523131",
			3118 => x"fe523131",
			3119 => x"01000b1c",
			3120 => x"0e005210",
			3121 => x"0b001408",
			3122 => x"00008304",
			3123 => x"01bd3131",
			3124 => x"fe793131",
			3125 => x"01000804",
			3126 => x"00003131",
			3127 => x"fe473131",
			3128 => x"0d001708",
			3129 => x"0000b504",
			3130 => x"01093131",
			3131 => x"ffe43131",
			3132 => x"020e3131",
			3133 => x"02008f0c",
			3134 => x"0b001908",
			3135 => x"03001804",
			3136 => x"017f3131",
			3137 => x"02013131",
			3138 => x"ff663131",
			3139 => x"04002d08",
			3140 => x"0b001604",
			3141 => x"00c03131",
			3142 => x"fe073131",
			3143 => x"01623131",
			3144 => x"fe643131",
			3145 => x"0000bc04",
			3146 => x"00ad3131",
			3147 => x"fe623131",
			3148 => x"07001604",
			3149 => x"e77b31dd",
			3150 => x"0200bb3c",
			3151 => x"05002714",
			3152 => x"0c001408",
			3153 => x"08001804",
			3154 => x"d66631dd",
			3155 => x"e95431dd",
			3156 => x"0c001504",
			3157 => x"d88d31dd",
			3158 => x"04001d04",
			3159 => x"d65831dd",
			3160 => x"d78a31dd",
			3161 => x"08001c18",
			3162 => x"0d00140c",
			3163 => x"01000908",
			3164 => x"0000a604",
			3165 => x"d93b31dd",
			3166 => x"d65f31dd",
			3167 => x"dca531dd",
			3168 => x"0e005104",
			3169 => x"daad31dd",
			3170 => x"0000b404",
			3171 => x"e85b31dd",
			3172 => x"de5531dd",
			3173 => x"0c001e0c",
			3174 => x"0200ac08",
			3175 => x"0c001704",
			3176 => x"ea8631dd",
			3177 => x"e59831dd",
			3178 => x"de9531dd",
			3179 => x"d66431dd",
			3180 => x"0e007214",
			3181 => x"0f008e10",
			3182 => x"0a002c04",
			3183 => x"d93131dd",
			3184 => x"0a004808",
			3185 => x"04003d04",
			3186 => x"d65c31dd",
			3187 => x"da3831dd",
			3188 => x"d65931dd",
			3189 => x"dc2731dd",
			3190 => x"d65831dd",
			3191 => x"0000be44",
			3192 => x"01000504",
			3193 => x"ff8432b1",
			3194 => x"0e005224",
			3195 => x"00008314",
			3196 => x"0c00190c",
			3197 => x"04000a04",
			3198 => x"ffd432b1",
			3199 => x"01000704",
			3200 => x"000732b1",
			3201 => x"009832b1",
			3202 => x"01001604",
			3203 => x"ffb432b1",
			3204 => x"001432b1",
			3205 => x"01000b08",
			3206 => x"08001904",
			3207 => x"000132b1",
			3208 => x"ff4832b1",
			3209 => x"0e004804",
			3210 => x"fffa32b1",
			3211 => x"005132b1",
			3212 => x"0d001918",
			3213 => x"0200a80c",
			3214 => x"0c001a08",
			3215 => x"0d001304",
			3216 => x"001c32b1",
			3217 => x"00f732b1",
			3218 => x"fff132b1",
			3219 => x"06006504",
			3220 => x"ff6232b1",
			3221 => x"0b001604",
			3222 => x"ffeb32b1",
			3223 => x"008a32b1",
			3224 => x"ffa332b1",
			3225 => x"0e006304",
			3226 => x"ff1d32b1",
			3227 => x"06007910",
			3228 => x"0a004304",
			3229 => x"008f32b1",
			3230 => x"05005b04",
			3231 => x"ff8432b1",
			3232 => x"0f007804",
			3233 => x"ffe332b1",
			3234 => x"005e32b1",
			3235 => x"07002c10",
			3236 => x"04001f04",
			3237 => x"ff9f32b1",
			3238 => x"02010204",
			3239 => x"006832b1",
			3240 => x"07002b04",
			3241 => x"ffad32b1",
			3242 => x"001832b1",
			3243 => x"ff5932b1",
			3244 => x"00009e30",
			3245 => x"08001604",
			3246 => x"ff5a33a5",
			3247 => x"04003628",
			3248 => x"0c00160c",
			3249 => x"01000908",
			3250 => x"00006504",
			3251 => x"006833a5",
			3252 => x"ff6633a5",
			3253 => x"00df33a5",
			3254 => x"01000b0c",
			3255 => x"00009408",
			3256 => x"07002704",
			3257 => x"ff2933a5",
			3258 => x"001c33a5",
			3259 => x"002133a5",
			3260 => x"07002908",
			3261 => x"0c001b04",
			3262 => x"00bd33a5",
			3263 => x"ffd233a5",
			3264 => x"08001f04",
			3265 => x"000533a5",
			3266 => x"ff8733a5",
			3267 => x"00d633a5",
			3268 => x"0e005718",
			3269 => x"0100090c",
			3270 => x"04003308",
			3271 => x"04002104",
			3272 => x"fff233a5",
			3273 => x"006533a5",
			3274 => x"ff8e33a5",
			3275 => x"0d001704",
			3276 => x"fee833a5",
			3277 => x"0d001a04",
			3278 => x"002c33a5",
			3279 => x"ffae33a5",
			3280 => x"0000b20c",
			3281 => x"01000904",
			3282 => x"ffda33a5",
			3283 => x"03003a04",
			3284 => x"00fa33a5",
			3285 => x"002733a5",
			3286 => x"0d00130c",
			3287 => x"06008c04",
			3288 => x"ff0133a5",
			3289 => x"00010e04",
			3290 => x"007e33a5",
			3291 => x"ffb333a5",
			3292 => x"06006b0c",
			3293 => x"0d001704",
			3294 => x"ff2833a5",
			3295 => x"05005804",
			3296 => x"007133a5",
			3297 => x"ff9f33a5",
			3298 => x"06007008",
			3299 => x"0200c304",
			3300 => x"010333a5",
			3301 => x"ffca33a5",
			3302 => x"06007504",
			3303 => x"ff2b33a5",
			3304 => x"002633a5",
			3305 => x"0500485c",
			3306 => x"0b001738",
			3307 => x"02008e18",
			3308 => x"0d001310",
			3309 => x"0c001104",
			3310 => x"010d34a9",
			3311 => x"08001904",
			3312 => x"feb834a9",
			3313 => x"0c001404",
			3314 => x"00e334a9",
			3315 => x"ff9a34a9",
			3316 => x"06003804",
			3317 => x"003634a9",
			3318 => x"012834a9",
			3319 => x"0e006508",
			3320 => x"04002d04",
			3321 => x"fe9534a9",
			3322 => x"ffee34a9",
			3323 => x"08001b08",
			3324 => x"03003104",
			3325 => x"febd34a9",
			3326 => x"004934a9",
			3327 => x"08001f08",
			3328 => x"06008e04",
			3329 => x"014634a9",
			3330 => x"ff6334a9",
			3331 => x"08002004",
			3332 => x"fee034a9",
			3333 => x"009a34a9",
			3334 => x"00009e18",
			3335 => x"0e004e14",
			3336 => x"09001e08",
			3337 => x"0b001804",
			3338 => x"ff9d34a9",
			3339 => x"00c234a9",
			3340 => x"01001004",
			3341 => x"fe9434a9",
			3342 => x"0d001c04",
			3343 => x"005f34a9",
			3344 => x"ffc534a9",
			3345 => x"00fe34a9",
			3346 => x"07002604",
			3347 => x"005734a9",
			3348 => x"05004604",
			3349 => x"fe9134a9",
			3350 => x"ffa034a9",
			3351 => x"0e005204",
			3352 => x"ff2634a9",
			3353 => x"05004904",
			3354 => x"015b34a9",
			3355 => x"08001b0c",
			3356 => x"0d001508",
			3357 => x"0b001804",
			3358 => x"fe9834a9",
			3359 => x"ffb234a9",
			3360 => x"005934a9",
			3361 => x"04003908",
			3362 => x"03003a04",
			3363 => x"004c34a9",
			3364 => x"fef534a9",
			3365 => x"03003b04",
			3366 => x"000334a9",
			3367 => x"05005d04",
			3368 => x"015d34a9",
			3369 => x"ff6c34a9",
			3370 => x"06008d5c",
			3371 => x"07002720",
			3372 => x"0300381c",
			3373 => x"0c001a18",
			3374 => x"0c001810",
			3375 => x"06004408",
			3376 => x"01000504",
			3377 => x"feda3565",
			3378 => x"01053565",
			3379 => x"01000c04",
			3380 => x"fef33565",
			3381 => x"00da3565",
			3382 => x"04002004",
			3383 => x"ff0e3565",
			3384 => x"017a3565",
			3385 => x"fe9e3565",
			3386 => x"fe623565",
			3387 => x"05004820",
			3388 => x"09001e0c",
			3389 => x"07002b08",
			3390 => x"07002904",
			3391 => x"00ca3565",
			3392 => x"ff423565",
			3393 => x"01793565",
			3394 => x"0000b20c",
			3395 => x"04002608",
			3396 => x"07002d04",
			3397 => x"fe953565",
			3398 => x"00233565",
			3399 => x"01023565",
			3400 => x"07002a04",
			3401 => x"ff4a3565",
			3402 => x"fe533565",
			3403 => x"09002008",
			3404 => x"01000504",
			3405 => x"fed93565",
			3406 => x"01943565",
			3407 => x"09002108",
			3408 => x"01000804",
			3409 => x"00833565",
			3410 => x"fef83565",
			3411 => x"0200cc08",
			3412 => x"0a004804",
			3413 => x"013b3565",
			3414 => x"ff893565",
			3415 => x"febf3565",
			3416 => x"fe8b3565",
			3417 => x"05004858",
			3418 => x"0b001738",
			3419 => x"02008e18",
			3420 => x"05001208",
			3421 => x"07001704",
			3422 => x"005d3671",
			3423 => x"fed93671",
			3424 => x"08001604",
			3425 => x"ff2f3671",
			3426 => x"05003c08",
			3427 => x"0c001704",
			3428 => x"014c3671",
			3429 => x"ffdb3671",
			3430 => x"001d3671",
			3431 => x"0e006508",
			3432 => x"04002d04",
			3433 => x"fe8c3671",
			3434 => x"ffe93671",
			3435 => x"08001b08",
			3436 => x"03003104",
			3437 => x"feb33671",
			3438 => x"00503671",
			3439 => x"08001f08",
			3440 => x"06008e04",
			3441 => x"01523671",
			3442 => x"ff5b3671",
			3443 => x"08002004",
			3444 => x"fed23671",
			3445 => x"00963671",
			3446 => x"00009e18",
			3447 => x"0e004e14",
			3448 => x"09001e08",
			3449 => x"0b001804",
			3450 => x"ff993671",
			3451 => x"00d03671",
			3452 => x"01001004",
			3453 => x"fe8b3671",
			3454 => x"0d001c04",
			3455 => x"00623671",
			3456 => x"ffc13671",
			3457 => x"01083671",
			3458 => x"0a004004",
			3459 => x"fe9c3671",
			3460 => x"005a3671",
			3461 => x"07002704",
			3462 => x"ff473671",
			3463 => x"05004904",
			3464 => x"01763671",
			3465 => x"08001b0c",
			3466 => x"0e005f04",
			3467 => x"feb23671",
			3468 => x"0000d004",
			3469 => x"00e33671",
			3470 => x"fecb3671",
			3471 => x"01000a0c",
			3472 => x"0d001404",
			3473 => x"00333671",
			3474 => x"0a004804",
			3475 => x"01893671",
			3476 => x"ffa73671",
			3477 => x"0000c008",
			3478 => x"0a004204",
			3479 => x"00063671",
			3480 => x"01403671",
			3481 => x"0f009604",
			3482 => x"fee53671",
			3483 => x"00af3671",
			3484 => x"0d001320",
			3485 => x"0300351c",
			3486 => x"0a003718",
			3487 => x"0c001108",
			3488 => x"00007504",
			3489 => x"00fa3785",
			3490 => x"fffb3785",
			3491 => x"08001904",
			3492 => x"fec33785",
			3493 => x"0c001608",
			3494 => x"06007b04",
			3495 => x"00bf3785",
			3496 => x"ffcc3785",
			3497 => x"ff0f3785",
			3498 => x"01223785",
			3499 => x"fe9f3785",
			3500 => x"0c001930",
			3501 => x"0d00192c",
			3502 => x"0f00891c",
			3503 => x"0a002c0c",
			3504 => x"0c001808",
			3505 => x"03002204",
			3506 => x"006d3785",
			3507 => x"01643785",
			3508 => x"ffbd3785",
			3509 => x"0c001808",
			3510 => x"06005304",
			3511 => x"fffb3785",
			3512 => x"ff603785",
			3513 => x"09001f04",
			3514 => x"00083785",
			3515 => x"00f03785",
			3516 => x"01000808",
			3517 => x"03002d04",
			3518 => x"ffd63785",
			3519 => x"00be3785",
			3520 => x"03002404",
			3521 => x"00623785",
			3522 => x"fec83785",
			3523 => x"ff1d3785",
			3524 => x"0a004224",
			3525 => x"0000ae14",
			3526 => x"0e005610",
			3527 => x"08001d08",
			3528 => x"01000804",
			3529 => x"ffda3785",
			3530 => x"feca3785",
			3531 => x"07002704",
			3532 => x"ffaf3785",
			3533 => x"00d73785",
			3534 => x"00dc3785",
			3535 => x"0d001708",
			3536 => x"01000c04",
			3537 => x"fe9f3785",
			3538 => x"ffc23785",
			3539 => x"07002c04",
			3540 => x"00a23785",
			3541 => x"ff853785",
			3542 => x"0a004304",
			3543 => x"013c3785",
			3544 => x"0e006c0c",
			3545 => x"0000be04",
			3546 => x"00b03785",
			3547 => x"08001f04",
			3548 => x"fef73785",
			3549 => x"003b3785",
			3550 => x"0a004804",
			3551 => x"00fb3785",
			3552 => x"ffd53785",
			3553 => x"07003058",
			3554 => x"04004550",
			3555 => x"03003530",
			3556 => x"09001f20",
			3557 => x"04002510",
			3558 => x"08001b08",
			3559 => x"0c001104",
			3560 => x"00983839",
			3561 => x"fecd3839",
			3562 => x"0c001504",
			3563 => x"01033839",
			3564 => x"ffe03839",
			3565 => x"07002508",
			3566 => x"04002b04",
			3567 => x"00473839",
			3568 => x"ff3e3839",
			3569 => x"02010204",
			3570 => x"013e3839",
			3571 => x"ffc93839",
			3572 => x"0b001704",
			3573 => x"00713839",
			3574 => x"0000a108",
			3575 => x"02008e04",
			3576 => x"ff333839",
			3577 => x"00613839",
			3578 => x"fec33839",
			3579 => x"09001f08",
			3580 => x"07002904",
			3581 => x"fea53839",
			3582 => x"00333839",
			3583 => x"08001b08",
			3584 => x"09002004",
			3585 => x"00423839",
			3586 => x"ff013839",
			3587 => x"0200bb08",
			3588 => x"0e005504",
			3589 => x"ffe53839",
			3590 => x"01003839",
			3591 => x"07002c04",
			3592 => x"00673839",
			3593 => x"fef03839",
			3594 => x"03004704",
			3595 => x"00fd3839",
			3596 => x"ffe83839",
			3597 => x"ff133839",
			3598 => x"06008d68",
			3599 => x"0c001a3c",
			3600 => x"0a004338",
			3601 => x"0000811c",
			3602 => x"0100070c",
			3603 => x"08001804",
			3604 => x"fe8e390f",
			3605 => x"0b001604",
			3606 => x"00a3390f",
			3607 => x"fed4390f",
			3608 => x"0e003908",
			3609 => x"0b001504",
			3610 => x"016f390f",
			3611 => x"fe7b390f",
			3612 => x"05002b04",
			3613 => x"0142390f",
			3614 => x"01f5390f",
			3615 => x"0e004e0c",
			3616 => x"01000b08",
			3617 => x"01000604",
			3618 => x"0031390f",
			3619 => x"fe1c390f",
			3620 => x"014e390f",
			3621 => x"05003708",
			3622 => x"05002d04",
			3623 => x"008a390f",
			3624 => x"fee0390f",
			3625 => x"07002704",
			3626 => x"ffbe390f",
			3627 => x"014a390f",
			3628 => x"fe67390f",
			3629 => x"03003a18",
			3630 => x"0e005610",
			3631 => x"0000a208",
			3632 => x"00009604",
			3633 => x"fe66390f",
			3634 => x"0029390f",
			3635 => x"0000ab04",
			3636 => x"fcd0390f",
			3637 => x"fe85390f",
			3638 => x"06006304",
			3639 => x"0100390f",
			3640 => x"fdd1390f",
			3641 => x"0000d010",
			3642 => x"0e00620c",
			3643 => x"0000b908",
			3644 => x"0a004504",
			3645 => x"0168390f",
			3646 => x"00a6390f",
			3647 => x"fe66390f",
			3648 => x"01d7390f",
			3649 => x"fe5b390f",
			3650 => x"fe6e390f",
			3651 => x"0800180c",
			3652 => x"00003904",
			3653 => x"00743969",
			3654 => x"04003604",
			3655 => x"fe833969",
			3656 => x"ffed3969",
			3657 => x"07003020",
			3658 => x"0000fa18",
			3659 => x"0e006d10",
			3660 => x"01000504",
			3661 => x"fea23969",
			3662 => x"0e006608",
			3663 => x"06007004",
			3664 => x"00363969",
			3665 => x"fef03969",
			3666 => x"00e53969",
			3667 => x"0e007404",
			3668 => x"feb03969",
			3669 => x"00993969",
			3670 => x"05003804",
			3671 => x"ff043969",
			3672 => x"01873969",
			3673 => x"fea83969",
			3674 => x"0800180c",
			3675 => x"00003904",
			3676 => x"006a39cd",
			3677 => x"04003604",
			3678 => x"fe8a39cd",
			3679 => x"ffe539cd",
			3680 => x"07003024",
			3681 => x"0000fa1c",
			3682 => x"0e006d14",
			3683 => x"01000504",
			3684 => x"fead39cd",
			3685 => x"0e006508",
			3686 => x"06007004",
			3687 => x"002939cd",
			3688 => x"fea939cd",
			3689 => x"08001b04",
			3690 => x"001239cd",
			3691 => x"014e39cd",
			3692 => x"0e007404",
			3693 => x"fec839cd",
			3694 => x"009439cd",
			3695 => x"05003804",
			3696 => x"ff0e39cd",
			3697 => x"017839cd",
			3698 => x"feb139cd",
			3699 => x"02010230",
			3700 => x"0000fa28",
			3701 => x"01000504",
			3702 => x"fea43a41",
			3703 => x"0e006d1c",
			3704 => x"0b001910",
			3705 => x"03003e08",
			3706 => x"0e004e04",
			3707 => x"ffe33a41",
			3708 => x"006f3a41",
			3709 => x"04003e04",
			3710 => x"fed13a41",
			3711 => x"00383a41",
			3712 => x"0c001a04",
			3713 => x"00903a41",
			3714 => x"07002904",
			3715 => x"fec33a41",
			3716 => x"ffd63a41",
			3717 => x"0b001404",
			3718 => x"00f43a41",
			3719 => x"fe8a3a41",
			3720 => x"0e007404",
			3721 => x"01253a41",
			3722 => x"ff9e3a41",
			3723 => x"01000608",
			3724 => x"0d001304",
			3725 => x"ff693a41",
			3726 => x"007a3a41",
			3727 => x"fea83a41",
			3728 => x"0b001934",
			3729 => x"08001808",
			3730 => x"00004304",
			3731 => x"00053ae5",
			3732 => x"ffb03ae5",
			3733 => x"02010224",
			3734 => x"0500120c",
			3735 => x"04000d08",
			3736 => x"06001d04",
			3737 => x"00043ae5",
			3738 => x"ffe43ae5",
			3739 => x"00063ae5",
			3740 => x"0a004510",
			3741 => x"01000508",
			3742 => x"07002904",
			3743 => x"000f3ae5",
			3744 => x"ffdc3ae5",
			3745 => x"0e004e04",
			3746 => x"00143ae5",
			3747 => x"005b3ae5",
			3748 => x"04003e04",
			3749 => x"ffe23ae5",
			3750 => x"00143ae5",
			3751 => x"01000604",
			3752 => x"00093ae5",
			3753 => x"ffd73ae5",
			3754 => x"0c001a08",
			3755 => x"03002e04",
			3756 => x"ffec3ae5",
			3757 => x"00303ae5",
			3758 => x"04004c10",
			3759 => x"09001f04",
			3760 => x"00153ae5",
			3761 => x"0200ef04",
			3762 => x"ff713ae5",
			3763 => x"0e007e04",
			3764 => x"00103ae5",
			3765 => x"fff93ae5",
			3766 => x"0200c904",
			3767 => x"00213ae5",
			3768 => x"fff43ae5",
			3769 => x"0000b540",
			3770 => x"0c001a28",
			3771 => x"0800180c",
			3772 => x"00003704",
			3773 => x"003e3bc9",
			3774 => x"06005c04",
			3775 => x"ff6f3bc9",
			3776 => x"fff73bc9",
			3777 => x"0e004e10",
			3778 => x"0f00540c",
			3779 => x"04000a04",
			3780 => x"ff9a3bc9",
			3781 => x"01000704",
			3782 => x"ffdc3bc9",
			3783 => x"00b03bc9",
			3784 => x"ff823bc9",
			3785 => x"0200a808",
			3786 => x"07002904",
			3787 => x"00ef3bc9",
			3788 => x"00493bc9",
			3789 => x"ffff3bc9",
			3790 => x"03003a10",
			3791 => x"09001f08",
			3792 => x"09001e04",
			3793 => x"ffc93bc9",
			3794 => x"004c3bc9",
			3795 => x"0b001804",
			3796 => x"001f3bc9",
			3797 => x"ff1e3bc9",
			3798 => x"0a004504",
			3799 => x"00bd3bc9",
			3800 => x"fff23bc9",
			3801 => x"05004818",
			3802 => x"0f009008",
			3803 => x"01001104",
			3804 => x"fefb3bc9",
			3805 => x"00433bc9",
			3806 => x"05003f0c",
			3807 => x"06008d08",
			3808 => x"04001e04",
			3809 => x"ffdf3bc9",
			3810 => x"00b13bc9",
			3811 => x"ff8f3bc9",
			3812 => x"ff5a3bc9",
			3813 => x"06006b0c",
			3814 => x"0d001704",
			3815 => x"ff433bc9",
			3816 => x"0d001b04",
			3817 => x"ffff3bc9",
			3818 => x"fffa3bc9",
			3819 => x"07002f0c",
			3820 => x"04003c04",
			3821 => x"00053bc9",
			3822 => x"0d001404",
			3823 => x"ffe83bc9",
			3824 => x"00c03bc9",
			3825 => x"ffbe3bc9",
			3826 => x"0000ae34",
			3827 => x"0e005224",
			3828 => x"0000831c",
			3829 => x"03001008",
			3830 => x"04000e04",
			3831 => x"ffc53cb5",
			3832 => x"00003cb5",
			3833 => x"09001e0c",
			3834 => x"08001804",
			3835 => x"fff73cb5",
			3836 => x"01000704",
			3837 => x"fffd3cb5",
			3838 => x"007b3cb5",
			3839 => x"01001404",
			3840 => x"ffd73cb5",
			3841 => x"00043cb5",
			3842 => x"01000b04",
			3843 => x"ff8e3cb5",
			3844 => x"00253cb5",
			3845 => x"05003508",
			3846 => x"0c001504",
			3847 => x"00293cb5",
			3848 => x"ffb13cb5",
			3849 => x"05004e04",
			3850 => x"00963cb5",
			3851 => x"fff13cb5",
			3852 => x"05004820",
			3853 => x"04001a0c",
			3854 => x"09001a04",
			3855 => x"ffea3cb5",
			3856 => x"0c001704",
			3857 => x"003c3cb5",
			3858 => x"fff33cb5",
			3859 => x"0100120c",
			3860 => x"01000808",
			3861 => x"01000704",
			3862 => x"ffcf3cb5",
			3863 => x"000c3cb5",
			3864 => x"ff583cb5",
			3865 => x"01001304",
			3866 => x"00183cb5",
			3867 => x"fff73cb5",
			3868 => x"06006b0c",
			3869 => x"03003a04",
			3870 => x"00173cb5",
			3871 => x"08001f04",
			3872 => x"ffab3cb5",
			3873 => x"00003cb5",
			3874 => x"0a004308",
			3875 => x"08001d04",
			3876 => x"00653cb5",
			3877 => x"fff23cb5",
			3878 => x"05005908",
			3879 => x"0f009804",
			3880 => x"ffb13cb5",
			3881 => x"00143cb5",
			3882 => x"03004904",
			3883 => x"00473cb5",
			3884 => x"ffe13cb5",
			3885 => x"07002f30",
			3886 => x"0e00722c",
			3887 => x"00002504",
			3888 => x"fe5d3d29",
			3889 => x"01000710",
			3890 => x"0600760c",
			3891 => x"01000504",
			3892 => x"fe493d29",
			3893 => x"0000a904",
			3894 => x"00763d29",
			3895 => x"fe423d29",
			3896 => x"01a93d29",
			3897 => x"0b001a10",
			3898 => x"0a004508",
			3899 => x"05001204",
			3900 => x"ff9a3d29",
			3901 => x"017f3d29",
			3902 => x"04004304",
			3903 => x"ff843d29",
			3904 => x"fe4a3d29",
			3905 => x"06005b04",
			3906 => x"fe603d29",
			3907 => x"01773d29",
			3908 => x"fe5b3d29",
			3909 => x"0c001408",
			3910 => x"04001804",
			3911 => x"fe893d29",
			3912 => x"01403d29",
			3913 => x"fe5b3d29",
			3914 => x"05004338",
			3915 => x"0b001730",
			3916 => x"08001b10",
			3917 => x"0c001104",
			3918 => x"004c3ded",
			3919 => x"0f009e04",
			3920 => x"ff573ded",
			3921 => x"03003104",
			3922 => x"ffe83ded",
			3923 => x"00323ded",
			3924 => x"0d001618",
			3925 => x"0d00130c",
			3926 => x"02005c04",
			3927 => x"002f3ded",
			3928 => x"0e006804",
			3929 => x"ffc23ded",
			3930 => x"00123ded",
			3931 => x"01000904",
			3932 => x"fff53ded",
			3933 => x"06008104",
			3934 => x"00b63ded",
			3935 => x"fffc3ded",
			3936 => x"0000eb04",
			3937 => x"ffc33ded",
			3938 => x"00293ded",
			3939 => x"08001904",
			3940 => x"00073ded",
			3941 => x"ff5f3ded",
			3942 => x"0a004520",
			3943 => x"0b001810",
			3944 => x"0300390c",
			3945 => x"09001e04",
			3946 => x"ffad3ded",
			3947 => x"04003704",
			3948 => x"00963ded",
			3949 => x"00143ded",
			3950 => x"ff8e3ded",
			3951 => x"01000704",
			3952 => x"ffe53ded",
			3953 => x"07003008",
			3954 => x"03003a04",
			3955 => x"00293ded",
			3956 => x"00af3ded",
			3957 => x"fff33ded",
			3958 => x"07002e04",
			3959 => x"ff903ded",
			3960 => x"09002504",
			3961 => x"003a3ded",
			3962 => x"ffdb3ded",
			3963 => x"0e00773c",
			3964 => x"0500120c",
			3965 => x"04000504",
			3966 => x"00693e69",
			3967 => x"01000e04",
			3968 => x"fe403e69",
			3969 => x"fffd3e69",
			3970 => x"08001814",
			3971 => x"06006510",
			3972 => x"06005c0c",
			3973 => x"05001b04",
			3974 => x"00383e69",
			3975 => x"00009904",
			3976 => x"fe9e3e69",
			3977 => x"ff523e69",
			3978 => x"00e23e69",
			3979 => x"fe7a3e69",
			3980 => x"0c001508",
			3981 => x"00008904",
			3982 => x"018f3e69",
			3983 => x"008c3e69",
			3984 => x"05002504",
			3985 => x"fe8a3e69",
			3986 => x"0f008808",
			3987 => x"0000d604",
			3988 => x"00143e69",
			3989 => x"fe6f3e69",
			3990 => x"01000904",
			3991 => x"01ad3e69",
			3992 => x"ffa33e69",
			3993 => x"fe833e69",
			3994 => x"0200bb3c",
			3995 => x"0e005e30",
			3996 => x"0000ae20",
			3997 => x"08001604",
			3998 => x"ffa23f2d",
			3999 => x"0e005110",
			4000 => x"0c001608",
			4001 => x"0f004b04",
			4002 => x"007b3f2d",
			4003 => x"ffe73f2d",
			4004 => x"01000b04",
			4005 => x"ffa73f2d",
			4006 => x"00243f2d",
			4007 => x"04002304",
			4008 => x"ffda3f2d",
			4009 => x"05004e04",
			4010 => x"009e3f2d",
			4011 => x"00143f2d",
			4012 => x"0a003e08",
			4013 => x"0d001704",
			4014 => x"ff6e3f2d",
			4015 => x"00153f2d",
			4016 => x"03004004",
			4017 => x"00403f2d",
			4018 => x"ffe93f2d",
			4019 => x"04003608",
			4020 => x"01000904",
			4021 => x"ffc13f2d",
			4022 => x"00293f2d",
			4023 => x"00a83f2d",
			4024 => x"0700290c",
			4025 => x"0a002804",
			4026 => x"ffb53f2d",
			4027 => x"0b001504",
			4028 => x"00883f2d",
			4029 => x"fff73f2d",
			4030 => x"0a002704",
			4031 => x"002f3f2d",
			4032 => x"0000fa08",
			4033 => x"01000404",
			4034 => x"fffe3f2d",
			4035 => x"ff3b3f2d",
			4036 => x"00010404",
			4037 => x"003e3f2d",
			4038 => x"01000608",
			4039 => x"01000504",
			4040 => x"fff93f2d",
			4041 => x"00013f2d",
			4042 => x"ffae3f2d",
			4043 => x"07002c50",
			4044 => x"04001714",
			4045 => x"0c00130c",
			4046 => x"00009408",
			4047 => x"08001904",
			4048 => x"027a3ff9",
			4049 => x"03e53ff9",
			4050 => x"fe643ff9",
			4051 => x"0c001404",
			4052 => x"ff893ff9",
			4053 => x"fe503ff9",
			4054 => x"08001910",
			4055 => x"09001e08",
			4056 => x"05003e04",
			4057 => x"fe4a3ff9",
			4058 => x"ff2c3ff9",
			4059 => x"05004b04",
			4060 => x"04a93ff9",
			4061 => x"fe463ff9",
			4062 => x"0000b518",
			4063 => x"0c001b10",
			4064 => x"01000b08",
			4065 => x"0e004e04",
			4066 => x"014e3ff9",
			4067 => x"03b73ff9",
			4068 => x"0b001604",
			4069 => x"049f3ff9",
			4070 => x"03963ff9",
			4071 => x"03003404",
			4072 => x"fe403ff9",
			4073 => x"02763ff9",
			4074 => x"0d00150c",
			4075 => x"06007804",
			4076 => x"fe413ff9",
			4077 => x"06009804",
			4078 => x"03263ff9",
			4079 => x"fe5b3ff9",
			4080 => x"06006404",
			4081 => x"fe653ff9",
			4082 => x"04163ff9",
			4083 => x"07002f14",
			4084 => x"05004e0c",
			4085 => x"04002204",
			4086 => x"fe513ff9",
			4087 => x"0b001604",
			4088 => x"ffc33ff9",
			4089 => x"fe513ff9",
			4090 => x"0000ca04",
			4091 => x"048e3ff9",
			4092 => x"fff33ff9",
			4093 => x"fe503ff9",
			4094 => x"0000ba4c",
			4095 => x"0e004e30",
			4096 => x"00008320",
			4097 => x"09001e14",
			4098 => x"0500120c",
			4099 => x"04000604",
			4100 => x"001840e5",
			4101 => x"04000b04",
			4102 => x"ffce40e5",
			4103 => x"ffff40e5",
			4104 => x"08001804",
			4105 => x"fffe40e5",
			4106 => x"007440e5",
			4107 => x"01001408",
			4108 => x"0d001304",
			4109 => x"000240e5",
			4110 => x"ffcd40e5",
			4111 => x"000540e5",
			4112 => x"01000b08",
			4113 => x"08001904",
			4114 => x"000140e5",
			4115 => x"ff7c40e5",
			4116 => x"08002004",
			4117 => x"fffe40e5",
			4118 => x"001440e5",
			4119 => x"08002318",
			4120 => x"08001b10",
			4121 => x"05004c0c",
			4122 => x"05004408",
			4123 => x"05001f04",
			4124 => x"001140e5",
			4125 => x"ffc840e5",
			4126 => x"006b40e5",
			4127 => x"ffa740e5",
			4128 => x"0c001a04",
			4129 => x"009440e5",
			4130 => x"002540e5",
			4131 => x"ffca40e5",
			4132 => x"0d00150c",
			4133 => x"0f008604",
			4134 => x"ff7d40e5",
			4135 => x"06008204",
			4136 => x"002840e5",
			4137 => x"ffb740e5",
			4138 => x"0a004314",
			4139 => x"09001c04",
			4140 => x"ffca40e5",
			4141 => x"07002e08",
			4142 => x"0d001804",
			4143 => x"007d40e5",
			4144 => x"ffee40e5",
			4145 => x"05004a04",
			4146 => x"ffd040e5",
			4147 => x"001240e5",
			4148 => x"05005904",
			4149 => x"ffac40e5",
			4150 => x"05005e04",
			4151 => x"004240e5",
			4152 => x"ffd340e5",
			4153 => x"08001d48",
			4154 => x"0e005524",
			4155 => x"03003520",
			4156 => x"0e004d18",
			4157 => x"0100090c",
			4158 => x"02002b08",
			4159 => x"0d001304",
			4160 => x"002641c1",
			4161 => x"fff841c1",
			4162 => x"ff2341c1",
			4163 => x"0b001508",
			4164 => x"01000c04",
			4165 => x"00b241c1",
			4166 => x"000441c1",
			4167 => x"ff6a41c1",
			4168 => x"0000a604",
			4169 => x"00ca41c1",
			4170 => x"ff9a41c1",
			4171 => x"ff2e41c1",
			4172 => x"0500380c",
			4173 => x"01000b04",
			4174 => x"fef241c1",
			4175 => x"07002a04",
			4176 => x"009f41c1",
			4177 => x"ff8341c1",
			4178 => x"0a004514",
			4179 => x"04003e10",
			4180 => x"09002008",
			4181 => x"0e005b04",
			4182 => x"ffc141c1",
			4183 => x"00d341c1",
			4184 => x"0200bb04",
			4185 => x"000e41c1",
			4186 => x"ff1541c1",
			4187 => x"00f641c1",
			4188 => x"ff5d41c1",
			4189 => x"0200b014",
			4190 => x"0d001908",
			4191 => x"05001904",
			4192 => x"ffd641c1",
			4193 => x"010741c1",
			4194 => x"07002908",
			4195 => x"06004304",
			4196 => x"ffed41c1",
			4197 => x"006841c1",
			4198 => x"ff4b41c1",
			4199 => x"05002d10",
			4200 => x"0500290c",
			4201 => x"07002f04",
			4202 => x"ff7541c1",
			4203 => x"03002604",
			4204 => x"003641c1",
			4205 => x"fffa41c1",
			4206 => x"00c241c1",
			4207 => x"ff2f41c1",
			4208 => x"0000b22c",
			4209 => x"04004028",
			4210 => x"04003620",
			4211 => x"0b001718",
			4212 => x"0d00130c",
			4213 => x"0c001104",
			4214 => x"005a4295",
			4215 => x"08001b04",
			4216 => x"ff7f4295",
			4217 => x"00164295",
			4218 => x"06003808",
			4219 => x"0e002504",
			4220 => x"000c4295",
			4221 => x"fff94295",
			4222 => x"00834295",
			4223 => x"01001604",
			4224 => x"ff714295",
			4225 => x"00064295",
			4226 => x"0e005004",
			4227 => x"fff54295",
			4228 => x"00df4295",
			4229 => x"ff8b4295",
			4230 => x"0e006514",
			4231 => x"01001210",
			4232 => x"0b001808",
			4233 => x"04003e04",
			4234 => x"ff424295",
			4235 => x"fff84295",
			4236 => x"0000c004",
			4237 => x"00424295",
			4238 => x"ff964295",
			4239 => x"00224295",
			4240 => x"06007910",
			4241 => x"0f007b08",
			4242 => x"0f007704",
			4243 => x"00224295",
			4244 => x"ffbb4295",
			4245 => x"0c001b04",
			4246 => x"007b4295",
			4247 => x"ffe54295",
			4248 => x"07002c10",
			4249 => x"05002904",
			4250 => x"ff9d4295",
			4251 => x"0d001308",
			4252 => x"0d001204",
			4253 => x"00304295",
			4254 => x"ffbc4295",
			4255 => x"00694295",
			4256 => x"05002308",
			4257 => x"0b001404",
			4258 => x"00214295",
			4259 => x"fffb4295",
			4260 => x"ff794295",
			4261 => x"0d00131c",
			4262 => x"00008810",
			4263 => x"05001208",
			4264 => x"02002904",
			4265 => x"00124361",
			4266 => x"ffca4361",
			4267 => x"0d001104",
			4268 => x"00054361",
			4269 => x"004a4361",
			4270 => x"06008c04",
			4271 => x"ff7d4361",
			4272 => x"00010e04",
			4273 => x"002c4361",
			4274 => x"ffed4361",
			4275 => x"0d001940",
			4276 => x"08001b14",
			4277 => x"0d001710",
			4278 => x"0900200c",
			4279 => x"04002908",
			4280 => x"07002104",
			4281 => x"00064361",
			4282 => x"ffd34361",
			4283 => x"003b4361",
			4284 => x"ff924361",
			4285 => x"00314361",
			4286 => x"07002714",
			4287 => x"03002c10",
			4288 => x"0c001808",
			4289 => x"04001d04",
			4290 => x"00014361",
			4291 => x"00614361",
			4292 => x"06004004",
			4293 => x"ffea4361",
			4294 => x"00024361",
			4295 => x"ffab4361",
			4296 => x"0200ac08",
			4297 => x"06005304",
			4298 => x"fffb4361",
			4299 => x"00984361",
			4300 => x"0e006508",
			4301 => x"0b001804",
			4302 => x"ffb34361",
			4303 => x"fffd4361",
			4304 => x"08001f04",
			4305 => x"00554361",
			4306 => x"ffde4361",
			4307 => x"07002908",
			4308 => x"06004404",
			4309 => x"fffb4361",
			4310 => x"00184361",
			4311 => x"ffa84361",
			4312 => x"0000ae40",
			4313 => x"0e00522c",
			4314 => x"0b001208",
			4315 => x"00004904",
			4316 => x"006c4455",
			4317 => x"fff34455",
			4318 => x"01000b10",
			4319 => x"0400340c",
			4320 => x"08001d04",
			4321 => x"ff5e4455",
			4322 => x"08001f04",
			4323 => x"ffef4455",
			4324 => x"00114455",
			4325 => x"ffec4455",
			4326 => x"0400170c",
			4327 => x"05001804",
			4328 => x"ffd94455",
			4329 => x"05001b04",
			4330 => x"00064455",
			4331 => x"fffb4455",
			4332 => x"0c001b04",
			4333 => x"00804455",
			4334 => x"ffe84455",
			4335 => x"04002308",
			4336 => x"0c001504",
			4337 => x"003c4455",
			4338 => x"ffad4455",
			4339 => x"05005008",
			4340 => x"04003604",
			4341 => x"002f4455",
			4342 => x"00d84455",
			4343 => x"fff24455",
			4344 => x"0e00651c",
			4345 => x"04004414",
			4346 => x"01001210",
			4347 => x"08001604",
			4348 => x"00214455",
			4349 => x"07002d08",
			4350 => x"0c001b04",
			4351 => x"ff454455",
			4352 => x"ffe54455",
			4353 => x"00114455",
			4354 => x"002b4455",
			4355 => x"07002f04",
			4356 => x"003e4455",
			4357 => x"ffe34455",
			4358 => x"0000d60c",
			4359 => x"0f008904",
			4360 => x"00924455",
			4361 => x"07002e04",
			4362 => x"ffd54455",
			4363 => x"000f4455",
			4364 => x"07002c10",
			4365 => x"0300310c",
			4366 => x"07002b04",
			4367 => x"ff914455",
			4368 => x"01000804",
			4369 => x"fff94455",
			4370 => x"003b4455",
			4371 => x"00674455",
			4372 => x"ff5c4455",
			4373 => x"0d001540",
			4374 => x"0300352c",
			4375 => x"05004424",
			4376 => x"0b001410",
			4377 => x"08001604",
			4378 => x"ffbc4561",
			4379 => x"04000d04",
			4380 => x"ffdb4561",
			4381 => x"0e007104",
			4382 => x"00904561",
			4383 => x"ffe14561",
			4384 => x"0d001304",
			4385 => x"ff5c4561",
			4386 => x"07002808",
			4387 => x"01000b04",
			4388 => x"ff824561",
			4389 => x"00134561",
			4390 => x"0e007204",
			4391 => x"00744561",
			4392 => x"ffea4561",
			4393 => x"08001b04",
			4394 => x"00a84561",
			4395 => x"ffeb4561",
			4396 => x"0b001808",
			4397 => x"07002b04",
			4398 => x"ff2e4561",
			4399 => x"ffec4561",
			4400 => x"04003c04",
			4401 => x"ffb64561",
			4402 => x"0c001b04",
			4403 => x"00784561",
			4404 => x"ffdd4561",
			4405 => x"07002920",
			4406 => x"0c001a10",
			4407 => x"03002208",
			4408 => x"07001f04",
			4409 => x"00124561",
			4410 => x"ffdc4561",
			4411 => x"0e004d04",
			4412 => x"00224561",
			4413 => x"00e74561",
			4414 => x"0000a90c",
			4415 => x"09002104",
			4416 => x"ff7e4561",
			4417 => x"09002204",
			4418 => x"00064561",
			4419 => x"fff74561",
			4420 => x"00484561",
			4421 => x"04003e18",
			4422 => x"0f008e10",
			4423 => x"0000b208",
			4424 => x"00009704",
			4425 => x"ffc34561",
			4426 => x"00204561",
			4427 => x"06007004",
			4428 => x"ffff4561",
			4429 => x"ff454561",
			4430 => x"07002e04",
			4431 => x"00654561",
			4432 => x"ffca4561",
			4433 => x"0a004804",
			4434 => x"00814561",
			4435 => x"04004d04",
			4436 => x"ffbe4561",
			4437 => x"04005a04",
			4438 => x"00094561",
			4439 => x"fff94561",
			4440 => x"0a004358",
			4441 => x"0400343c",
			4442 => x"0b00172c",
			4443 => x"0d001314",
			4444 => x"02005c08",
			4445 => x"0c001404",
			4446 => x"005e462d",
			4447 => x"ffed462d",
			4448 => x"06008c04",
			4449 => x"ff8c462d",
			4450 => x"0f00a904",
			4451 => x"0029462d",
			4452 => x"ffed462d",
			4453 => x"0d001610",
			4454 => x"06008008",
			4455 => x"01000904",
			4456 => x"ffec462d",
			4457 => x"00ac462d",
			4458 => x"03002f04",
			4459 => x"ffb8462d",
			4460 => x"001a462d",
			4461 => x"0000eb04",
			4462 => x"ffba462d",
			4463 => x"002b462d",
			4464 => x"04003108",
			4465 => x"08001904",
			4466 => x"0008462d",
			4467 => x"ff61462d",
			4468 => x"04003204",
			4469 => x"0023462d",
			4470 => x"ffeb462d",
			4471 => x"0c001804",
			4472 => x"ffd6462d",
			4473 => x"0000ae08",
			4474 => x"0a003e04",
			4475 => x"009b462d",
			4476 => x"0016462d",
			4477 => x"0e006108",
			4478 => x"0c001904",
			4479 => x"0013462d",
			4480 => x"ff88462d",
			4481 => x"09002204",
			4482 => x"007a462d",
			4483 => x"fff8462d",
			4484 => x"0e006c08",
			4485 => x"0000b904",
			4486 => x"0009462d",
			4487 => x"ff5e462d",
			4488 => x"01000904",
			4489 => x"0036462d",
			4490 => x"fff7462d",
			4491 => x"0000b54c",
			4492 => x"0e005234",
			4493 => x"00008324",
			4494 => x"09001e18",
			4495 => x"0500120c",
			4496 => x"04000604",
			4497 => x"00184729",
			4498 => x"0d001304",
			4499 => x"ffc14729",
			4500 => x"00054729",
			4501 => x"0c001908",
			4502 => x"01000704",
			4503 => x"fffc4729",
			4504 => x"00804729",
			4505 => x"fff54729",
			4506 => x"01001608",
			4507 => x"0d001304",
			4508 => x"00024729",
			4509 => x"ffc74729",
			4510 => x"00044729",
			4511 => x"01000d08",
			4512 => x"0e004d04",
			4513 => x"ff744729",
			4514 => x"ffe64729",
			4515 => x"0e004704",
			4516 => x"fff94729",
			4517 => x"00294729",
			4518 => x"08002314",
			4519 => x"08001b0c",
			4520 => x"03003508",
			4521 => x"0f007a04",
			4522 => x"00394729",
			4523 => x"ffec4729",
			4524 => x"ffcd4729",
			4525 => x"0c001a04",
			4526 => x"00a34729",
			4527 => x"00134729",
			4528 => x"ffb94729",
			4529 => x"06007514",
			4530 => x"01001210",
			4531 => x"0e00680c",
			4532 => x"0d001704",
			4533 => x"ff4a4729",
			4534 => x"05005804",
			4535 => x"00204729",
			4536 => x"ffe54729",
			4537 => x"002b4729",
			4538 => x"00274729",
			4539 => x"04003118",
			4540 => x"07002908",
			4541 => x"0a002804",
			4542 => x"ffda4729",
			4543 => x"00404729",
			4544 => x"0a002704",
			4545 => x"00274729",
			4546 => x"01000808",
			4547 => x"01000504",
			4548 => x"ffda4729",
			4549 => x"00154729",
			4550 => x"ff694729",
			4551 => x"0c001b04",
			4552 => x"00694729",
			4553 => x"ffdd4729",
			4554 => x"02009730",
			4555 => x"0e004820",
			4556 => x"07001704",
			4557 => x"004e481d",
			4558 => x"08001d10",
			4559 => x"01000a04",
			4560 => x"ff78481d",
			4561 => x"01000c08",
			4562 => x"01000b04",
			4563 => x"0000481d",
			4564 => x"0012481d",
			4565 => x"ffe0481d",
			4566 => x"05001e04",
			4567 => x"ffe3481d",
			4568 => x"0c001a04",
			4569 => x"0047481d",
			4570 => x"fffa481d",
			4571 => x"0100120c",
			4572 => x"08001904",
			4573 => x"000f481d",
			4574 => x"07002504",
			4575 => x"0000481d",
			4576 => x"00ac481d",
			4577 => x"fff0481d",
			4578 => x"0e005a18",
			4579 => x"0d00150c",
			4580 => x"03003508",
			4581 => x"01000704",
			4582 => x"0017481d",
			4583 => x"ffde481d",
			4584 => x"ff71481d",
			4585 => x"0c001a04",
			4586 => x"0048481d",
			4587 => x"0a003b04",
			4588 => x"0005481d",
			4589 => x"ff8b481d",
			4590 => x"0200b70c",
			4591 => x"03002f08",
			4592 => x"0e007204",
			4593 => x"ffde481d",
			4594 => x"0018481d",
			4595 => x"0082481d",
			4596 => x"0700290c",
			4597 => x"0a002804",
			4598 => x"ffb8481d",
			4599 => x"0a003404",
			4600 => x"0079481d",
			4601 => x"0003481d",
			4602 => x"01000610",
			4603 => x"0200d908",
			4604 => x"06007104",
			4605 => x"ffdd481d",
			4606 => x"0061481d",
			4607 => x"03003304",
			4608 => x"0017481d",
			4609 => x"ffac481d",
			4610 => x"0a002704",
			4611 => x"0023481d",
			4612 => x"04004c04",
			4613 => x"ff59481d",
			4614 => x"0016481d",
			4615 => x"0000c038",
			4616 => x"00002504",
			4617 => x"fe5848c1",
			4618 => x"01000714",
			4619 => x"01000504",
			4620 => x"fe4048c1",
			4621 => x"0000a90c",
			4622 => x"0e004d08",
			4623 => x"00004f04",
			4624 => x"011448c1",
			4625 => x"fe4548c1",
			4626 => x"025348c1",
			4627 => x"fe3848c1",
			4628 => x"0b001a18",
			4629 => x"0c00150c",
			4630 => x"08001904",
			4631 => x"017e48c1",
			4632 => x"0e004204",
			4633 => x"029b48c1",
			4634 => x"039048c1",
			4635 => x"05002504",
			4636 => x"fe5a48c1",
			4637 => x"0d001304",
			4638 => x"fff448c1",
			4639 => x"020448c1",
			4640 => x"04002804",
			4641 => x"fe5a48c1",
			4642 => x"011148c1",
			4643 => x"0e007218",
			4644 => x"0f007604",
			4645 => x"fe5248c1",
			4646 => x"07002f10",
			4647 => x"0e006504",
			4648 => x"feeb48c1",
			4649 => x"0b001604",
			4650 => x"ff4548c1",
			4651 => x"0e006804",
			4652 => x"013548c1",
			4653 => x"034e48c1",
			4654 => x"fe5c48c1",
			4655 => x"fe5748c1",
			4656 => x"0d001324",
			4657 => x"03003520",
			4658 => x"0300331c",
			4659 => x"0c001108",
			4660 => x"00004104",
			4661 => x"00c449a5",
			4662 => x"000749a5",
			4663 => x"0600440c",
			4664 => x"0e002d04",
			4665 => x"ff9249a5",
			4666 => x"02006b04",
			4667 => x"006849a5",
			4668 => x"ffd049a5",
			4669 => x"01000b04",
			4670 => x"ff0449a5",
			4671 => x"ffef49a5",
			4672 => x"00c449a5",
			4673 => x"fee149a5",
			4674 => x"0000ae2c",
			4675 => x"0e005120",
			4676 => x"01000b14",
			4677 => x"0b001708",
			4678 => x"0a002a04",
			4679 => x"006d49a5",
			4680 => x"ffb549a5",
			4681 => x"01000808",
			4682 => x"01000704",
			4683 => x"ffba49a5",
			4684 => x"001349a5",
			4685 => x"fef349a5",
			4686 => x"0c001b08",
			4687 => x"05001604",
			4688 => x"fff449a5",
			4689 => x"00f549a5",
			4690 => x"ffac49a5",
			4691 => x"05003504",
			4692 => x"ffc449a5",
			4693 => x"07002b04",
			4694 => x"012649a5",
			4695 => x"001249a5",
			4696 => x"06006508",
			4697 => x"0a004204",
			4698 => x"fec849a5",
			4699 => x"004749a5",
			4700 => x"09001c0c",
			4701 => x"04001808",
			4702 => x"0c001504",
			4703 => x"003b49a5",
			4704 => x"fff549a5",
			4705 => x"ff0a49a5",
			4706 => x"0700300c",
			4707 => x"09001d04",
			4708 => x"00fe49a5",
			4709 => x"04003904",
			4710 => x"ffea49a5",
			4711 => x"008e49a5",
			4712 => x"ff5349a5",
			4713 => x"00009e2c",
			4714 => x"08001604",
			4715 => x"ffa94a89",
			4716 => x"06005524",
			4717 => x"00008318",
			4718 => x"0c001910",
			4719 => x"05001208",
			4720 => x"0a000a04",
			4721 => x"000e4a89",
			4722 => x"ffce4a89",
			4723 => x"01000704",
			4724 => x"00044a89",
			4725 => x"009e4a89",
			4726 => x"01001604",
			4727 => x"ffc24a89",
			4728 => x"00004a89",
			4729 => x"01000b08",
			4730 => x"00009304",
			4731 => x"ff884a89",
			4732 => x"fffc4a89",
			4733 => x"00124a89",
			4734 => x"008d4a89",
			4735 => x"04003e34",
			4736 => x"0e006510",
			4737 => x"0d001708",
			4738 => x"05005004",
			4739 => x"ff564a89",
			4740 => x"fff94a89",
			4741 => x"05003704",
			4742 => x"ffa54a89",
			4743 => x"004a4a89",
			4744 => x"03002410",
			4745 => x"0500280c",
			4746 => x"0e007604",
			4747 => x"ffbb4a89",
			4748 => x"0000d804",
			4749 => x"001e4a89",
			4750 => x"fff84a89",
			4751 => x"00724a89",
			4752 => x"0d001208",
			4753 => x"06009a04",
			4754 => x"00414a89",
			4755 => x"fff64a89",
			4756 => x"04003b08",
			4757 => x"04003104",
			4758 => x"ff674a89",
			4759 => x"ffe44a89",
			4760 => x"000b4a89",
			4761 => x"0a004808",
			4762 => x"03003e04",
			4763 => x"fff34a89",
			4764 => x"00664a89",
			4765 => x"04004d04",
			4766 => x"ffa14a89",
			4767 => x"04005a04",
			4768 => x"00044a89",
			4769 => x"fffa4a89",
			4770 => x"04004748",
			4771 => x"04004040",
			4772 => x"03003e34",
			4773 => x"04003420",
			4774 => x"0b001710",
			4775 => x"08001b08",
			4776 => x"0c001104",
			4777 => x"00be4b3d",
			4778 => x"ff514b3d",
			4779 => x"0a003704",
			4780 => x"007d4b3d",
			4781 => x"fefc4b3d",
			4782 => x"04003108",
			4783 => x"08001904",
			4784 => x"00114b3d",
			4785 => x"fed14b3d",
			4786 => x"03003504",
			4787 => x"00934b3d",
			4788 => x"ff8e4b3d",
			4789 => x"04003504",
			4790 => x"015c4b3d",
			4791 => x"0000ae08",
			4792 => x"0f005d04",
			4793 => x"ffb54b3d",
			4794 => x"01614b3d",
			4795 => x"0e005b04",
			4796 => x"fe934b3d",
			4797 => x"004c4b3d",
			4798 => x"0c001b04",
			4799 => x"fedc4b3d",
			4800 => x"0e006004",
			4801 => x"00bb4b3d",
			4802 => x"ff6c4b3d",
			4803 => x"08001c04",
			4804 => x"fea34b3d",
			4805 => x"00424b3d",
			4806 => x"0d001504",
			4807 => x"ff264b3d",
			4808 => x"05006304",
			4809 => x"01714b3d",
			4810 => x"0f007208",
			4811 => x"06006a04",
			4812 => x"ffeb4b3d",
			4813 => x"00694b3d",
			4814 => x"ff4a4b3d",
			4815 => x"00008318",
			4816 => x"05001208",
			4817 => x"07001804",
			4818 => x"00244c09",
			4819 => x"ff694c09",
			4820 => x"0c001908",
			4821 => x"08001804",
			4822 => x"ffff4c09",
			4823 => x"00f54c09",
			4824 => x"01001604",
			4825 => x"ff8e4c09",
			4826 => x"001c4c09",
			4827 => x"0e004d08",
			4828 => x"08001f04",
			4829 => x"ff024c09",
			4830 => x"00164c09",
			4831 => x"05003828",
			4832 => x"01000b0c",
			4833 => x"05002208",
			4834 => x"05002104",
			4835 => x"ffc54c09",
			4836 => x"00204c09",
			4837 => x"fee74c09",
			4838 => x"0d00160c",
			4839 => x"05002204",
			4840 => x"ff8d4c09",
			4841 => x"0a002d04",
			4842 => x"01074c09",
			4843 => x"ffa84c09",
			4844 => x"0000eb08",
			4845 => x"0f006504",
			4846 => x"00424c09",
			4847 => x"ff024c09",
			4848 => x"02010204",
			4849 => x"00734c09",
			4850 => x"ffdb4c09",
			4851 => x"00009e04",
			4852 => x"00e34c09",
			4853 => x"06007510",
			4854 => x"0000c008",
			4855 => x"0e005c04",
			4856 => x"ffb94c09",
			4857 => x"00fe4c09",
			4858 => x"08001f04",
			4859 => x"ff074c09",
			4860 => x"00214c09",
			4861 => x"08001f08",
			4862 => x"0c001b04",
			4863 => x"00a64c09",
			4864 => x"ffc34c09",
			4865 => x"ff864c09",
			4866 => x"0e007240",
			4867 => x"0c001e3c",
			4868 => x"08001810",
			4869 => x"09001e08",
			4870 => x"04000a04",
			4871 => x"ffae4c8d",
			4872 => x"fe5b4c8d",
			4873 => x"0b001704",
			4874 => x"01944c8d",
			4875 => x"fe5e4c8d",
			4876 => x"0c001610",
			4877 => x"00008908",
			4878 => x"05001304",
			4879 => x"003d4c8d",
			4880 => x"01e44c8d",
			4881 => x"0d001304",
			4882 => x"fe694c8d",
			4883 => x"006f4c8d",
			4884 => x"05003710",
			4885 => x"0b001608",
			4886 => x"01000b04",
			4887 => x"fe3a4c8d",
			4888 => x"00fb4c8d",
			4889 => x"05003104",
			4890 => x"fe3c4c8d",
			4891 => x"ff624c8d",
			4892 => x"0e004d04",
			4893 => x"ff694c8d",
			4894 => x"00009e04",
			4895 => x"02074c8d",
			4896 => x"00a14c8d",
			4897 => x"fe684c8d",
			4898 => x"fe634c8d",
			4899 => x"0000b240",
			4900 => x"0e005230",
			4901 => x"0000831c",
			4902 => x"05001208",
			4903 => x"07001704",
			4904 => x"00464d91",
			4905 => x"ff3c4d91",
			4906 => x"0c001a10",
			4907 => x"0e003808",
			4908 => x"0c001504",
			4909 => x"00db4d91",
			4910 => x"ff764d91",
			4911 => x"09001c04",
			4912 => x"00154d91",
			4913 => x"012a4d91",
			4914 => x"ff794d91",
			4915 => x"0d00150c",
			4916 => x"05004708",
			4917 => x"05004104",
			4918 => x"ff2c4d91",
			4919 => x"00564d91",
			4920 => x"feea4d91",
			4921 => x"0f005204",
			4922 => x"ffa94d91",
			4923 => x"00ad4d91",
			4924 => x"0400360c",
			4925 => x"0a003208",
			4926 => x"0d001304",
			4927 => x"fffd4d91",
			4928 => x"00cd4d91",
			4929 => x"ff814d91",
			4930 => x"01384d91",
			4931 => x"0600660c",
			4932 => x"09002304",
			4933 => x"fee24d91",
			4934 => x"08002304",
			4935 => x"00314d91",
			4936 => x"fffb4d91",
			4937 => x"06007018",
			4938 => x"0d001408",
			4939 => x"05005404",
			4940 => x"ff314d91",
			4941 => x"001c4d91",
			4942 => x"0a004504",
			4943 => x"01324d91",
			4944 => x"06006b04",
			4945 => x"ff874d91",
			4946 => x"0e006604",
			4947 => x"00524d91",
			4948 => x"fffa4d91",
			4949 => x"0e006504",
			4950 => x"fec94d91",
			4951 => x"07002c0c",
			4952 => x"05002804",
			4953 => x"ff144d91",
			4954 => x"02010204",
			4955 => x"00d94d91",
			4956 => x"ffb34d91",
			4957 => x"04003c08",
			4958 => x"0c001404",
			4959 => x"00304d91",
			4960 => x"fece4d91",
			4961 => x"0f008104",
			4962 => x"00954d91",
			4963 => x"ffa04d91",
			4964 => x"00009e2c",
			4965 => x"08001604",
			4966 => x"ff6e4e5d",
			4967 => x"04003624",
			4968 => x"0c00160c",
			4969 => x"04000d04",
			4970 => x"ffce4e5d",
			4971 => x"02008004",
			4972 => x"00d44e5d",
			4973 => x"000b4e5d",
			4974 => x"0d00150c",
			4975 => x"01000b08",
			4976 => x"09002004",
			4977 => x"ff304e5d",
			4978 => x"fffc4e5d",
			4979 => x"00214e5d",
			4980 => x"05002f08",
			4981 => x"09001e04",
			4982 => x"00044e5d",
			4983 => x"ff9b4e5d",
			4984 => x"00744e5d",
			4985 => x"00c24e5d",
			4986 => x"04002514",
			4987 => x"0e006504",
			4988 => x"ff094e5d",
			4989 => x"0f008b04",
			4990 => x"00a14e5d",
			4991 => x"0c001704",
			4992 => x"ff2c4e5d",
			4993 => x"03002404",
			4994 => x"00614e5d",
			4995 => x"ffcc4e5d",
			4996 => x"0e005204",
			4997 => x"ff4b4e5d",
			4998 => x"0000ae08",
			4999 => x"0a003e04",
			5000 => x"00d24e5d",
			5001 => x"ffcc4e5d",
			5002 => x"04003e0c",
			5003 => x"0e005b04",
			5004 => x"ff0d4e5d",
			5005 => x"03003b04",
			5006 => x"004b4e5d",
			5007 => x"ff534e5d",
			5008 => x"0d001508",
			5009 => x"08001904",
			5010 => x"ffa84e5d",
			5011 => x"00094e5d",
			5012 => x"07002f04",
			5013 => x"00d74e5d",
			5014 => x"ffb34e5d",
			5015 => x"0d001324",
			5016 => x"03003520",
			5017 => x"0300331c",
			5018 => x"00008814",
			5019 => x"05001208",
			5020 => x"04000b04",
			5021 => x"ff3c4f21",
			5022 => x"fff54f21",
			5023 => x"0c001608",
			5024 => x"08001804",
			5025 => x"ffd84f21",
			5026 => x"01004f21",
			5027 => x"ff724f21",
			5028 => x"0a003604",
			5029 => x"fed44f21",
			5030 => x"ffcc4f21",
			5031 => x"00e24f21",
			5032 => x"fecb4f21",
			5033 => x"0700303c",
			5034 => x"09002124",
			5035 => x"05004b1c",
			5036 => x"0f00690c",
			5037 => x"0e004e08",
			5038 => x"0b001704",
			5039 => x"00a94f21",
			5040 => x"fef04f21",
			5041 => x"01094f21",
			5042 => x"0e007008",
			5043 => x"03003404",
			5044 => x"ff7d4f21",
			5045 => x"004f4f21",
			5046 => x"06009104",
			5047 => x"00da4f21",
			5048 => x"ffa94f21",
			5049 => x"03004004",
			5050 => x"ff514f21",
			5051 => x"00564f21",
			5052 => x"0a003e10",
			5053 => x"07002b0c",
			5054 => x"0000a208",
			5055 => x"0a002d04",
			5056 => x"ffcf4f21",
			5057 => x"00a64f21",
			5058 => x"ffc44f21",
			5059 => x"ff374f21",
			5060 => x"0a004804",
			5061 => x"010d4f21",
			5062 => x"ffac4f21",
			5063 => x"ff2c4f21",
			5064 => x"0e00723c",
			5065 => x"04004734",
			5066 => x"04004330",
			5067 => x"0000ae1c",
			5068 => x"0e005110",
			5069 => x"00009e08",
			5070 => x"0c001a04",
			5071 => x"00904f9d",
			5072 => x"fe9f4f9d",
			5073 => x"0d001704",
			5074 => x"fe064f9d",
			5075 => x"00d94f9d",
			5076 => x"04003608",
			5077 => x"0f006404",
			5078 => x"01074f9d",
			5079 => x"ffcc4f9d",
			5080 => x"01ab4f9d",
			5081 => x"0e005b04",
			5082 => x"fe214f9d",
			5083 => x"03003e08",
			5084 => x"05002804",
			5085 => x"fed84f9d",
			5086 => x"00824f9d",
			5087 => x"0000cc04",
			5088 => x"ff5a4f9d",
			5089 => x"fe654f9d",
			5090 => x"fe5d4f9d",
			5091 => x"03004904",
			5092 => x"01c84f9d",
			5093 => x"fead4f9d",
			5094 => x"fe714f9d",
			5095 => x"08001b24",
			5096 => x"0c001104",
			5097 => x"004a5071",
			5098 => x"0f009e18",
			5099 => x"05004404",
			5100 => x"ff4a5071",
			5101 => x"05004c08",
			5102 => x"0000b404",
			5103 => x"00925071",
			5104 => x"ffe75071",
			5105 => x"03004104",
			5106 => x"ff595071",
			5107 => x"03004704",
			5108 => x"000b5071",
			5109 => x"ffec5071",
			5110 => x"04002804",
			5111 => x"ffe25071",
			5112 => x"00395071",
			5113 => x"06008640",
			5114 => x"0d001934",
			5115 => x"07002718",
			5116 => x"0b001508",
			5117 => x"05003204",
			5118 => x"00875071",
			5119 => x"fff75071",
			5120 => x"0d001508",
			5121 => x"0b001804",
			5122 => x"ff685071",
			5123 => x"fffb5071",
			5124 => x"09001e04",
			5125 => x"ffe65071",
			5126 => x"00395071",
			5127 => x"0b00190c",
			5128 => x"0d001304",
			5129 => x"fffa5071",
			5130 => x"05002204",
			5131 => x"fff75071",
			5132 => x"00a85071",
			5133 => x"0200bd08",
			5134 => x"02009c04",
			5135 => x"ffbd5071",
			5136 => x"00785071",
			5137 => x"0e006c04",
			5138 => x"ffa75071",
			5139 => x"00125071",
			5140 => x"07002908",
			5141 => x"06004404",
			5142 => x"fff85071",
			5143 => x"00215071",
			5144 => x"ff8d5071",
			5145 => x"01000604",
			5146 => x"00145071",
			5147 => x"ff815071",
			5148 => x"06008664",
			5149 => x"08001b20",
			5150 => x"0000c71c",
			5151 => x"0500440c",
			5152 => x"0c001104",
			5153 => x"00ed514d",
			5154 => x"01000a04",
			5155 => x"fea4514d",
			5156 => x"ff94514d",
			5157 => x"05004c08",
			5158 => x"0000ab04",
			5159 => x"013b514d",
			5160 => x"005b514d",
			5161 => x"0f006a04",
			5162 => x"feb5514d",
			5163 => x"0028514d",
			5164 => x"fecd514d",
			5165 => x"0e004e24",
			5166 => x"0c001608",
			5167 => x"0f005204",
			5168 => x"0109514d",
			5169 => x"0022514d",
			5170 => x"08001f10",
			5171 => x"07002708",
			5172 => x"0d001504",
			5173 => x"fe90514d",
			5174 => x"ffc5514d",
			5175 => x"08001d04",
			5176 => x"ff68514d",
			5177 => x"006c514d",
			5178 => x"06004004",
			5179 => x"ff98514d",
			5180 => x"0b001b04",
			5181 => x"00d7514d",
			5182 => x"fff3514d",
			5183 => x"0d001814",
			5184 => x"00009f04",
			5185 => x"0168514d",
			5186 => x"0e005a08",
			5187 => x"0e005604",
			5188 => x"ff44514d",
			5189 => x"fff9514d",
			5190 => x"0200ae04",
			5191 => x"0169514d",
			5192 => x"0052514d",
			5193 => x"0e005b08",
			5194 => x"08002404",
			5195 => x"00e1514d",
			5196 => x"ff56514d",
			5197 => x"fecd514d",
			5198 => x"01000808",
			5199 => x"0b001604",
			5200 => x"ff19514d",
			5201 => x"00a7514d",
			5202 => x"feb3514d",
			5203 => x"06008d50",
			5204 => x"0d001944",
			5205 => x"01000b24",
			5206 => x"0000fa20",
			5207 => x"05004410",
			5208 => x"07002108",
			5209 => x"0c001704",
			5210 => x"009c51f1",
			5211 => x"fe7b51f1",
			5212 => x"09001c04",
			5213 => x"ffa351f1",
			5214 => x"fe6151f1",
			5215 => x"03003508",
			5216 => x"08001b04",
			5217 => x"026251f1",
			5218 => x"ffe351f1",
			5219 => x"0d001404",
			5220 => x"fef551f1",
			5221 => x"009151f1",
			5222 => x"018e51f1",
			5223 => x"0200a114",
			5224 => x"0c001a0c",
			5225 => x"04000d04",
			5226 => x"ffb851f1",
			5227 => x"0d001204",
			5228 => x"00de51f1",
			5229 => x"01b351f1",
			5230 => x"06002d04",
			5231 => x"fee051f1",
			5232 => x"001851f1",
			5233 => x"0e005b04",
			5234 => x"fe4c51f1",
			5235 => x"0200c904",
			5236 => x"00fb51f1",
			5237 => x"ff6951f1",
			5238 => x"07002908",
			5239 => x"06004004",
			5240 => x"fee251f1",
			5241 => x"016351f1",
			5242 => x"fe3b51f1",
			5243 => x"fe6b51f1",
			5244 => x"04004760",
			5245 => x"00009e1c",
			5246 => x"08001604",
			5247 => x"feb252bd",
			5248 => x"06005510",
			5249 => x"0b001204",
			5250 => x"016252bd",
			5251 => x"04001204",
			5252 => x"fe8852bd",
			5253 => x"00008304",
			5254 => x"009e52bd",
			5255 => x"ff3652bd",
			5256 => x"0c001804",
			5257 => x"004952bd",
			5258 => x"016752bd",
			5259 => x"0e005a14",
			5260 => x"0000ae10",
			5261 => x"0000a90c",
			5262 => x"08001b04",
			5263 => x"005b52bd",
			5264 => x"0d001704",
			5265 => x"fe8a52bd",
			5266 => x"00d452bd",
			5267 => x"00bd52bd",
			5268 => x"fe3c52bd",
			5269 => x"05003718",
			5270 => x"0300240c",
			5271 => x"09001c08",
			5272 => x"0200aa04",
			5273 => x"006d52bd",
			5274 => x"fe9852bd",
			5275 => x"013e52bd",
			5276 => x"04001b08",
			5277 => x"0f00ad04",
			5278 => x"00b352bd",
			5279 => x"ff2652bd",
			5280 => x"fe5352bd",
			5281 => x"0200bb0c",
			5282 => x"0d001404",
			5283 => x"003752bd",
			5284 => x"06006604",
			5285 => x"00c952bd",
			5286 => x"019552bd",
			5287 => x"0f008804",
			5288 => x"fe6b52bd",
			5289 => x"01000904",
			5290 => x"011c52bd",
			5291 => x"ff2452bd",
			5292 => x"07002f04",
			5293 => x"012c52bd",
			5294 => x"fefa52bd",
			5295 => x"07003054",
			5296 => x"0400454c",
			5297 => x"03003530",
			5298 => x"09001f20",
			5299 => x"04002510",
			5300 => x"08001b08",
			5301 => x"0c001104",
			5302 => x"00905369",
			5303 => x"feda5369",
			5304 => x"0a002c04",
			5305 => x"00815369",
			5306 => x"ff2d5369",
			5307 => x"07002508",
			5308 => x"0f005304",
			5309 => x"002e5369",
			5310 => x"ff375369",
			5311 => x"02010204",
			5312 => x"012d5369",
			5313 => x"ffcc5369",
			5314 => x"0b001704",
			5315 => x"00625369",
			5316 => x"0000a108",
			5317 => x"02008e04",
			5318 => x"ff3f5369",
			5319 => x"005a5369",
			5320 => x"fed05369",
			5321 => x"0d00140c",
			5322 => x"04003604",
			5323 => x"febb5369",
			5324 => x"0000b204",
			5325 => x"000e5369",
			5326 => x"ff0c5369",
			5327 => x"08001c08",
			5328 => x"06006504",
			5329 => x"ff6c5369",
			5330 => x"008d5369",
			5331 => x"0000c604",
			5332 => x"011d5369",
			5333 => x"ff5a5369",
			5334 => x"03004704",
			5335 => x"00eb5369",
			5336 => x"ffee5369",
			5337 => x"ff1c5369",
			5338 => x"0700304c",
			5339 => x"04004748",
			5340 => x"00009e20",
			5341 => x"08001b0c",
			5342 => x"0c001104",
			5343 => x"00f65405",
			5344 => x"05002d04",
			5345 => x"fe8b5405",
			5346 => x"ffe45405",
			5347 => x"06005510",
			5348 => x"0b001508",
			5349 => x"05001804",
			5350 => x"00525405",
			5351 => x"01325405",
			5352 => x"08001f04",
			5353 => x"feeb5405",
			5354 => x"008f5405",
			5355 => x"01455405",
			5356 => x"0e005a14",
			5357 => x"0000ad10",
			5358 => x"0e005108",
			5359 => x"0d001704",
			5360 => x"fe655405",
			5361 => x"00785405",
			5362 => x"04003404",
			5363 => x"ff435405",
			5364 => x"009b5405",
			5365 => x"fe545405",
			5366 => x"0200a604",
			5367 => x"01515405",
			5368 => x"05002808",
			5369 => x"07002e04",
			5370 => x"fe675405",
			5371 => x"007a5405",
			5372 => x"07002904",
			5373 => x"00d65405",
			5374 => x"ffa15405",
			5375 => x"00ec5405",
			5376 => x"fea05405",
			5377 => x"08001808",
			5378 => x"03001304",
			5379 => x"003b54c1",
			5380 => x"ff6054c1",
			5381 => x"07003054",
			5382 => x"01000b30",
			5383 => x"0400341c",
			5384 => x"0d00120c",
			5385 => x"04000e04",
			5386 => x"ffc654c1",
			5387 => x"07002904",
			5388 => x"008e54c1",
			5389 => x"ffe854c1",
			5390 => x"07002008",
			5391 => x"0c001704",
			5392 => x"005854c1",
			5393 => x"ffd054c1",
			5394 => x"0e007004",
			5395 => x"ff4254c1",
			5396 => x"002654c1",
			5397 => x"0c001804",
			5398 => x"ff9854c1",
			5399 => x"0c001a08",
			5400 => x"0a004304",
			5401 => x"00a554c1",
			5402 => x"ffad54c1",
			5403 => x"0a004204",
			5404 => x"ffb154c1",
			5405 => x"005354c1",
			5406 => x"0d001918",
			5407 => x"0500280c",
			5408 => x"0c001404",
			5409 => x"005854c1",
			5410 => x"0200a104",
			5411 => x"000554c1",
			5412 => x"ff7854c1",
			5413 => x"0a002f04",
			5414 => x"00e054c1",
			5415 => x"05003704",
			5416 => x"ffb054c1",
			5417 => x"005154c1",
			5418 => x"07002908",
			5419 => x"06003f04",
			5420 => x"fff554c1",
			5421 => x"004654c1",
			5422 => x"ff7954c1",
			5423 => x"ff7f54c1",
			5424 => x"06008d68",
			5425 => x"0c001a3c",
			5426 => x"0a004338",
			5427 => x"0000811c",
			5428 => x"0100070c",
			5429 => x"08001804",
			5430 => x"fe965597",
			5431 => x"0b001604",
			5432 => x"00975597",
			5433 => x"fedf5597",
			5434 => x"0e003908",
			5435 => x"0b001504",
			5436 => x"01615597",
			5437 => x"fe845597",
			5438 => x"05002b04",
			5439 => x"01365597",
			5440 => x"01e65597",
			5441 => x"0e004e0c",
			5442 => x"01000b08",
			5443 => x"01000604",
			5444 => x"002a5597",
			5445 => x"fe345597",
			5446 => x"013e5597",
			5447 => x"04002508",
			5448 => x"05002c04",
			5449 => x"008f5597",
			5450 => x"feab5597",
			5451 => x"03003904",
			5452 => x"012f5597",
			5453 => x"00055597",
			5454 => x"fe6f5597",
			5455 => x"03003a18",
			5456 => x"0e005610",
			5457 => x"0000a208",
			5458 => x"00009604",
			5459 => x"fe6b5597",
			5460 => x"00205597",
			5461 => x"0000ab04",
			5462 => x"fd0e5597",
			5463 => x"fe915597",
			5464 => x"06006304",
			5465 => x"00f45597",
			5466 => x"fdde5597",
			5467 => x"0000d010",
			5468 => x"0e00620c",
			5469 => x"0000b908",
			5470 => x"0a004504",
			5471 => x"01575597",
			5472 => x"009f5597",
			5473 => x"fe6d5597",
			5474 => x"01b15597",
			5475 => x"fe635597",
			5476 => x"fe705597",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1757, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3651, initial_addr_3'length));
	end generate gen_rom_7;

	gen_rom_8: if SELECT_ROM = 8 generate
		bank <= (
			0 => x"0400331c",
			1 => x"04002e10",
			2 => x"0500420c",
			3 => x"04002b04",
			4 => x"d95a0095",
			5 => x"01000a04",
			6 => x"db900095",
			7 => x"d95d0095",
			8 => x"db910095",
			9 => x"08001c04",
			10 => x"e36b0095",
			11 => x"0000f904",
			12 => x"da7c0095",
			13 => x"d95f0095",
			14 => x"0b001e24",
			15 => x"0000b514",
			16 => x"0d00140c",
			17 => x"07002504",
			18 => x"e92f0095",
			19 => x"0000a804",
			20 => x"e0f00095",
			21 => x"e42b0095",
			22 => x"07002904",
			23 => x"de990095",
			24 => x"d9640095",
			25 => x"01000d0c",
			26 => x"0a004508",
			27 => x"0d001404",
			28 => x"e9f10095",
			29 => x"e2b50095",
			30 => x"ea770095",
			31 => x"de7a0095",
			32 => x"0b001f04",
			33 => x"ddbb0095",
			34 => x"0b002004",
			35 => x"da5d0095",
			36 => x"d95b0095",
			37 => x"0e006b34",
			38 => x"0c001810",
			39 => x"0d001108",
			40 => x"01000704",
			41 => x"ff250129",
			42 => x"005d0129",
			43 => x"05003c04",
			44 => x"ff690129",
			45 => x"01370129",
			46 => x"00009e08",
			47 => x"08001904",
			48 => x"ffd20129",
			49 => x"fea20129",
			50 => x"0d001308",
			51 => x"09002004",
			52 => x"fed40129",
			53 => x"01140129",
			54 => x"0e005708",
			55 => x"0a003704",
			56 => x"ff280129",
			57 => x"01060129",
			58 => x"0000ae04",
			59 => x"fea20129",
			60 => x"0000c704",
			61 => x"ffeb0129",
			62 => x"01010129",
			63 => x"0c001b0c",
			64 => x"08001908",
			65 => x"08001804",
			66 => x"ff980129",
			67 => x"00120129",
			68 => x"fe930129",
			69 => x"01001008",
			70 => x"03006a04",
			71 => x"01040129",
			72 => x"ffc60129",
			73 => x"ff110129",
			74 => x"0000ed34",
			75 => x"0b001714",
			76 => x"04002b04",
			77 => x"ffbd01ad",
			78 => x"04003e0c",
			79 => x"05004908",
			80 => x"05004404",
			81 => x"009401ad",
			82 => x"ffba01ad",
			83 => x"00dd01ad",
			84 => x"ffea01ad",
			85 => x"02009704",
			86 => x"ff5601ad",
			87 => x"0000a808",
			88 => x"08001d04",
			89 => x"00a101ad",
			90 => x"fff601ad",
			91 => x"0c001908",
			92 => x"07002b04",
			93 => x"ff4f01ad",
			94 => x"004601ad",
			95 => x"0000ad04",
			96 => x"ff8e01ad",
			97 => x"0e006704",
			98 => x"007801ad",
			99 => x"ffbe01ad",
			100 => x"05005008",
			101 => x"03003d04",
			102 => x"ff6401ad",
			103 => x"000401ad",
			104 => x"0a005404",
			105 => x"003b01ad",
			106 => x"ffd001ad",
			107 => x"04002b04",
			108 => x"fe6201f9",
			109 => x"02010620",
			110 => x"0a005c1c",
			111 => x"0a004710",
			112 => x"07002504",
			113 => x"01b801f9",
			114 => x"02009704",
			115 => x"fe3101f9",
			116 => x"01000904",
			117 => x"00d001f9",
			118 => x"ffd201f9",
			119 => x"08001d04",
			120 => x"01be01f9",
			121 => x"06007804",
			122 => x"000401f9",
			123 => x"01de01f9",
			124 => x"fe7301f9",
			125 => x"fe5901f9",
			126 => x"0d001638",
			127 => x"06005c0c",
			128 => x"07002508",
			129 => x"05003c04",
			130 => x"ffea0285",
			131 => x"00480285",
			132 => x"ffa30285",
			133 => x"0e005c10",
			134 => x"0000a204",
			135 => x"ffdd0285",
			136 => x"0a003904",
			137 => x"ffe80285",
			138 => x"0a004204",
			139 => x"00970285",
			140 => x"ffed0285",
			141 => x"0200bb08",
			142 => x"05004804",
			143 => x"00050285",
			144 => x"ff940285",
			145 => x"0900200c",
			146 => x"0e006504",
			147 => x"00200285",
			148 => x"0b001704",
			149 => x"00110285",
			150 => x"ffb30285",
			151 => x"08001d04",
			152 => x"006f0285",
			153 => x"fff30285",
			154 => x"01000704",
			155 => x"00040285",
			156 => x"0f008104",
			157 => x"ffb40285",
			158 => x"02010304",
			159 => x"001e0285",
			160 => x"ffda0285",
			161 => x"05003c04",
			162 => x"fe9102f9",
			163 => x"0d00151c",
			164 => x"03003508",
			165 => x"03003204",
			166 => x"00a702f9",
			167 => x"fef102f9",
			168 => x"0100090c",
			169 => x"0f006404",
			170 => x"006d02f9",
			171 => x"0c001804",
			172 => x"003e02f9",
			173 => x"019802f9",
			174 => x"0000b904",
			175 => x"ffef02f9",
			176 => x"012702f9",
			177 => x"0b001908",
			178 => x"08001b04",
			179 => x"ffd302f9",
			180 => x"fe6d02f9",
			181 => x"04003604",
			182 => x"fec002f9",
			183 => x"03003d04",
			184 => x"017c02f9",
			185 => x"0200b904",
			186 => x"fe9902f9",
			187 => x"01000b04",
			188 => x"014902f9",
			189 => x"ffac02f9",
			190 => x"0e00653c",
			191 => x"0000a218",
			192 => x"09001d08",
			193 => x"05003c04",
			194 => x"ffe903bd",
			195 => x"004c03bd",
			196 => x"0c001808",
			197 => x"0e004904",
			198 => x"001103bd",
			199 => x"ffff03bd",
			200 => x"08001904",
			201 => x"000303bd",
			202 => x"ff8b03bd",
			203 => x"0500450c",
			204 => x"06006908",
			205 => x"03003104",
			206 => x"000603bd",
			207 => x"ffc403bd",
			208 => x"001103bd",
			209 => x"0d00170c",
			210 => x"07002c08",
			211 => x"04003704",
			212 => x"001203bd",
			213 => x"007e03bd",
			214 => x"fff103bd",
			215 => x"0200b904",
			216 => x"ffd203bd",
			217 => x"04006604",
			218 => x"001c03bd",
			219 => x"fff603bd",
			220 => x"0000d608",
			221 => x"07003004",
			222 => x"ff9303bd",
			223 => x"000403bd",
			224 => x"0000fa10",
			225 => x"03003508",
			226 => x"0200d804",
			227 => x"001703bd",
			228 => x"ffdd03bd",
			229 => x"03005c04",
			230 => x"006703bd",
			231 => x"fff403bd",
			232 => x"05005008",
			233 => x"03003d04",
			234 => x"ffb903bd",
			235 => x"000203bd",
			236 => x"03005304",
			237 => x"001403bd",
			238 => x"ffef03bd",
			239 => x"05003c04",
			240 => x"fe5c0419",
			241 => x"01001024",
			242 => x"03005c20",
			243 => x"0a004514",
			244 => x"07002508",
			245 => x"03003304",
			246 => x"02a00419",
			247 => x"01df0419",
			248 => x"02009704",
			249 => x"fedd0419",
			250 => x"0d001704",
			251 => x"01340419",
			252 => x"ff7a0419",
			253 => x"05006508",
			254 => x"08001d04",
			255 => x"02040419",
			256 => x"00f70419",
			257 => x"027e0419",
			258 => x"fe670419",
			259 => x"08002204",
			260 => x"ff730419",
			261 => x"fe570419",
			262 => x"08001d3c",
			263 => x"0a004534",
			264 => x"0600641c",
			265 => x"05004510",
			266 => x"0b001608",
			267 => x"05003c04",
			268 => x"ffdc04bd",
			269 => x"007104bd",
			270 => x"09001c04",
			271 => x"000404bd",
			272 => x"ff6804bd",
			273 => x"06005904",
			274 => x"fff204bd",
			275 => x"0d001404",
			276 => x"00b204bd",
			277 => x"003c04bd",
			278 => x"0200bb08",
			279 => x"0d001304",
			280 => x"001504bd",
			281 => x"ff2504bd",
			282 => x"0900200c",
			283 => x"06007804",
			284 => x"001b04bd",
			285 => x"01000504",
			286 => x"001404bd",
			287 => x"ff5204bd",
			288 => x"008c04bd",
			289 => x"09002504",
			290 => x"00c504bd",
			291 => x"fffb04bd",
			292 => x"09001f08",
			293 => x"0a003604",
			294 => x"ffe704bd",
			295 => x"004f04bd",
			296 => x"05005e08",
			297 => x"03004604",
			298 => x"ff3f04bd",
			299 => x"fff904bd",
			300 => x"0a005904",
			301 => x"004704bd",
			302 => x"ffc304bd",
			303 => x"04002b04",
			304 => x"fe650519",
			305 => x"02010124",
			306 => x"0a005c20",
			307 => x"07002f18",
			308 => x"0d001710",
			309 => x"0e006508",
			310 => x"0000b404",
			311 => x"00570519",
			312 => x"01540519",
			313 => x"04003c04",
			314 => x"00a90519",
			315 => x"ff070519",
			316 => x"0200b904",
			317 => x"fe340519",
			318 => x"fff10519",
			319 => x"06007404",
			320 => x"012e0519",
			321 => x"01bd0519",
			322 => x"fe7f0519",
			323 => x"05005204",
			324 => x"fe590519",
			325 => x"00750519",
			326 => x"08001f40",
			327 => x"0a003614",
			328 => x"07002508",
			329 => x"05003b04",
			330 => x"ffb105ad",
			331 => x"008605ad",
			332 => x"09002004",
			333 => x"ff2305ad",
			334 => x"09002104",
			335 => x"000a05ad",
			336 => x"fffb05ad",
			337 => x"0a004218",
			338 => x"0d001714",
			339 => x"0f006308",
			340 => x"01000804",
			341 => x"ff6d05ad",
			342 => x"007d05ad",
			343 => x"08001804",
			344 => x"ffba05ad",
			345 => x"0a003b04",
			346 => x"000f05ad",
			347 => x"00ef05ad",
			348 => x"ff9605ad",
			349 => x"0a004304",
			350 => x"ff4605ad",
			351 => x"01000404",
			352 => x"ff8305ad",
			353 => x"0000be04",
			354 => x"ffef05ad",
			355 => x"03005504",
			356 => x"00da05ad",
			357 => x"ffea05ad",
			358 => x"04004a04",
			359 => x"ff3205ad",
			360 => x"05008104",
			361 => x"003d05ad",
			362 => x"ffc105ad",
			363 => x"01000938",
			364 => x"08001b1c",
			365 => x"05004918",
			366 => x"07002910",
			367 => x"07002308",
			368 => x"09001a04",
			369 => x"fff00661",
			370 => x"00260661",
			371 => x"06005f04",
			372 => x"ff9c0661",
			373 => x"ffff0661",
			374 => x"0000f204",
			375 => x"004c0661",
			376 => x"ffe50661",
			377 => x"00be0661",
			378 => x"05004d14",
			379 => x"0f00640c",
			380 => x"01000808",
			381 => x"08001c04",
			382 => x"000b0661",
			383 => x"ffb60661",
			384 => x"00260661",
			385 => x"05004204",
			386 => x"fff60661",
			387 => x"007f0661",
			388 => x"0c001b04",
			389 => x"ff8a0661",
			390 => x"002a0661",
			391 => x"09001e08",
			392 => x"05003f04",
			393 => x"ffd70661",
			394 => x"006e0661",
			395 => x"04004314",
			396 => x"0000c704",
			397 => x"ff350661",
			398 => x"0201030c",
			399 => x"03003a08",
			400 => x"0000dd04",
			401 => x"00050661",
			402 => x"ffe90661",
			403 => x"00460661",
			404 => x"ffce0661",
			405 => x"0a005904",
			406 => x"004f0661",
			407 => x"ffd40661",
			408 => x"0d001538",
			409 => x"05004924",
			410 => x"0d001310",
			411 => x"07002308",
			412 => x"05003c04",
			413 => x"ffee072d",
			414 => x"002a072d",
			415 => x"07002c04",
			416 => x"ff98072d",
			417 => x"0001072d",
			418 => x"00009e0c",
			419 => x"0e004b08",
			420 => x"07002204",
			421 => x"0000072d",
			422 => x"000e072d",
			423 => x"ffdb072d",
			424 => x"04002d04",
			425 => x"ffed072d",
			426 => x"004f072d",
			427 => x"0d00140c",
			428 => x"04003e04",
			429 => x"007c072d",
			430 => x"01000704",
			431 => x"ffdf072d",
			432 => x"001e072d",
			433 => x"08001b04",
			434 => x"0018072d",
			435 => x"ffe2072d",
			436 => x"06006208",
			437 => x"0c001604",
			438 => x"ffff072d",
			439 => x"ff84072d",
			440 => x"0b00190c",
			441 => x"0b001708",
			442 => x"06008704",
			443 => x"000f072d",
			444 => x"fff6072d",
			445 => x"ffb1072d",
			446 => x"04004b0c",
			447 => x"08002208",
			448 => x"0a003b04",
			449 => x"fff0072d",
			450 => x"007f072d",
			451 => x"ffe1072d",
			452 => x"0e007108",
			453 => x"01000a04",
			454 => x"000a072d",
			455 => x"ffc3072d",
			456 => x"07003c04",
			457 => x"001b072d",
			458 => x"fffa072d",
			459 => x"08001d3c",
			460 => x"0a003614",
			461 => x"0700240c",
			462 => x"07002004",
			463 => x"ffe207d1",
			464 => x"09001a04",
			465 => x"fffd07d1",
			466 => x"002607d1",
			467 => x"09002004",
			468 => x"ff8107d1",
			469 => x"000d07d1",
			470 => x"0d001720",
			471 => x"09002118",
			472 => x"01000810",
			473 => x"03003b08",
			474 => x"0a003b04",
			475 => x"006207d1",
			476 => x"ff7307d1",
			477 => x"04003e04",
			478 => x"00ad07d1",
			479 => x"fff107d1",
			480 => x"06006404",
			481 => x"00bc07d1",
			482 => x"fffb07d1",
			483 => x"0200bc04",
			484 => x"ff8f07d1",
			485 => x"008f07d1",
			486 => x"03004104",
			487 => x"ffa607d1",
			488 => x"000e07d1",
			489 => x"0d001304",
			490 => x"002407d1",
			491 => x"0f007204",
			492 => x"ff5207d1",
			493 => x"0e006504",
			494 => x"007007d1",
			495 => x"05005e04",
			496 => x"ff9207d1",
			497 => x"05008104",
			498 => x"001107d1",
			499 => x"ffe507d1",
			500 => x"04002b04",
			501 => x"fe5d0835",
			502 => x"01001028",
			503 => x"04006624",
			504 => x"0a004514",
			505 => x"07002508",
			506 => x"0a003604",
			507 => x"025b0835",
			508 => x"01d70835",
			509 => x"02009704",
			510 => x"fef00835",
			511 => x"0000ed04",
			512 => x"010d0835",
			513 => x"ff520835",
			514 => x"0200cc08",
			515 => x"08001c04",
			516 => x"01f50835",
			517 => x"004e0835",
			518 => x"07003604",
			519 => x"01e10835",
			520 => x"02540835",
			521 => x"fe680835",
			522 => x"08002204",
			523 => x"ffa80835",
			524 => x"fe5a0835",
			525 => x"05003c04",
			526 => x"fe630889",
			527 => x"02010624",
			528 => x"0b002020",
			529 => x"0a004818",
			530 => x"09001d08",
			531 => x"05004404",
			532 => x"01700889",
			533 => x"022e0889",
			534 => x"0000b408",
			535 => x"04003804",
			536 => x"fec40889",
			537 => x"00410889",
			538 => x"0e006304",
			539 => x"01520889",
			540 => x"000a0889",
			541 => x"0f007204",
			542 => x"009e0889",
			543 => x"01b60889",
			544 => x"fe750889",
			545 => x"fe5d0889",
			546 => x"05003e04",
			547 => x"fe66091d",
			548 => x"08001d24",
			549 => x"0e005a10",
			550 => x"05004908",
			551 => x"09001d04",
			552 => x"0205091d",
			553 => x"ffbe091d",
			554 => x"0e005604",
			555 => x"023d091d",
			556 => x"010f091d",
			557 => x"0000be04",
			558 => x"fea9091d",
			559 => x"0e006204",
			560 => x"01aa091d",
			561 => x"07002c04",
			562 => x"fe85091d",
			563 => x"0200c904",
			564 => x"ff78091d",
			565 => x"0169091d",
			566 => x"05004f10",
			567 => x"0a003b08",
			568 => x"0a003904",
			569 => x"fe80091d",
			570 => x"00b8091d",
			571 => x"03004004",
			572 => x"fe2f091d",
			573 => x"ffcb091d",
			574 => x"0f007708",
			575 => x"04004904",
			576 => x"ffd4091d",
			577 => x"fe39091d",
			578 => x"0a005908",
			579 => x"0e007c04",
			580 => x"01a7091d",
			581 => x"00cb091d",
			582 => x"feb3091d",
			583 => x"04002b04",
			584 => x"fecf0999",
			585 => x"09001e0c",
			586 => x"05004708",
			587 => x"07002504",
			588 => x"00bc0999",
			589 => x"ff240999",
			590 => x"015f0999",
			591 => x"08001b10",
			592 => x"05004c08",
			593 => x"0000be04",
			594 => x"feff0999",
			595 => x"00be0999",
			596 => x"0c001b04",
			597 => x"01330999",
			598 => x"ffe80999",
			599 => x"01000808",
			600 => x"04003c04",
			601 => x"00010999",
			602 => x"fecf0999",
			603 => x"04003b0c",
			604 => x"0000b504",
			605 => x"fea10999",
			606 => x"04003404",
			607 => x"ff4a0999",
			608 => x"008c0999",
			609 => x"01000904",
			610 => x"01280999",
			611 => x"04004304",
			612 => x"ff350999",
			613 => x"00b00999",
			614 => x"0000ed44",
			615 => x"09001e0c",
			616 => x"05003c04",
			617 => x"ff9b0a3d",
			618 => x"0d001204",
			619 => x"00190a3d",
			620 => x"01000a3d",
			621 => x"0000b41c",
			622 => x"0e005514",
			623 => x"05004b10",
			624 => x"07002b08",
			625 => x"01000504",
			626 => x"004e0a3d",
			627 => x"fee90a3d",
			628 => x"01000c04",
			629 => x"005b0a3d",
			630 => x"fffb0a3d",
			631 => x"00cd0a3d",
			632 => x"05004704",
			633 => x"00470a3d",
			634 => x"fed40a3d",
			635 => x"0e005f0c",
			636 => x"0d001704",
			637 => x"010d0a3d",
			638 => x"07002c04",
			639 => x"ffa80a3d",
			640 => x"00300a3d",
			641 => x"0000c704",
			642 => x"ff210a3d",
			643 => x"07002b04",
			644 => x"ffaf0a3d",
			645 => x"0d001804",
			646 => x"01160a3d",
			647 => x"ffe70a3d",
			648 => x"05005008",
			649 => x"03003d04",
			650 => x"ff1e0a3d",
			651 => x"00020a3d",
			652 => x"03005304",
			653 => x"00370a3d",
			654 => x"ffc70a3d",
			655 => x"04002b04",
			656 => x"fe650aa1",
			657 => x"0800232c",
			658 => x"05004914",
			659 => x"07002508",
			660 => x"08001904",
			661 => x"01120aa1",
			662 => x"01c60aa1",
			663 => x"0d001304",
			664 => x"fe610aa1",
			665 => x"0000ae04",
			666 => x"ff690aa1",
			667 => x"00ee0aa1",
			668 => x"0e005704",
			669 => x"01cd0aa1",
			670 => x"0000b204",
			671 => x"fe550aa1",
			672 => x"0e005f08",
			673 => x"05005404",
			674 => x"01e00aa1",
			675 => x"013c0aa1",
			676 => x"0000c704",
			677 => x"fe640aa1",
			678 => x"010a0aa1",
			679 => x"fe850aa1",
			680 => x"0200ee4c",
			681 => x"0000c724",
			682 => x"06006a1c",
			683 => x"09001d08",
			684 => x"05003c04",
			685 => x"ff320b4d",
			686 => x"01960b4d",
			687 => x"0000b50c",
			688 => x"0e005a08",
			689 => x"02009804",
			690 => x"ff420b4d",
			691 => x"00760b4d",
			692 => x"fe820b4d",
			693 => x"06005f04",
			694 => x"ff040b4d",
			695 => x"013b0b4d",
			696 => x"0d001304",
			697 => x"ffe90b4d",
			698 => x"fe760b4d",
			699 => x"0000dd14",
			700 => x"0d001808",
			701 => x"04002d04",
			702 => x"ffa20b4d",
			703 => x"01990b4d",
			704 => x"01000b04",
			705 => x"00ad0b4d",
			706 => x"07003204",
			707 => x"ff030b4d",
			708 => x"00010b4d",
			709 => x"07002b04",
			710 => x"fe960b4d",
			711 => x"0300590c",
			712 => x"01001008",
			713 => x"04003104",
			714 => x"ffd20b4d",
			715 => x"01660b4d",
			716 => x"ffaf0b4d",
			717 => x"ff4a0b4d",
			718 => x"03003d04",
			719 => x"fe890b4d",
			720 => x"01001004",
			721 => x"00dc0b4d",
			722 => x"ff200b4d",
			723 => x"0400310c",
			724 => x"04002b04",
			725 => x"fe4b0bc1",
			726 => x"0000f104",
			727 => x"02db0bc1",
			728 => x"fe490bc1",
			729 => x"0d001b2c",
			730 => x"04006128",
			731 => x"0500490c",
			732 => x"07002504",
			733 => x"03fe0bc1",
			734 => x"0f006704",
			735 => x"fe8e0bc1",
			736 => x"02470bc1",
			737 => x"0000b90c",
			738 => x"01000908",
			739 => x"08001b04",
			740 => x"04970bc1",
			741 => x"02b00bc1",
			742 => x"ffbe0bc1",
			743 => x"09002308",
			744 => x"0e006204",
			745 => x"03eb0bc1",
			746 => x"02ac0bc1",
			747 => x"01000c04",
			748 => x"03ca0bc1",
			749 => x"04e90bc1",
			750 => x"fe4e0bc1",
			751 => x"fe4c0bc1",
			752 => x"0500410c",
			753 => x"05003c04",
			754 => x"fe410c4d",
			755 => x"0000df04",
			756 => x"03710c4d",
			757 => x"fe3e0c4d",
			758 => x"0d001b30",
			759 => x"03005c2c",
			760 => x"0000b414",
			761 => x"0c001808",
			762 => x"0b001504",
			763 => x"08790c4d",
			764 => x"05c70c4d",
			765 => x"0d001404",
			766 => x"03a10c4d",
			767 => x"07002904",
			768 => x"00dd0c4d",
			769 => x"fe470c4d",
			770 => x"01000c10",
			771 => x"0200b908",
			772 => x"0e005b04",
			773 => x"07390c4d",
			774 => x"02920c4d",
			775 => x"09002004",
			776 => x"05bb0c4d",
			777 => x"06f60c4d",
			778 => x"05005204",
			779 => x"02e20c4d",
			780 => x"05d80c4d",
			781 => x"fe4b0c4d",
			782 => x"0b001f08",
			783 => x"0600ac04",
			784 => x"002d0c4d",
			785 => x"fe460c4d",
			786 => x"fe420c4d",
			787 => x"04002b04",
			788 => x"fe720cd9",
			789 => x"0b001714",
			790 => x"0500490c",
			791 => x"03003304",
			792 => x"014e0cd9",
			793 => x"0a003b04",
			794 => x"005e0cd9",
			795 => x"ff150cd9",
			796 => x"07002904",
			797 => x"01c50cd9",
			798 => x"00b70cd9",
			799 => x"05004f14",
			800 => x"0000ae04",
			801 => x"fe5b0cd9",
			802 => x"0e005b04",
			803 => x"01350cd9",
			804 => x"07002c04",
			805 => x"fedc0cd9",
			806 => x"0a004204",
			807 => x"00e50cd9",
			808 => x"fe8c0cd9",
			809 => x"09002108",
			810 => x"0f006f04",
			811 => x"01650cd9",
			812 => x"00660cd9",
			813 => x"0f00810c",
			814 => x"0e006808",
			815 => x"0200b904",
			816 => x"ff010cd9",
			817 => x"00fc0cd9",
			818 => x"fe310cd9",
			819 => x"01001004",
			820 => x"01740cd9",
			821 => x"feff0cd9",
			822 => x"0d001534",
			823 => x"03003920",
			824 => x"07002508",
			825 => x"05003c04",
			826 => x"ffd90dad",
			827 => x"00870dad",
			828 => x"0000b50c",
			829 => x"09001d04",
			830 => x"003e0dad",
			831 => x"0c001b04",
			832 => x"ff360dad",
			833 => x"001f0dad",
			834 => x"0000df08",
			835 => x"04002d04",
			836 => x"fff80dad",
			837 => x"008a0dad",
			838 => x"ff940dad",
			839 => x"0900210c",
			840 => x"0e005d04",
			841 => x"00c70dad",
			842 => x"06006d04",
			843 => x"ffed0dad",
			844 => x"00440dad",
			845 => x"08001b04",
			846 => x"00420dad",
			847 => x"ffaf0dad",
			848 => x"01000708",
			849 => x"08001d04",
			850 => x"007c0dad",
			851 => x"ffc40dad",
			852 => x"0a004724",
			853 => x"02009c10",
			854 => x"0700290c",
			855 => x"07002808",
			856 => x"09001d04",
			857 => x"001f0dad",
			858 => x"ffda0dad",
			859 => x"005d0dad",
			860 => x"ffda0dad",
			861 => x"0b001608",
			862 => x"09001e04",
			863 => x"fff40dad",
			864 => x"00130dad",
			865 => x"06007604",
			866 => x"ff0c0dad",
			867 => x"09002104",
			868 => x"ffc50dad",
			869 => x"00190dad",
			870 => x"0a005908",
			871 => x"0f00a204",
			872 => x"006a0dad",
			873 => x"fffe0dad",
			874 => x"ffc30dad",
			875 => x"0b001720",
			876 => x"05004918",
			877 => x"07002508",
			878 => x"05003c04",
			879 => x"ffc20e79",
			880 => x"00a70e79",
			881 => x"0200ad04",
			882 => x"ff280e79",
			883 => x"0200e208",
			884 => x"03002904",
			885 => x"ffeb0e79",
			886 => x"00a10e79",
			887 => x"ff990e79",
			888 => x"05004f04",
			889 => x"00d40e79",
			890 => x"00040e79",
			891 => x"05005124",
			892 => x"0000ae0c",
			893 => x"09001d04",
			894 => x"00680e79",
			895 => x"03003d04",
			896 => x"fef00e79",
			897 => x"00040e79",
			898 => x"0e005b08",
			899 => x"0200ba04",
			900 => x"00eb0e79",
			901 => x"ffc20e79",
			902 => x"0f007c04",
			903 => x"ff470e79",
			904 => x"03003a04",
			905 => x"ff620e79",
			906 => x"0a004204",
			907 => x"009a0e79",
			908 => x"ffe00e79",
			909 => x"09002108",
			910 => x"0e005d04",
			911 => x"00f30e79",
			912 => x"00020e79",
			913 => x"0200b904",
			914 => x"ff3c0e79",
			915 => x"0e00690c",
			916 => x"08001f04",
			917 => x"00ac0e79",
			918 => x"01000b04",
			919 => x"000d0e79",
			920 => x"ffbc0e79",
			921 => x"0f008104",
			922 => x"ff5a0e79",
			923 => x"0a005904",
			924 => x"00630e79",
			925 => x"ffe10e79",
			926 => x"0d001544",
			927 => x"05004930",
			928 => x"0d00131c",
			929 => x"07002308",
			930 => x"05003c04",
			931 => x"ffee0f5d",
			932 => x"00290f5d",
			933 => x"07002c0c",
			934 => x"05003d08",
			935 => x"05003404",
			936 => x"fff40f5d",
			937 => x"000c0f5d",
			938 => x"ff960f5d",
			939 => x"03002e04",
			940 => x"fffc0f5d",
			941 => x"00060f5d",
			942 => x"00009e0c",
			943 => x"0e004b08",
			944 => x"07002204",
			945 => x"00000f5d",
			946 => x"000d0f5d",
			947 => x"ffdb0f5d",
			948 => x"04002d04",
			949 => x"ffed0f5d",
			950 => x"004c0f5d",
			951 => x"0d00140c",
			952 => x"04003e04",
			953 => x"00780f5d",
			954 => x"01000704",
			955 => x"ffe00f5d",
			956 => x"001d0f5d",
			957 => x"08001b04",
			958 => x"00180f5d",
			959 => x"ffe40f5d",
			960 => x"06006208",
			961 => x"0c001604",
			962 => x"00000f5d",
			963 => x"ff890f5d",
			964 => x"0b00190c",
			965 => x"0b001708",
			966 => x"06008704",
			967 => x"000e0f5d",
			968 => x"fff60f5d",
			969 => x"ffb40f5d",
			970 => x"04004b0c",
			971 => x"08002208",
			972 => x"0a003b04",
			973 => x"fff00f5d",
			974 => x"007a0f5d",
			975 => x"ffe20f5d",
			976 => x"0e007108",
			977 => x"01000a04",
			978 => x"000a0f5d",
			979 => x"ffc50f5d",
			980 => x"07003c04",
			981 => x"001a0f5d",
			982 => x"fffa0f5d",
			983 => x"04002b04",
			984 => x"fe880fd1",
			985 => x"0000f528",
			986 => x"09001d04",
			987 => x"01820fd1",
			988 => x"02009808",
			989 => x"09001f04",
			990 => x"ffe10fd1",
			991 => x"fed60fd1",
			992 => x"0a00420c",
			993 => x"08001904",
			994 => x"ffb00fd1",
			995 => x"0d001704",
			996 => x"01080fd1",
			997 => x"ff530fd1",
			998 => x"0000d608",
			999 => x"0e006504",
			1000 => x"000d0fd1",
			1001 => x"fee20fd1",
			1002 => x"0f007804",
			1003 => x"ff3d0fd1",
			1004 => x"01560fd1",
			1005 => x"03003d04",
			1006 => x"fe990fd1",
			1007 => x"01000d04",
			1008 => x"01070fd1",
			1009 => x"0a004804",
			1010 => x"ffec0fd1",
			1011 => x"ff080fd1",
			1012 => x"05004114",
			1013 => x"04002e0c",
			1014 => x"05003e04",
			1015 => x"fe59105d",
			1016 => x"03003304",
			1017 => x"0018105d",
			1018 => x"fe5e105d",
			1019 => x"03003304",
			1020 => x"013b105d",
			1021 => x"fe31105d",
			1022 => x"0b002030",
			1023 => x"0201062c",
			1024 => x"05004f14",
			1025 => x"09001d04",
			1026 => x"02c1105d",
			1027 => x"0000b408",
			1028 => x"0e005a04",
			1029 => x"003a105d",
			1030 => x"fdfb105d",
			1031 => x"0b001704",
			1032 => x"02ab105d",
			1033 => x"00d6105d",
			1034 => x"0f008110",
			1035 => x"08001c08",
			1036 => x"0e005a04",
			1037 => x"029e105d",
			1038 => x"01f6105d",
			1039 => x"0000c504",
			1040 => x"ffad105d",
			1041 => x"015e105d",
			1042 => x"0d001904",
			1043 => x"0233105d",
			1044 => x"02d0105d",
			1045 => x"fe34105d",
			1046 => x"fe5d105d",
			1047 => x"0d00153c",
			1048 => x"03003928",
			1049 => x"07002508",
			1050 => x"05003c04",
			1051 => x"ffda1139",
			1052 => x"00841139",
			1053 => x"0700280c",
			1054 => x"09001d08",
			1055 => x"0e006b04",
			1056 => x"00381139",
			1057 => x"fffb1139",
			1058 => x"ff401139",
			1059 => x"0000df10",
			1060 => x"0200a608",
			1061 => x"06005d04",
			1062 => x"001d1139",
			1063 => x"ffb01139",
			1064 => x"03002f04",
			1065 => x"fffb1139",
			1066 => x"00951139",
			1067 => x"ff9d1139",
			1068 => x"0900210c",
			1069 => x"0e005d04",
			1070 => x"00b81139",
			1071 => x"06006d04",
			1072 => x"ffee1139",
			1073 => x"003f1139",
			1074 => x"08001b04",
			1075 => x"00411139",
			1076 => x"ffb21139",
			1077 => x"01000708",
			1078 => x"08001d04",
			1079 => x"00771139",
			1080 => x"ffc71139",
			1081 => x"0a004720",
			1082 => x"02009c0c",
			1083 => x"07002908",
			1084 => x"00008f04",
			1085 => x"fff41139",
			1086 => x"00551139",
			1087 => x"ffdb1139",
			1088 => x"0b001608",
			1089 => x"09001e04",
			1090 => x"fff51139",
			1091 => x"00131139",
			1092 => x"06007604",
			1093 => x"ff171139",
			1094 => x"06008a04",
			1095 => x"00181139",
			1096 => x"ffc71139",
			1097 => x"0a005908",
			1098 => x"0f00a204",
			1099 => x"00661139",
			1100 => x"ffff1139",
			1101 => x"ffc51139",
			1102 => x"08001d40",
			1103 => x"0a003614",
			1104 => x"0700240c",
			1105 => x"07002004",
			1106 => x"ffe311f5",
			1107 => x"09001a04",
			1108 => x"fffd11f5",
			1109 => x"002611f5",
			1110 => x"09002004",
			1111 => x"ff8611f5",
			1112 => x"000d11f5",
			1113 => x"0d001724",
			1114 => x"0b00170c",
			1115 => x"08001604",
			1116 => x"ffe711f5",
			1117 => x"00010104",
			1118 => x"00a711f5",
			1119 => x"ffef11f5",
			1120 => x"05005210",
			1121 => x"0e005b08",
			1122 => x"0c001904",
			1123 => x"ffe111f5",
			1124 => x"007a11f5",
			1125 => x"0000d004",
			1126 => x"ff7111f5",
			1127 => x"fff911f5",
			1128 => x"08001b04",
			1129 => x"00b511f5",
			1130 => x"000411f5",
			1131 => x"03004104",
			1132 => x"ffaa11f5",
			1133 => x"000e11f5",
			1134 => x"0d001304",
			1135 => x"002511f5",
			1136 => x"0f007204",
			1137 => x"ff5a11f5",
			1138 => x"0e006504",
			1139 => x"006b11f5",
			1140 => x"05005e0c",
			1141 => x"0c001e04",
			1142 => x"ff8a11f5",
			1143 => x"0c001f04",
			1144 => x"001811f5",
			1145 => x"fff111f5",
			1146 => x"0c002104",
			1147 => x"001c11f5",
			1148 => x"ffdd11f5",
			1149 => x"05003c04",
			1150 => x"fe5f1261",
			1151 => x"0100102c",
			1152 => x"03005c28",
			1153 => x"0a00481c",
			1154 => x"0d00150c",
			1155 => x"0000f208",
			1156 => x"09001d04",
			1157 => x"02651261",
			1158 => x"01211261",
			1159 => x"ff1f1261",
			1160 => x"0b001908",
			1161 => x"05004b04",
			1162 => x"ff991261",
			1163 => x"fe241261",
			1164 => x"0000d204",
			1165 => x"ffd71261",
			1166 => x"01c61261",
			1167 => x"0000ca04",
			1168 => x"014e1261",
			1169 => x"05006504",
			1170 => x"01d31261",
			1171 => x"023b1261",
			1172 => x"fe6d1261",
			1173 => x"07003104",
			1174 => x"00191261",
			1175 => x"fe5a1261",
			1176 => x"04002b04",
			1177 => x"fe6d12f5",
			1178 => x"0e00652c",
			1179 => x"0d001514",
			1180 => x"0000b20c",
			1181 => x"07002708",
			1182 => x"08001b04",
			1183 => x"007512f5",
			1184 => x"01d412f5",
			1185 => x"ff2f12f5",
			1186 => x"09001f04",
			1187 => x"00c912f5",
			1188 => x"01b512f5",
			1189 => x"04003c08",
			1190 => x"04003204",
			1191 => x"ffc212f5",
			1192 => x"fe6212f5",
			1193 => x"03003e04",
			1194 => x"015612f5",
			1195 => x"0200ba04",
			1196 => x"fe4012f5",
			1197 => x"0f006f04",
			1198 => x"ff0f12f5",
			1199 => x"017412f5",
			1200 => x"07002b04",
			1201 => x"fdda12f5",
			1202 => x"0000d604",
			1203 => x"feff12f5",
			1204 => x"0001100c",
			1205 => x"0c002208",
			1206 => x"0000f504",
			1207 => x"01af12f5",
			1208 => x"00bb12f5",
			1209 => x"fec712f5",
			1210 => x"05004f04",
			1211 => x"fe8812f5",
			1212 => x"ff9512f5",
			1213 => x"04002b04",
			1214 => x"fe6e1379",
			1215 => x"0d001520",
			1216 => x"0200d81c",
			1217 => x"0f007c18",
			1218 => x"0700270c",
			1219 => x"03003908",
			1220 => x"04003404",
			1221 => x"01931379",
			1222 => x"ffe91379",
			1223 => x"01f81379",
			1224 => x"0000b204",
			1225 => x"ff3b1379",
			1226 => x"0e006104",
			1227 => x"01a51379",
			1228 => x"ff601379",
			1229 => x"01b61379",
			1230 => x"ff021379",
			1231 => x"0b001908",
			1232 => x"08001c04",
			1233 => x"ff311379",
			1234 => x"fdf81379",
			1235 => x"0a003b04",
			1236 => x"fe7a1379",
			1237 => x"03003b08",
			1238 => x"04003504",
			1239 => x"fee01379",
			1240 => x"02651379",
			1241 => x"0000c304",
			1242 => x"fe4c1379",
			1243 => x"0d001b04",
			1244 => x"00f51379",
			1245 => x"fecf1379",
			1246 => x"04002b04",
			1247 => x"fea0140d",
			1248 => x"08001d2c",
			1249 => x"0a004524",
			1250 => x"06006414",
			1251 => x"01000808",
			1252 => x"0e005204",
			1253 => x"ff64140d",
			1254 => x"007f140d",
			1255 => x"09001e04",
			1256 => x"0167140d",
			1257 => x"06006004",
			1258 => x"003b140d",
			1259 => x"00e8140d",
			1260 => x"0000be04",
			1261 => x"fe98140d",
			1262 => x"0000e108",
			1263 => x"05005004",
			1264 => x"017b140d",
			1265 => x"ffa8140d",
			1266 => x"ff2e140d",
			1267 => x"09002504",
			1268 => x"0168140d",
			1269 => x"0031140d",
			1270 => x"0c001a04",
			1271 => x"0029140d",
			1272 => x"05005e0c",
			1273 => x"07003304",
			1274 => x"fe95140d",
			1275 => x"00011204",
			1276 => x"0089140d",
			1277 => x"ff4d140d",
			1278 => x"0a005904",
			1279 => x"00bb140d",
			1280 => x"0d001b04",
			1281 => x"fff4140d",
			1282 => x"ff38140d",
			1283 => x"0b001714",
			1284 => x"0500490c",
			1285 => x"05004408",
			1286 => x"05003c04",
			1287 => x"ff8a14b9",
			1288 => x"009114b9",
			1289 => x"ff8814b9",
			1290 => x"05004f04",
			1291 => x"00c814b9",
			1292 => x"000514b9",
			1293 => x"08001804",
			1294 => x"005a14b9",
			1295 => x"0c001914",
			1296 => x"09001d04",
			1297 => x"005b14b9",
			1298 => x"07002c08",
			1299 => x"0f005c04",
			1300 => x"ffe314b9",
			1301 => x"ff0b14b9",
			1302 => x"06009d04",
			1303 => x"005914b9",
			1304 => x"fff314b9",
			1305 => x"03003b10",
			1306 => x"0400390c",
			1307 => x"0b001808",
			1308 => x"0f006d04",
			1309 => x"fff814b9",
			1310 => x"005e14b9",
			1311 => x"ff5714b9",
			1312 => x"00de14b9",
			1313 => x"07002f0c",
			1314 => x"0a004808",
			1315 => x"04003c04",
			1316 => x"002814b9",
			1317 => x"ff2814b9",
			1318 => x"003014b9",
			1319 => x"0d001b08",
			1320 => x"03005c04",
			1321 => x"008c14b9",
			1322 => x"fff014b9",
			1323 => x"0000e704",
			1324 => x"000f14b9",
			1325 => x"ffb514b9",
			1326 => x"0200ee54",
			1327 => x"0500513c",
			1328 => x"0a004234",
			1329 => x"08001918",
			1330 => x"07002b10",
			1331 => x"0b001508",
			1332 => x"0d001004",
			1333 => x"ff6a1575",
			1334 => x"00c91575",
			1335 => x"09001d04",
			1336 => x"004e1575",
			1337 => x"fece1575",
			1338 => x"0000cc04",
			1339 => x"fff61575",
			1340 => x"00f01575",
			1341 => x"0000ae0c",
			1342 => x"07002708",
			1343 => x"05004604",
			1344 => x"ff651575",
			1345 => x"01021575",
			1346 => x"fe871575",
			1347 => x"0e005b08",
			1348 => x"0000c404",
			1349 => x"01911575",
			1350 => x"ffc01575",
			1351 => x"0000c404",
			1352 => x"ff291575",
			1353 => x"01011575",
			1354 => x"08001b04",
			1355 => x"00881575",
			1356 => x"fe7a1575",
			1357 => x"08001c0c",
			1358 => x"09002104",
			1359 => x"01851575",
			1360 => x"06007004",
			1361 => x"ffe81575",
			1362 => x"00c51575",
			1363 => x"0000c504",
			1364 => x"fec11575",
			1365 => x"03005c04",
			1366 => x"010a1575",
			1367 => x"ff6a1575",
			1368 => x"03003d04",
			1369 => x"fea81575",
			1370 => x"01001004",
			1371 => x"00bb1575",
			1372 => x"ff5c1575",
			1373 => x"0e00653c",
			1374 => x"09001e18",
			1375 => x"05004514",
			1376 => x"07002510",
			1377 => x"05003e0c",
			1378 => x"0c001508",
			1379 => x"05002904",
			1380 => x"ff9b1669",
			1381 => x"005e1669",
			1382 => x"ff621669",
			1383 => x"011f1669",
			1384 => x"ff0e1669",
			1385 => x"01731669",
			1386 => x"06005704",
			1387 => x"febe1669",
			1388 => x"0200b914",
			1389 => x"0600640c",
			1390 => x"08001d08",
			1391 => x"0c001904",
			1392 => x"ffee1669",
			1393 => x"00f01669",
			1394 => x"fec01669",
			1395 => x"01000904",
			1396 => x"ffbe1669",
			1397 => x"fea81669",
			1398 => x"0b001c08",
			1399 => x"0200c904",
			1400 => x"01651669",
			1401 => x"00311669",
			1402 => x"ff7c1669",
			1403 => x"07002b0c",
			1404 => x"03003108",
			1405 => x"03002c04",
			1406 => x"ff9c1669",
			1407 => x"00a31669",
			1408 => x"fe7f1669",
			1409 => x"08001d1c",
			1410 => x"0000cd04",
			1411 => x"fedb1669",
			1412 => x"0200ee0c",
			1413 => x"04004308",
			1414 => x"03003104",
			1415 => x"fff51669",
			1416 => x"01671669",
			1417 => x"fffe1669",
			1418 => x"07003304",
			1419 => x"ff071669",
			1420 => x"08001c04",
			1421 => x"ffd91669",
			1422 => x"005e1669",
			1423 => x"0300460c",
			1424 => x"0c001e04",
			1425 => x"fe951669",
			1426 => x"0c001f04",
			1427 => x"00331669",
			1428 => x"ff8a1669",
			1429 => x"0a005904",
			1430 => x"00bc1669",
			1431 => x"01000b04",
			1432 => x"fff71669",
			1433 => x"ff6c1669",
			1434 => x"05003c04",
			1435 => x"feab1707",
			1436 => x"09001d08",
			1437 => x"0000b404",
			1438 => x"017c1707",
			1439 => x"ff5e1707",
			1440 => x"05005124",
			1441 => x"0a004218",
			1442 => x"0300390c",
			1443 => x"04003908",
			1444 => x"05004304",
			1445 => x"005e1707",
			1446 => x"fec51707",
			1447 => x"00981707",
			1448 => x"08001f08",
			1449 => x"0b001804",
			1450 => x"014c1707",
			1451 => x"002c1707",
			1452 => x"fee51707",
			1453 => x"08001b04",
			1454 => x"00731707",
			1455 => x"06008a04",
			1456 => x"fe651707",
			1457 => x"00231707",
			1458 => x"08001c0c",
			1459 => x"09002104",
			1460 => x"018c1707",
			1461 => x"04004704",
			1462 => x"00a41707",
			1463 => x"ffb61707",
			1464 => x"0000c504",
			1465 => x"feb81707",
			1466 => x"0a005908",
			1467 => x"04003f04",
			1468 => x"00341707",
			1469 => x"012a1707",
			1470 => x"01000b04",
			1471 => x"fff91707",
			1472 => x"ff321707",
			1473 => x"04002e10",
			1474 => x"0500420c",
			1475 => x"04002b04",
			1476 => x"fe571779",
			1477 => x"09001f04",
			1478 => x"ffb21779",
			1479 => x"fe5c1779",
			1480 => x"fffb1779",
			1481 => x"0d001b20",
			1482 => x"0400611c",
			1483 => x"0a004510",
			1484 => x"0d00180c",
			1485 => x"07002504",
			1486 => x"02881779",
			1487 => x"0000b404",
			1488 => x"003f1779",
			1489 => x"01d31779",
			1490 => x"fee41779",
			1491 => x"08001d04",
			1492 => x"025f1779",
			1493 => x"09002504",
			1494 => x"00b91779",
			1495 => x"028d1779",
			1496 => x"fe641779",
			1497 => x"01000e08",
			1498 => x"0200d904",
			1499 => x"fe6c1779",
			1500 => x"01741779",
			1501 => x"fe5a1779",
			1502 => x"08001c30",
			1503 => x"09002018",
			1504 => x"0400340c",
			1505 => x"0000df08",
			1506 => x"04002b04",
			1507 => x"ffd61825",
			1508 => x"00981825",
			1509 => x"ffaf1825",
			1510 => x"0a004508",
			1511 => x"0f005d04",
			1512 => x"001d1825",
			1513 => x"ff4f1825",
			1514 => x"003f1825",
			1515 => x"09002108",
			1516 => x"0c001b04",
			1517 => x"00af1825",
			1518 => x"fffd1825",
			1519 => x"0200c60c",
			1520 => x"09002204",
			1521 => x"ff8f1825",
			1522 => x"01000804",
			1523 => x"00311825",
			1524 => x"fffb1825",
			1525 => x"006a1825",
			1526 => x"0000af10",
			1527 => x"0600540c",
			1528 => x"09001f08",
			1529 => x"00008804",
			1530 => x"fffa1825",
			1531 => x"002f1825",
			1532 => x"fff01825",
			1533 => x"ff4f1825",
			1534 => x"0d001508",
			1535 => x"05004404",
			1536 => x"ffec1825",
			1537 => x"007a1825",
			1538 => x"05005e08",
			1539 => x"03004604",
			1540 => x"ff821825",
			1541 => x"00001825",
			1542 => x"0a005904",
			1543 => x"003e1825",
			1544 => x"ffd71825",
			1545 => x"0d00152c",
			1546 => x"0300391c",
			1547 => x"07002508",
			1548 => x"05003c04",
			1549 => x"ff8a18d1",
			1550 => x"011818d1",
			1551 => x"0200a604",
			1552 => x"feb318d1",
			1553 => x"0000df0c",
			1554 => x"0000b504",
			1555 => x"ffb618d1",
			1556 => x"04002d04",
			1557 => x"ffea18d1",
			1558 => x"010118d1",
			1559 => x"fed918d1",
			1560 => x"04003c08",
			1561 => x"08001904",
			1562 => x"008118d1",
			1563 => x"016b18d1",
			1564 => x"05005204",
			1565 => x"ff5618d1",
			1566 => x"011718d1",
			1567 => x"0b001910",
			1568 => x"0b001608",
			1569 => x"01000b04",
			1570 => x"008018d1",
			1571 => x"ffaf18d1",
			1572 => x"01000704",
			1573 => x"ffb418d1",
			1574 => x"fea318d1",
			1575 => x"03003b08",
			1576 => x"04003504",
			1577 => x"ff5018d1",
			1578 => x"014e18d1",
			1579 => x"0a004304",
			1580 => x"fed518d1",
			1581 => x"08001f08",
			1582 => x"04004d04",
			1583 => x"00ff18d1",
			1584 => x"ffdd18d1",
			1585 => x"01000b04",
			1586 => x"002018d1",
			1587 => x"ff3818d1",
			1588 => x"0e006b38",
			1589 => x"0c001810",
			1590 => x"0d001108",
			1591 => x"01000704",
			1592 => x"ff31196d",
			1593 => x"0058196d",
			1594 => x"05003c04",
			1595 => x"ff6f196d",
			1596 => x"012a196d",
			1597 => x"00009e08",
			1598 => x"08001904",
			1599 => x"ffcb196d",
			1600 => x"feaa196d",
			1601 => x"0d001308",
			1602 => x"09002004",
			1603 => x"fee8196d",
			1604 => x"010b196d",
			1605 => x"01000708",
			1606 => x"0b001804",
			1607 => x"0132196d",
			1608 => x"0059196d",
			1609 => x"0e005108",
			1610 => x"0200a004",
			1611 => x"0146196d",
			1612 => x"ffec196d",
			1613 => x"0c001a04",
			1614 => x"ff42196d",
			1615 => x"003e196d",
			1616 => x"0c001b0c",
			1617 => x"08001908",
			1618 => x"08001804",
			1619 => x"ff9c196d",
			1620 => x"000d196d",
			1621 => x"fe9f196d",
			1622 => x"01001008",
			1623 => x"03006a04",
			1624 => x"00f8196d",
			1625 => x"ffca196d",
			1626 => x"ff1b196d",
			1627 => x"03003514",
			1628 => x"07002508",
			1629 => x"05003c04",
			1630 => x"ffd71a09",
			1631 => x"006c1a09",
			1632 => x"01000508",
			1633 => x"0000e204",
			1634 => x"00321a09",
			1635 => x"fff21a09",
			1636 => x"ff451a09",
			1637 => x"08001c18",
			1638 => x"0000f714",
			1639 => x"0900210c",
			1640 => x"09002008",
			1641 => x"09001f04",
			1642 => x"006f1a09",
			1643 => x"ffac1a09",
			1644 => x"00b71a09",
			1645 => x"0200c604",
			1646 => x"ffbd1a09",
			1647 => x"006c1a09",
			1648 => x"ffbc1a09",
			1649 => x"0f007210",
			1650 => x"0a003d04",
			1651 => x"000b1a09",
			1652 => x"0200b004",
			1653 => x"ff641a09",
			1654 => x"0200cb04",
			1655 => x"00161a09",
			1656 => x"ffe71a09",
			1657 => x"0e006504",
			1658 => x"004c1a09",
			1659 => x"0f008104",
			1660 => x"ffb31a09",
			1661 => x"00010f08",
			1662 => x"03006704",
			1663 => x"004f1a09",
			1664 => x"fff81a09",
			1665 => x"ffd91a09",
			1666 => x"0d001530",
			1667 => x"0300351c",
			1668 => x"07002508",
			1669 => x"05003c04",
			1670 => x"ffe91abd",
			1671 => x"003f1abd",
			1672 => x"01000508",
			1673 => x"09001e04",
			1674 => x"fff91abd",
			1675 => x"00301abd",
			1676 => x"0c001904",
			1677 => x"ff901abd",
			1678 => x"09002004",
			1679 => x"fffd1abd",
			1680 => x"00091abd",
			1681 => x"0900210c",
			1682 => x"08001c08",
			1683 => x"0c001904",
			1684 => x"00a21abd",
			1685 => x"000e1abd",
			1686 => x"000b1abd",
			1687 => x"0000c704",
			1688 => x"ffb41abd",
			1689 => x"00391abd",
			1690 => x"0b001910",
			1691 => x"01000704",
			1692 => x"000a1abd",
			1693 => x"0b001608",
			1694 => x"05003304",
			1695 => x"fff61abd",
			1696 => x"00151abd",
			1697 => x"ff751abd",
			1698 => x"0a003b04",
			1699 => x"ffc21abd",
			1700 => x"03003e08",
			1701 => x"04003604",
			1702 => x"fff01abd",
			1703 => x"007a1abd",
			1704 => x"0200b904",
			1705 => x"ffaa1abd",
			1706 => x"0a005908",
			1707 => x"00010a04",
			1708 => x"00451abd",
			1709 => x"fffa1abd",
			1710 => x"ffdf1abd",
			1711 => x"0e00653c",
			1712 => x"0000a218",
			1713 => x"09001d08",
			1714 => x"05003c04",
			1715 => x"ffea1b89",
			1716 => x"004c1b89",
			1717 => x"0c001808",
			1718 => x"0e004904",
			1719 => x"00111b89",
			1720 => x"00001b89",
			1721 => x"08001904",
			1722 => x"00031b89",
			1723 => x"ff8f1b89",
			1724 => x"0500450c",
			1725 => x"06006908",
			1726 => x"03003104",
			1727 => x"00061b89",
			1728 => x"ffc61b89",
			1729 => x"00111b89",
			1730 => x"0d00170c",
			1731 => x"07002c08",
			1732 => x"08001804",
			1733 => x"00081b89",
			1734 => x"00721b89",
			1735 => x"fff11b89",
			1736 => x"0200b904",
			1737 => x"ffd21b89",
			1738 => x"07003304",
			1739 => x"001b1b89",
			1740 => x"fff61b89",
			1741 => x"0000d60c",
			1742 => x"05004d08",
			1743 => x"07002e04",
			1744 => x"00001b89",
			1745 => x"00041b89",
			1746 => x"ff971b89",
			1747 => x"0000fa10",
			1748 => x"03003508",
			1749 => x"0200d804",
			1750 => x"00171b89",
			1751 => x"ffde1b89",
			1752 => x"03005c04",
			1753 => x"00631b89",
			1754 => x"fff41b89",
			1755 => x"05005008",
			1756 => x"03003d04",
			1757 => x"ffbb1b89",
			1758 => x"00021b89",
			1759 => x"03005304",
			1760 => x"00131b89",
			1761 => x"ffef1b89",
			1762 => x"04002e10",
			1763 => x"0500420c",
			1764 => x"04002b04",
			1765 => x"fe541c0d",
			1766 => x"0b001704",
			1767 => x"ff871c0d",
			1768 => x"fe591c0d",
			1769 => x"fff41c0d",
			1770 => x"0d001b28",
			1771 => x"04006124",
			1772 => x"0a004718",
			1773 => x"0d00150c",
			1774 => x"0e006508",
			1775 => x"0b001804",
			1776 => x"02611c0d",
			1777 => x"01251c0d",
			1778 => x"010d1c0d",
			1779 => x"0000d008",
			1780 => x"03003d04",
			1781 => x"00481c0d",
			1782 => x"fde41c0d",
			1783 => x"01b71c0d",
			1784 => x"0c001e08",
			1785 => x"0a004804",
			1786 => x"01f01c0d",
			1787 => x"027d1c0d",
			1788 => x"02d61c0d",
			1789 => x"fe5f1c0d",
			1790 => x"01000e08",
			1791 => x"0f007704",
			1792 => x"fe671c0d",
			1793 => x"019f1c0d",
			1794 => x"fe571c0d",
			1795 => x"05004b2c",
			1796 => x"07002508",
			1797 => x"05003e04",
			1798 => x"ffdd1cb1",
			1799 => x"00641cb1",
			1800 => x"0000ab0c",
			1801 => x"09001d04",
			1802 => x"00251cb1",
			1803 => x"01000504",
			1804 => x"001c1cb1",
			1805 => x"ff3d1cb1",
			1806 => x"0200d20c",
			1807 => x"0f006404",
			1808 => x"ffde1cb1",
			1809 => x"04002d04",
			1810 => x"fff01cb1",
			1811 => x"00871cb1",
			1812 => x"01000504",
			1813 => x"000e1cb1",
			1814 => x"0a004204",
			1815 => x"ff851cb1",
			1816 => x"000f1cb1",
			1817 => x"08001b0c",
			1818 => x"03004104",
			1819 => x"009d1cb1",
			1820 => x"03004504",
			1821 => x"ffd51cb1",
			1822 => x"00211cb1",
			1823 => x"06005d04",
			1824 => x"003c1cb1",
			1825 => x"0000b504",
			1826 => x"ff6f1cb1",
			1827 => x"0e006508",
			1828 => x"04004d04",
			1829 => x"00701cb1",
			1830 => x"ffdd1cb1",
			1831 => x"0200cd04",
			1832 => x"ff9e1cb1",
			1833 => x"0d001b04",
			1834 => x"00431cb1",
			1835 => x"ffd41cb1",
			1836 => x"05003e08",
			1837 => x"05003c04",
			1838 => x"fe5b1d1d",
			1839 => x"ff481d1d",
			1840 => x"0d001b24",
			1841 => x"00011020",
			1842 => x"09001d04",
			1843 => x"02831d1d",
			1844 => x"0000b410",
			1845 => x"0e005508",
			1846 => x"05004b04",
			1847 => x"ffa61d1d",
			1848 => x"029c1d1d",
			1849 => x"0c001a04",
			1850 => x"fe031d1d",
			1851 => x"003e1d1d",
			1852 => x"03005c08",
			1853 => x"0a004704",
			1854 => x"01681d1d",
			1855 => x"01fc1d1d",
			1856 => x"fe7e1d1d",
			1857 => x"fee41d1d",
			1858 => x"01000d08",
			1859 => x"03007c04",
			1860 => x"01771d1d",
			1861 => x"fe761d1d",
			1862 => x"fe5c1d1d",
			1863 => x"08001d2c",
			1864 => x"0a004524",
			1865 => x"0a00421c",
			1866 => x"05004914",
			1867 => x"0000df10",
			1868 => x"0f006608",
			1869 => x"09001d04",
			1870 => x"008b1db9",
			1871 => x"ff3c1db9",
			1872 => x"01000904",
			1873 => x"00bd1db9",
			1874 => x"ffaf1db9",
			1875 => x"ff631db9",
			1876 => x"0e005c04",
			1877 => x"00a71db9",
			1878 => x"00041db9",
			1879 => x"08001b04",
			1880 => x"001a1db9",
			1881 => x"ff431db9",
			1882 => x"09002504",
			1883 => x"00bf1db9",
			1884 => x"fffb1db9",
			1885 => x"09001f08",
			1886 => x"0a003604",
			1887 => x"ffe81db9",
			1888 => x"004e1db9",
			1889 => x"05005e14",
			1890 => x"07002f04",
			1891 => x"ff3c1db9",
			1892 => x"03003a04",
			1893 => x"ffd81db9",
			1894 => x"03004908",
			1895 => x"07003704",
			1896 => x"001b1db9",
			1897 => x"fffa1db9",
			1898 => x"fff41db9",
			1899 => x"0a005904",
			1900 => x"00441db9",
			1901 => x"ffc51db9",
			1902 => x"0e006530",
			1903 => x"0000b91c",
			1904 => x"06006418",
			1905 => x"08001d10",
			1906 => x"0000ad0c",
			1907 => x"0e005508",
			1908 => x"08001b04",
			1909 => x"ffad1e7d",
			1910 => x"00ad1e7d",
			1911 => x"ff211e7d",
			1912 => x"00c11e7d",
			1913 => x"09001d04",
			1914 => x"000e1e7d",
			1915 => x"fed91e7d",
			1916 => x"fedf1e7d",
			1917 => x"0f006604",
			1918 => x"ff641e7d",
			1919 => x"0200d00c",
			1920 => x"0d001604",
			1921 => x"01401e7d",
			1922 => x"07003504",
			1923 => x"00531e7d",
			1924 => x"ffc81e7d",
			1925 => x"ff9d1e7d",
			1926 => x"0a004824",
			1927 => x"08001b14",
			1928 => x"0000e108",
			1929 => x"0000d004",
			1930 => x"ff921e7d",
			1931 => x"010f1e7d",
			1932 => x"07002b04",
			1933 => x"fee51e7d",
			1934 => x"01000704",
			1935 => x"00781e7d",
			1936 => x"ff841e7d",
			1937 => x"0c001b08",
			1938 => x"0b001904",
			1939 => x"fe9b1e7d",
			1940 => x"ffcc1e7d",
			1941 => x"00010c04",
			1942 => x"005c1e7d",
			1943 => x"ff641e7d",
			1944 => x"0a005908",
			1945 => x"00010304",
			1946 => x"00cd1e7d",
			1947 => x"00121e7d",
			1948 => x"0d001b04",
			1949 => x"001d1e7d",
			1950 => x"ff791e7d",
			1951 => x"0d001428",
			1952 => x"05004920",
			1953 => x"0700250c",
			1954 => x"0d001004",
			1955 => x"ffea1f41",
			1956 => x"04002b04",
			1957 => x"fff41f41",
			1958 => x"00411f41",
			1959 => x"06005e04",
			1960 => x"ff9b1f41",
			1961 => x"0b001608",
			1962 => x"0d001304",
			1963 => x"ffd81f41",
			1964 => x"00031f41",
			1965 => x"06008104",
			1966 => x"003f1f41",
			1967 => x"fff61f41",
			1968 => x"09002104",
			1969 => x"007a1f41",
			1970 => x"00021f41",
			1971 => x"0000ca18",
			1972 => x"07002608",
			1973 => x"00008f04",
			1974 => x"fff31f41",
			1975 => x"00361f41",
			1976 => x"03003308",
			1977 => x"09001f04",
			1978 => x"ffdb1f41",
			1979 => x"00301f41",
			1980 => x"0a004704",
			1981 => x"ff5d1f41",
			1982 => x"000d1f41",
			1983 => x"0e006908",
			1984 => x"0f007304",
			1985 => x"ffe81f41",
			1986 => x"00651f41",
			1987 => x"0c001b0c",
			1988 => x"0a003908",
			1989 => x"0a003604",
			1990 => x"fff61f41",
			1991 => x"000a1f41",
			1992 => x"ffb41f41",
			1993 => x"0201020c",
			1994 => x"03005c08",
			1995 => x"0a003d04",
			1996 => x"fffe1f41",
			1997 => x"00471f41",
			1998 => x"fff11f41",
			1999 => x"ffe71f41",
			2000 => x"0000ed3c",
			2001 => x"00009e0c",
			2002 => x"0c001808",
			2003 => x"05003c04",
			2004 => x"ffbd1fcd",
			2005 => x"00ae1fcd",
			2006 => x"fef41fcd",
			2007 => x"04004724",
			2008 => x"0d001310",
			2009 => x"0900200c",
			2010 => x"05004e08",
			2011 => x"05004404",
			2012 => x"00361fcd",
			2013 => x"ff181fcd",
			2014 => x"00561fcd",
			2015 => x"00aa1fcd",
			2016 => x"01000704",
			2017 => x"00f51fcd",
			2018 => x"09002108",
			2019 => x"01000804",
			2020 => x"ff831fcd",
			2021 => x"00b21fcd",
			2022 => x"0200b904",
			2023 => x"ff1f1fcd",
			2024 => x"00611fcd",
			2025 => x"07003004",
			2026 => x"ff711fcd",
			2027 => x"03005c04",
			2028 => x"00811fcd",
			2029 => x"ffd11fcd",
			2030 => x"05005004",
			2031 => x"ff281fcd",
			2032 => x"0a004f04",
			2033 => x"004e1fcd",
			2034 => x"ffcb1fcd",
			2035 => x"0d00153c",
			2036 => x"0e006524",
			2037 => x"0000b418",
			2038 => x"0e005714",
			2039 => x"0500460c",
			2040 => x"07002508",
			2041 => x"05003c04",
			2042 => x"ffed2099",
			2043 => x"00302099",
			2044 => x"ffbc2099",
			2045 => x"09001f04",
			2046 => x"005f2099",
			2047 => x"00092099",
			2048 => x"ffb32099",
			2049 => x"07002708",
			2050 => x"09001c04",
			2051 => x"fff22099",
			2052 => x"00012099",
			2053 => x"00792099",
			2054 => x"07002b0c",
			2055 => x"03003108",
			2056 => x"03002c04",
			2057 => x"fffb2099",
			2058 => x"00112099",
			2059 => x"ffa62099",
			2060 => x"0000cd04",
			2061 => x"ffd12099",
			2062 => x"09001e04",
			2063 => x"fff02099",
			2064 => x"00502099",
			2065 => x"01000708",
			2066 => x"08001c04",
			2067 => x"00422099",
			2068 => x"ffea2099",
			2069 => x"0a004714",
			2070 => x"0b001608",
			2071 => x"06006f04",
			2072 => x"00152099",
			2073 => x"fff72099",
			2074 => x"07003004",
			2075 => x"ff5f2099",
			2076 => x"0f009f04",
			2077 => x"00162099",
			2078 => x"ffeb2099",
			2079 => x"0a00590c",
			2080 => x"0f007204",
			2081 => x"fffb2099",
			2082 => x"0f00a204",
			2083 => x"003e2099",
			2084 => x"fffd2099",
			2085 => x"ffdd2099",
			2086 => x"0100071c",
			2087 => x"05004914",
			2088 => x"0f006604",
			2089 => x"ffac2145",
			2090 => x"0000e108",
			2091 => x"0a002c04",
			2092 => x"fffb2145",
			2093 => x"00582145",
			2094 => x"07002e04",
			2095 => x"ffc22145",
			2096 => x"000a2145",
			2097 => x"04004304",
			2098 => x"00a62145",
			2099 => x"ffd42145",
			2100 => x"07002508",
			2101 => x"05003c04",
			2102 => x"ffed2145",
			2103 => x"005c2145",
			2104 => x"0a004724",
			2105 => x"0a003b0c",
			2106 => x"0e004d08",
			2107 => x"06004d04",
			2108 => x"ffe92145",
			2109 => x"00212145",
			2110 => x"ff762145",
			2111 => x"0900210c",
			2112 => x"01000804",
			2113 => x"ffb62145",
			2114 => x"04003804",
			2115 => x"fff72145",
			2116 => x"006f2145",
			2117 => x"0f007f04",
			2118 => x"ff792145",
			2119 => x"04003404",
			2120 => x"fff62145",
			2121 => x"00322145",
			2122 => x"0a005908",
			2123 => x"08002304",
			2124 => x"005a2145",
			2125 => x"fff62145",
			2126 => x"01000b04",
			2127 => x"00002145",
			2128 => x"ffda2145",
			2129 => x"0d001540",
			2130 => x"05004928",
			2131 => x"07002514",
			2132 => x"05003e10",
			2133 => x"01000704",
			2134 => x"ffad2219",
			2135 => x"01000808",
			2136 => x"08001904",
			2137 => x"002c2219",
			2138 => x"fffa2219",
			2139 => x"ffd92219",
			2140 => x"00be2219",
			2141 => x"06005e04",
			2142 => x"feda2219",
			2143 => x"0000df0c",
			2144 => x"01000908",
			2145 => x"03002f04",
			2146 => x"fff32219",
			2147 => x"01062219",
			2148 => x"ff932219",
			2149 => x"ff192219",
			2150 => x"04003c08",
			2151 => x"0000b504",
			2152 => x"00692219",
			2153 => x"01282219",
			2154 => x"05005308",
			2155 => x"04003e04",
			2156 => x"ffd22219",
			2157 => x"ff422219",
			2158 => x"09002104",
			2159 => x"00d62219",
			2160 => x"000d2219",
			2161 => x"0200b90c",
			2162 => x"01000704",
			2163 => x"004a2219",
			2164 => x"0c001604",
			2165 => x"fff82219",
			2166 => x"feaa2219",
			2167 => x"0b00190c",
			2168 => x"0b001708",
			2169 => x"0b001604",
			2170 => x"ffd12219",
			2171 => x"00072219",
			2172 => x"ff382219",
			2173 => x"01000d0c",
			2174 => x"03006108",
			2175 => x"04003404",
			2176 => x"ffec2219",
			2177 => x"01002219",
			2178 => x"ffdf2219",
			2179 => x"08002004",
			2180 => x"002f2219",
			2181 => x"ff562219",
			2182 => x"0a003614",
			2183 => x"07002510",
			2184 => x"07002004",
			2185 => x"ffd522c5",
			2186 => x"0c001708",
			2187 => x"0c001504",
			2188 => x"fffa22c5",
			2189 => x"004922c5",
			2190 => x"fff822c5",
			2191 => x"ff3822c5",
			2192 => x"08001d28",
			2193 => x"0d001620",
			2194 => x"05004910",
			2195 => x"0d001308",
			2196 => x"0a003904",
			2197 => x"002922c5",
			2198 => x"ff3422c5",
			2199 => x"0000ae04",
			2200 => x"ffee22c5",
			2201 => x"00a922c5",
			2202 => x"0e005604",
			2203 => x"00d622c5",
			2204 => x"0000b504",
			2205 => x"ff7422c5",
			2206 => x"09002004",
			2207 => x"ffeb22c5",
			2208 => x"00d222c5",
			2209 => x"06007604",
			2210 => x"ff8322c5",
			2211 => x"000d22c5",
			2212 => x"0f007208",
			2213 => x"06005804",
			2214 => x"002722c5",
			2215 => x"ff2922c5",
			2216 => x"0e006704",
			2217 => x"007722c5",
			2218 => x"0b001a04",
			2219 => x"ff7122c5",
			2220 => x"0d001c08",
			2221 => x"03006104",
			2222 => x"006422c5",
			2223 => x"ffea22c5",
			2224 => x"ffc722c5",
			2225 => x"0000ed44",
			2226 => x"09001e0c",
			2227 => x"05003c04",
			2228 => x"ffa02369",
			2229 => x"0d001204",
			2230 => x"001a2369",
			2231 => x"00f62369",
			2232 => x"0000b41c",
			2233 => x"0e005514",
			2234 => x"05004b10",
			2235 => x"07002b08",
			2236 => x"01000504",
			2237 => x"00492369",
			2238 => x"fef22369",
			2239 => x"01000c04",
			2240 => x"00562369",
			2241 => x"fffb2369",
			2242 => x"00bf2369",
			2243 => x"05004704",
			2244 => x"00412369",
			2245 => x"fedf2369",
			2246 => x"0e005f0c",
			2247 => x"0d001704",
			2248 => x"01062369",
			2249 => x"07002c04",
			2250 => x"ffab2369",
			2251 => x"002e2369",
			2252 => x"0000c704",
			2253 => x"ff2c2369",
			2254 => x"07002b04",
			2255 => x"ffba2369",
			2256 => x"0d001804",
			2257 => x"010b2369",
			2258 => x"ffeb2369",
			2259 => x"05005008",
			2260 => x"03003d04",
			2261 => x"ff282369",
			2262 => x"00022369",
			2263 => x"03005304",
			2264 => x"00342369",
			2265 => x"ffc82369",
			2266 => x"0500524c",
			2267 => x"0e005b24",
			2268 => x"0600621c",
			2269 => x"09001e10",
			2270 => x"00008104",
			2271 => x"ffd0242d",
			2272 => x"01000504",
			2273 => x"fff5242d",
			2274 => x"05003c04",
			2275 => x"fff5242d",
			2276 => x"0083242d",
			2277 => x"05004b08",
			2278 => x"06005d04",
			2279 => x"ff56242d",
			2280 => x"0014242d",
			2281 => x"0010242d",
			2282 => x"0000bc04",
			2283 => x"0072242d",
			2284 => x"0000242d",
			2285 => x"0100050c",
			2286 => x"0000d104",
			2287 => x"ffe9242d",
			2288 => x"0a003604",
			2289 => x"fff6242d",
			2290 => x"004c242d",
			2291 => x"0d00140c",
			2292 => x"03003508",
			2293 => x"01000a04",
			2294 => x"ffa8242d",
			2295 => x"0001242d",
			2296 => x"003f242d",
			2297 => x"0a00470c",
			2298 => x"0b001608",
			2299 => x"0b001504",
			2300 => x"fff4242d",
			2301 => x"0008242d",
			2302 => x"ff61242d",
			2303 => x"0002242d",
			2304 => x"08001c08",
			2305 => x"06007504",
			2306 => x"0094242d",
			2307 => x"fffd242d",
			2308 => x"07002f04",
			2309 => x"ffb3242d",
			2310 => x"0a005904",
			2311 => x"004e242d",
			2312 => x"01000b04",
			2313 => x"0001242d",
			2314 => x"ffd7242d",
			2315 => x"05003c04",
			2316 => x"fe7b24a9",
			2317 => x"09001e0c",
			2318 => x"05004708",
			2319 => x"07002504",
			2320 => x"017b24a9",
			2321 => x"ff1b24a9",
			2322 => x"01bf24a9",
			2323 => x"0000b410",
			2324 => x"0a003b04",
			2325 => x"fe6524a9",
			2326 => x"0e005504",
			2327 => x"008124a9",
			2328 => x"06006304",
			2329 => x"fe7624a9",
			2330 => x"001224a9",
			2331 => x"0b001708",
			2332 => x"04003b04",
			2333 => x"016f24a9",
			2334 => x"00c024a9",
			2335 => x"09002008",
			2336 => x"0000cc04",
			2337 => x"004c24a9",
			2338 => x"fe9024a9",
			2339 => x"0d001508",
			2340 => x"07002d04",
			2341 => x"019124a9",
			2342 => x"006a24a9",
			2343 => x"0f008104",
			2344 => x"ff8824a9",
			2345 => x"009e24a9",
			2346 => x"05003c04",
			2347 => x"fe692515",
			2348 => x"0201012c",
			2349 => x"09001e08",
			2350 => x"01000804",
			2351 => x"00612515",
			2352 => x"01f52515",
			2353 => x"0000c714",
			2354 => x"0e006210",
			2355 => x"05004b08",
			2356 => x"06005d04",
			2357 => x"fe3d2515",
			2358 => x"00652515",
			2359 => x"09002104",
			2360 => x"01752515",
			2361 => x"ff832515",
			2362 => x"fdfc2515",
			2363 => x"07002b04",
			2364 => x"ffca2515",
			2365 => x"0d001604",
			2366 => x"01c92515",
			2367 => x"0f007f04",
			2368 => x"ff772515",
			2369 => x"011c2515",
			2370 => x"05005204",
			2371 => x"fe662515",
			2372 => x"004e2515",
			2373 => x"0500410c",
			2374 => x"05003c04",
			2375 => x"fe4f25a1",
			2376 => x"0d001404",
			2377 => x"01c325a1",
			2378 => x"fe4a25a1",
			2379 => x"0d001b30",
			2380 => x"03005c2c",
			2381 => x"0000b414",
			2382 => x"0c001808",
			2383 => x"0f005b04",
			2384 => x"03c525a1",
			2385 => x"027625a1",
			2386 => x"0d001404",
			2387 => x"019c25a1",
			2388 => x"0b001904",
			2389 => x"fe4125a1",
			2390 => x"001325a1",
			2391 => x"0d00150c",
			2392 => x"0e006508",
			2393 => x"0b001804",
			2394 => x"037b25a1",
			2395 => x"02e525a1",
			2396 => x"027c25a1",
			2397 => x"0b001904",
			2398 => x"ff7e25a1",
			2399 => x"0200c704",
			2400 => x"022025a1",
			2401 => x"035125a1",
			2402 => x"fe6025a1",
			2403 => x"0b001f08",
			2404 => x"0600ac04",
			2405 => x"00a125a1",
			2406 => x"fe5c25a1",
			2407 => x"fe5125a1",
			2408 => x"05003c04",
			2409 => x"fe7d262d",
			2410 => x"0b001714",
			2411 => x"0500490c",
			2412 => x"03003304",
			2413 => x"0129262d",
			2414 => x"0d001304",
			2415 => x"feea262d",
			2416 => x"004f262d",
			2417 => x"05004f04",
			2418 => x"0162262d",
			2419 => x"0043262d",
			2420 => x"05004f14",
			2421 => x"01000704",
			2422 => x"ffe5262d",
			2423 => x"0000b504",
			2424 => x"fe65262d",
			2425 => x"0e005b04",
			2426 => x"00f2262d",
			2427 => x"05004504",
			2428 => x"ffc9262d",
			2429 => x"fe97262d",
			2430 => x"09002108",
			2431 => x"0b001804",
			2432 => x"0182262d",
			2433 => x"00a9262d",
			2434 => x"0f00810c",
			2435 => x"0e006808",
			2436 => x"0200b904",
			2437 => x"fe9b262d",
			2438 => x"00b9262d",
			2439 => x"fe55262d",
			2440 => x"01001004",
			2441 => x"015d262d",
			2442 => x"ff09262d",
			2443 => x"0d001530",
			2444 => x"03003920",
			2445 => x"07002508",
			2446 => x"05003e04",
			2447 => x"ffda2701",
			2448 => x"007a2701",
			2449 => x"0000b50c",
			2450 => x"09001d04",
			2451 => x"00382701",
			2452 => x"0c001b04",
			2453 => x"ff412701",
			2454 => x"001d2701",
			2455 => x"0000df08",
			2456 => x"04002e04",
			2457 => x"fff72701",
			2458 => x"00822701",
			2459 => x"ffa12701",
			2460 => x"04003c04",
			2461 => x"00b12701",
			2462 => x"08001b08",
			2463 => x"09002004",
			2464 => x"00042701",
			2465 => x"00862701",
			2466 => x"ffa92701",
			2467 => x"0b001914",
			2468 => x"0b001608",
			2469 => x"06006f04",
			2470 => x"00192701",
			2471 => x"fff12701",
			2472 => x"04002f08",
			2473 => x"0a003604",
			2474 => x"fff72701",
			2475 => x"00162701",
			2476 => x"ff3a2701",
			2477 => x"0a003b04",
			2478 => x"ff922701",
			2479 => x"04004614",
			2480 => x"01000e08",
			2481 => x"08001d04",
			2482 => x"00b72701",
			2483 => x"000a2701",
			2484 => x"06007004",
			2485 => x"ffd92701",
			2486 => x"0600a104",
			2487 => x"000d2701",
			2488 => x"fff32701",
			2489 => x"0f007204",
			2490 => x"ffa82701",
			2491 => x"0e006804",
			2492 => x"003e2701",
			2493 => x"0e007104",
			2494 => x"ffc62701",
			2495 => x"001e2701",
			2496 => x"04002b04",
			2497 => x"fe842785",
			2498 => x"0e005a18",
			2499 => x"08001d14",
			2500 => x"0f00630c",
			2501 => x"09001d04",
			2502 => x"01a92785",
			2503 => x"06005704",
			2504 => x"ff112785",
			2505 => x"00282785",
			2506 => x"03003d04",
			2507 => x"019c2785",
			2508 => x"ffc72785",
			2509 => x"ff0f2785",
			2510 => x"0000b908",
			2511 => x"0c001a04",
			2512 => x"fe852785",
			2513 => x"ff7c2785",
			2514 => x"0e006510",
			2515 => x"0d001504",
			2516 => x"01992785",
			2517 => x"06006804",
			2518 => x"fef32785",
			2519 => x"06006b04",
			2520 => x"01162785",
			2521 => x"fff82785",
			2522 => x"0000d604",
			2523 => x"ff122785",
			2524 => x"07002c04",
			2525 => x"ff382785",
			2526 => x"02010504",
			2527 => x"01482785",
			2528 => x"fee12785",
			2529 => x"0100093c",
			2530 => x"08001d2c",
			2531 => x"0000ed24",
			2532 => x"0300391c",
			2533 => x"0700280c",
			2534 => x"07002508",
			2535 => x"05003c04",
			2536 => x"fff02861",
			2537 => x"00402861",
			2538 => x"ff902861",
			2539 => x"06007808",
			2540 => x"0000ae04",
			2541 => x"fffe2861",
			2542 => x"007b2861",
			2543 => x"07002d04",
			2544 => x"ffcd2861",
			2545 => x"00152861",
			2546 => x"0c001b04",
			2547 => x"00bb2861",
			2548 => x"fff82861",
			2549 => x"07003204",
			2550 => x"ffd72861",
			2551 => x"ffff2861",
			2552 => x"07002704",
			2553 => x"00162861",
			2554 => x"0a003d08",
			2555 => x"09002204",
			2556 => x"000c2861",
			2557 => x"fffc2861",
			2558 => x"ffaf2861",
			2559 => x"04004320",
			2560 => x"0200be10",
			2561 => x"09001e0c",
			2562 => x"00008804",
			2563 => x"fff52861",
			2564 => x"06005604",
			2565 => x"003a2861",
			2566 => x"fffe2861",
			2567 => x"ff662861",
			2568 => x"0201010c",
			2569 => x"0a003b04",
			2570 => x"ffed2861",
			2571 => x"06006a04",
			2572 => x"fffe2861",
			2573 => x"00522861",
			2574 => x"ffd62861",
			2575 => x"04004b08",
			2576 => x"07003204",
			2577 => x"00542861",
			2578 => x"fffb2861",
			2579 => x"0e007104",
			2580 => x"ffbf2861",
			2581 => x"07003e04",
			2582 => x"001b2861",
			2583 => x"fffa2861",
			2584 => x"08001d4c",
			2585 => x"0100092c",
			2586 => x"05005224",
			2587 => x"0a004220",
			2588 => x"08001910",
			2589 => x"0000e008",
			2590 => x"07002804",
			2591 => x"ff97292d",
			2592 => x"00be292d",
			2593 => x"07002b04",
			2594 => x"ff3b292d",
			2595 => x"fff6292d",
			2596 => x"0000ae08",
			2597 => x"07002704",
			2598 => x"0079292d",
			2599 => x"ff52292d",
			2600 => x"05003c04",
			2601 => x"ffd9292d",
			2602 => x"0111292d",
			2603 => x"ff51292d",
			2604 => x"05005904",
			2605 => x"011b292d",
			2606 => x"002b292d",
			2607 => x"0700270c",
			2608 => x"0f005304",
			2609 => x"ffcc292d",
			2610 => x"05003704",
			2611 => x"fff8292d",
			2612 => x"00d5292d",
			2613 => x"0c001b0c",
			2614 => x"01000e08",
			2615 => x"07003004",
			2616 => x"fefa292d",
			2617 => x"0005292d",
			2618 => x"0024292d",
			2619 => x"0f006904",
			2620 => x"ffb0292d",
			2621 => x"0081292d",
			2622 => x"09001f08",
			2623 => x"0a003604",
			2624 => x"ffce292d",
			2625 => x"008a292d",
			2626 => x"05005e08",
			2627 => x"03004604",
			2628 => x"fef2292d",
			2629 => x"fff6292d",
			2630 => x"0f007204",
			2631 => x"ffa5292d",
			2632 => x"0a005904",
			2633 => x"00a3292d",
			2634 => x"ffc0292d",
			2635 => x"05003c04",
			2636 => x"fe612999",
			2637 => x"0800232c",
			2638 => x"03005c28",
			2639 => x"05004f14",
			2640 => x"07002508",
			2641 => x"03003304",
			2642 => x"022f2999",
			2643 => x"01972999",
			2644 => x"00009e04",
			2645 => x"fe902999",
			2646 => x"0000dd04",
			2647 => x"00c62999",
			2648 => x"fee12999",
			2649 => x"09002108",
			2650 => x"0000ba04",
			2651 => x"02522999",
			2652 => x"01a52999",
			2653 => x"0000c704",
			2654 => x"ff9e2999",
			2655 => x"0c001b04",
			2656 => x"00ef2999",
			2657 => x"01dd2999",
			2658 => x"fe732999",
			2659 => x"01001004",
			2660 => x"00002999",
			2661 => x"fe5f2999",
			2662 => x"05003e04",
			2663 => x"fe652a0d",
			2664 => x"02010130",
			2665 => x"09001e08",
			2666 => x"01000804",
			2667 => x"00a62a0d",
			2668 => x"021c2a0d",
			2669 => x"01000910",
			2670 => x"0a00450c",
			2671 => x"0e006508",
			2672 => x"0000ae04",
			2673 => x"ffed2a0d",
			2674 => x"01842a0d",
			2675 => x"ff852a0d",
			2676 => x"019e2a0d",
			2677 => x"0000c70c",
			2678 => x"04004308",
			2679 => x"0e005a04",
			2680 => x"ff502a0d",
			2681 => x"fe152a0d",
			2682 => x"00bd2a0d",
			2683 => x"0a005b08",
			2684 => x"07002f04",
			2685 => x"00692a0d",
			2686 => x"018b2a0d",
			2687 => x"fe932a0d",
			2688 => x"05005204",
			2689 => x"fe602a0d",
			2690 => x"00122a0d",
			2691 => x"0000ed58",
			2692 => x"01000928",
			2693 => x"08001d20",
			2694 => x"0600570c",
			2695 => x"0c001808",
			2696 => x"05003c04",
			2697 => x"ffee2ad9",
			2698 => x"005a2ad9",
			2699 => x"ff8f2ad9",
			2700 => x"09001e0c",
			2701 => x"06005f04",
			2702 => x"ffe42ad9",
			2703 => x"07002904",
			2704 => x"00102ad9",
			2705 => x"fffc2ad9",
			2706 => x"04004304",
			2707 => x"00bd2ad9",
			2708 => x"000d2ad9",
			2709 => x"01000804",
			2710 => x"ffbb2ad9",
			2711 => x"00222ad9",
			2712 => x"0200b918",
			2713 => x"0e005a14",
			2714 => x"08001c08",
			2715 => x"05003f04",
			2716 => x"fff02ad9",
			2717 => x"007d2ad9",
			2718 => x"0200a808",
			2719 => x"09001e04",
			2720 => x"00082ad9",
			2721 => x"ffb02ad9",
			2722 => x"00132ad9",
			2723 => x"ff532ad9",
			2724 => x"04004c10",
			2725 => x"08001f08",
			2726 => x"04003404",
			2727 => x"fff92ad9",
			2728 => x"008d2ad9",
			2729 => x"07003004",
			2730 => x"ffe12ad9",
			2731 => x"000b2ad9",
			2732 => x"0e006d04",
			2733 => x"ffcc2ad9",
			2734 => x"001c2ad9",
			2735 => x"05005008",
			2736 => x"03003d04",
			2737 => x"ff802ad9",
			2738 => x"00042ad9",
			2739 => x"03005304",
			2740 => x"002d2ad9",
			2741 => x"ffdf2ad9",
			2742 => x"05003c04",
			2743 => x"fe602b45",
			2744 => x"0100102c",
			2745 => x"03005c28",
			2746 => x"0a00481c",
			2747 => x"0d00150c",
			2748 => x"0000f208",
			2749 => x"09001d04",
			2750 => x"024c2b45",
			2751 => x"01012b45",
			2752 => x"ff302b45",
			2753 => x"0b001908",
			2754 => x"05004b04",
			2755 => x"ff9e2b45",
			2756 => x"fe412b45",
			2757 => x"0000d204",
			2758 => x"ffeb2b45",
			2759 => x"01a92b45",
			2760 => x"0000ca04",
			2761 => x"013a2b45",
			2762 => x"07003704",
			2763 => x"01ca2b45",
			2764 => x"02272b45",
			2765 => x"fe712b45",
			2766 => x"07003104",
			2767 => x"00232b45",
			2768 => x"fe5c2b45",
			2769 => x"05003c04",
			2770 => x"fe742bc1",
			2771 => x"09001d08",
			2772 => x"0000a404",
			2773 => x"01cb2bc1",
			2774 => x"ff5f2bc1",
			2775 => x"05004914",
			2776 => x"0f006604",
			2777 => x"fe712bc1",
			2778 => x"0000df04",
			2779 => x"00be2bc1",
			2780 => x"05004208",
			2781 => x"05004004",
			2782 => x"ff352bc1",
			2783 => x"00902bc1",
			2784 => x"fdfd2bc1",
			2785 => x"0e005a0c",
			2786 => x"09002108",
			2787 => x"01000804",
			2788 => x"00ab2bc1",
			2789 => x"01bb2bc1",
			2790 => x"00382bc1",
			2791 => x"0000b904",
			2792 => x"fea62bc1",
			2793 => x"0e006508",
			2794 => x"0200b904",
			2795 => x"00512bc1",
			2796 => x"018a2bc1",
			2797 => x"0200cc04",
			2798 => x"fee72bc1",
			2799 => x"00cd2bc1",
			2800 => x"05003c04",
			2801 => x"fe762c45",
			2802 => x"09001d08",
			2803 => x"0000a404",
			2804 => x"01c32c45",
			2805 => x"ff732c45",
			2806 => x"05004914",
			2807 => x"0f006608",
			2808 => x"01000904",
			2809 => x"fe5a2c45",
			2810 => x"feff2c45",
			2811 => x"05004708",
			2812 => x"0000f204",
			2813 => x"01652c45",
			2814 => x"feaa2c45",
			2815 => x"fed72c45",
			2816 => x"0e005c10",
			2817 => x"08001d0c",
			2818 => x"0d001408",
			2819 => x"0e005904",
			2820 => x"01cd2c45",
			2821 => x"00cc2c45",
			2822 => x"00d82c45",
			2823 => x"ff732c45",
			2824 => x"0000c004",
			2825 => x"fe6a2c45",
			2826 => x"0e006508",
			2827 => x"09002704",
			2828 => x"018a2c45",
			2829 => x"ff362c45",
			2830 => x"0200cc04",
			2831 => x"ff072c45",
			2832 => x"00bc2c45",
			2833 => x"0b001714",
			2834 => x"05003c04",
			2835 => x"ffbd2cf9",
			2836 => x"04003d0c",
			2837 => x"05004908",
			2838 => x"05004504",
			2839 => x"00522cf9",
			2840 => x"ffc32cf9",
			2841 => x"00972cf9",
			2842 => x"fff92cf9",
			2843 => x"05004f24",
			2844 => x"09001d04",
			2845 => x"00222cf9",
			2846 => x"0000ae08",
			2847 => x"01000504",
			2848 => x"001a2cf9",
			2849 => x"ff592cf9",
			2850 => x"06006508",
			2851 => x"0200b704",
			2852 => x"006e2cf9",
			2853 => x"ffe52cf9",
			2854 => x"01000c08",
			2855 => x"07002c04",
			2856 => x"ff9a2cf9",
			2857 => x"000c2cf9",
			2858 => x"01001004",
			2859 => x"001b2cf9",
			2860 => x"ffe42cf9",
			2861 => x"09002104",
			2862 => x"00592cf9",
			2863 => x"0000c708",
			2864 => x"0a004504",
			2865 => x"ff942cf9",
			2866 => x"00092cf9",
			2867 => x"01000b0c",
			2868 => x"03006108",
			2869 => x"0e006c04",
			2870 => x"00572cf9",
			2871 => x"00062cf9",
			2872 => x"fff82cf9",
			2873 => x"0f008104",
			2874 => x"ffd52cf9",
			2875 => x"08002304",
			2876 => x"00212cf9",
			2877 => x"ffe82cf9",
			2878 => x"04002b04",
			2879 => x"fe612d5d",
			2880 => x"0201052c",
			2881 => x"0a005c28",
			2882 => x"0a004518",
			2883 => x"0d001710",
			2884 => x"07002508",
			2885 => x"0d001204",
			2886 => x"016b2d5d",
			2887 => x"01f42d5d",
			2888 => x"02009704",
			2889 => x"fef62d5d",
			2890 => x"00c62d5d",
			2891 => x"0c001b04",
			2892 => x"fe0e2d5d",
			2893 => x"ffe02d5d",
			2894 => x"08001d04",
			2895 => x"01cb2d5d",
			2896 => x"0000d704",
			2897 => x"ff692d5d",
			2898 => x"05006104",
			2899 => x"01422d5d",
			2900 => x"01f82d5d",
			2901 => x"fe6f2d5d",
			2902 => x"fe572d5d",
			2903 => x"0b001720",
			2904 => x"05004918",
			2905 => x"07002508",
			2906 => x"05003c04",
			2907 => x"ffc92e21",
			2908 => x"00842e21",
			2909 => x"0000b404",
			2910 => x"ff412e21",
			2911 => x"0200e208",
			2912 => x"03002904",
			2913 => x"fff02e21",
			2914 => x"008f2e21",
			2915 => x"ffa92e21",
			2916 => x"05004f04",
			2917 => x"00c22e21",
			2918 => x"00052e21",
			2919 => x"08001804",
			2920 => x"00562e21",
			2921 => x"0c001914",
			2922 => x"09001d04",
			2923 => x"00572e21",
			2924 => x"07002c08",
			2925 => x"0f005c04",
			2926 => x"ffe62e21",
			2927 => x"ff162e21",
			2928 => x"06009d04",
			2929 => x"00572e21",
			2930 => x"fff32e21",
			2931 => x"03003b10",
			2932 => x"0400390c",
			2933 => x"0b001808",
			2934 => x"0f006d04",
			2935 => x"fff82e21",
			2936 => x"005c2e21",
			2937 => x"ff5e2e21",
			2938 => x"00d12e21",
			2939 => x"07002f0c",
			2940 => x"0a004808",
			2941 => x"04003c04",
			2942 => x"00252e21",
			2943 => x"ff382e21",
			2944 => x"00302e21",
			2945 => x"0d001b08",
			2946 => x"03005c04",
			2947 => x"00872e21",
			2948 => x"fff12e21",
			2949 => x"0000e704",
			2950 => x"000f2e21",
			2951 => x"ffb72e21",
			2952 => x"05003c04",
			2953 => x"fe802ecf",
			2954 => x"0b001714",
			2955 => x"0500490c",
			2956 => x"07002304",
			2957 => x"01682ecf",
			2958 => x"0000b704",
			2959 => x"fec52ecf",
			2960 => x"00db2ecf",
			2961 => x"07002904",
			2962 => x"01792ecf",
			2963 => x"008c2ecf",
			2964 => x"05005120",
			2965 => x"03003e18",
			2966 => x"0a003d0c",
			2967 => x"01000804",
			2968 => x"00b42ecf",
			2969 => x"0000b904",
			2970 => x"fe832ecf",
			2971 => x"ffa62ecf",
			2972 => x"0c001b04",
			2973 => x"fe812ecf",
			2974 => x"0600a104",
			2975 => x"ffdb2ecf",
			2976 => x"ff972ecf",
			2977 => x"04003604",
			2978 => x"014b2ecf",
			2979 => x"ffac2ecf",
			2980 => x"08001c0c",
			2981 => x"04004708",
			2982 => x"09002104",
			2983 => x"01cb2ecf",
			2984 => x"00b42ecf",
			2985 => x"ff612ecf",
			2986 => x"07002f04",
			2987 => x"fe9e2ecf",
			2988 => x"0a005908",
			2989 => x"06008c04",
			2990 => x"01632ecf",
			2991 => x"00252ecf",
			2992 => x"01000b04",
			2993 => x"fffd2ecf",
			2994 => x"fee92ecf",
			2995 => x"0d00152c",
			2996 => x"0300351c",
			2997 => x"07002508",
			2998 => x"05003c04",
			2999 => x"ffe92f71",
			3000 => x"00402f71",
			3001 => x"01000508",
			3002 => x"09001e04",
			3003 => x"fff92f71",
			3004 => x"00322f71",
			3005 => x"0c001904",
			3006 => x"ff8d2f71",
			3007 => x"09002004",
			3008 => x"fffd2f71",
			3009 => x"00092f71",
			3010 => x"0c001a08",
			3011 => x"08001c04",
			3012 => x"00972f71",
			3013 => x"00132f71",
			3014 => x"0c001b04",
			3015 => x"ffc72f71",
			3016 => x"002d2f71",
			3017 => x"0c001a0c",
			3018 => x"0b001608",
			3019 => x"06006f04",
			3020 => x"00162f71",
			3021 => x"fff52f71",
			3022 => x"ff822f71",
			3023 => x"08001d10",
			3024 => x"0400490c",
			3025 => x"0a003b08",
			3026 => x"07002a04",
			3027 => x"ffd52f71",
			3028 => x"00052f71",
			3029 => x"00732f71",
			3030 => x"ffd82f71",
			3031 => x"05005e04",
			3032 => x"ffbf2f71",
			3033 => x"0a005904",
			3034 => x"002a2f71",
			3035 => x"ffdf2f71",
			3036 => x"0100071c",
			3037 => x"05004914",
			3038 => x"0f006604",
			3039 => x"ffa93005",
			3040 => x"0000e108",
			3041 => x"0a002c04",
			3042 => x"fffb3005",
			3043 => x"005a3005",
			3044 => x"07002e04",
			3045 => x"ffc13005",
			3046 => x"000b3005",
			3047 => x"04004304",
			3048 => x"00ab3005",
			3049 => x"ffd23005",
			3050 => x"07002508",
			3051 => x"05003c04",
			3052 => x"ffec3005",
			3053 => x"005f3005",
			3054 => x"0a004718",
			3055 => x"0f005d08",
			3056 => x"0f005904",
			3057 => x"ffe53005",
			3058 => x"001c3005",
			3059 => x"0400400c",
			3060 => x"07002e04",
			3061 => x"ff8c3005",
			3062 => x"07003504",
			3063 => x"001a3005",
			3064 => x"ffea3005",
			3065 => x"fffa3005",
			3066 => x"0a005908",
			3067 => x"08002304",
			3068 => x"005d3005",
			3069 => x"fff63005",
			3070 => x"01000b04",
			3071 => x"00013005",
			3072 => x"ffd93005",
			3073 => x"0b001720",
			3074 => x"05004918",
			3075 => x"07002508",
			3076 => x"05003c04",
			3077 => x"ffc430b1",
			3078 => x"00a230b1",
			3079 => x"0200ad04",
			3080 => x"ff2f30b1",
			3081 => x"0200e208",
			3082 => x"03002904",
			3083 => x"ffec30b1",
			3084 => x"009c30b1",
			3085 => x"ff9d30b1",
			3086 => x"05004f04",
			3087 => x"00cc30b1",
			3088 => x"000730b1",
			3089 => x"05004f1c",
			3090 => x"0000ae08",
			3091 => x"09001d04",
			3092 => x"006230b1",
			3093 => x"fef230b1",
			3094 => x"0e005b08",
			3095 => x"0200ba04",
			3096 => x"00d330b1",
			3097 => x"ffc530b1",
			3098 => x"07002c04",
			3099 => x"ff6b30b1",
			3100 => x"08001c04",
			3101 => x"007730b1",
			3102 => x"ffb130b1",
			3103 => x"09002108",
			3104 => x"06006904",
			3105 => x"00f430b1",
			3106 => x"000330b1",
			3107 => x"07002f08",
			3108 => x"0a004804",
			3109 => x"ff5d30b1",
			3110 => x"004f30b1",
			3111 => x"0a005908",
			3112 => x"00010704",
			3113 => x"009930b1",
			3114 => x"000130b1",
			3115 => x"ffba30b1",
			3116 => x"0d001538",
			3117 => x"0300351c",
			3118 => x"07002508",
			3119 => x"05003e04",
			3120 => x"ff993175",
			3121 => x"00e13175",
			3122 => x"01000508",
			3123 => x"09001e04",
			3124 => x"ffa03175",
			3125 => x"00c53175",
			3126 => x"0c001904",
			3127 => x"feb53175",
			3128 => x"0000b504",
			3129 => x"ff6f3175",
			3130 => x"009b3175",
			3131 => x"09002114",
			3132 => x"01000408",
			3133 => x"0000c604",
			3134 => x"00613175",
			3135 => x"ff503175",
			3136 => x"0b001808",
			3137 => x"09001f04",
			3138 => x"01583175",
			3139 => x"00973175",
			3140 => x"00183175",
			3141 => x"0000c704",
			3142 => x"ff2e3175",
			3143 => x"00ba3175",
			3144 => x"0c001a10",
			3145 => x"0b001608",
			3146 => x"0a003204",
			3147 => x"ffb93175",
			3148 => x"00743175",
			3149 => x"09002104",
			3150 => x"feb03175",
			3151 => x"ffaa3175",
			3152 => x"08001d10",
			3153 => x"0a003b08",
			3154 => x"01000704",
			3155 => x"00223175",
			3156 => x"ff0c3175",
			3157 => x"04004904",
			3158 => x"012e3175",
			3159 => x"ff773175",
			3160 => x"04004804",
			3161 => x"ff0a3175",
			3162 => x"0a005904",
			3163 => x"006c3175",
			3164 => x"ff8a3175",
			3165 => x"0d001524",
			3166 => x"03003914",
			3167 => x"0a003d10",
			3168 => x"04002b04",
			3169 => x"ff403219",
			3170 => x"0e004d04",
			3171 => x"01093219",
			3172 => x"07002904",
			3173 => x"ff443219",
			3174 => x"00cb3219",
			3175 => x"ff543219",
			3176 => x"0d001408",
			3177 => x"01000504",
			3178 => x"ffff3219",
			3179 => x"01053219",
			3180 => x"0200c404",
			3181 => x"ff6d3219",
			3182 => x"006a3219",
			3183 => x"0b001910",
			3184 => x"0b001608",
			3185 => x"01000b04",
			3186 => x"006a3219",
			3187 => x"ffb83219",
			3188 => x"07002e04",
			3189 => x"fed03219",
			3190 => x"ffc33219",
			3191 => x"0a003b04",
			3192 => x"ff083219",
			3193 => x"03003b08",
			3194 => x"04003504",
			3195 => x"ffce3219",
			3196 => x"01203219",
			3197 => x"0200b904",
			3198 => x"ff2d3219",
			3199 => x"0d001b08",
			3200 => x"04004c04",
			3201 => x"00ce3219",
			3202 => x"ffdb3219",
			3203 => x"01000d04",
			3204 => x"00173219",
			3205 => x"ff773219",
			3206 => x"0d001534",
			3207 => x"0e00651c",
			3208 => x"05004610",
			3209 => x"06005f0c",
			3210 => x"07002408",
			3211 => x"05003904",
			3212 => x"ffee32d5",
			3213 => x"002632d5",
			3214 => x"ffbd32d5",
			3215 => x"001232d5",
			3216 => x"0b001804",
			3217 => x"006732d5",
			3218 => x"0000b904",
			3219 => x"ffdb32d5",
			3220 => x"002b32d5",
			3221 => x"07002b0c",
			3222 => x"03003108",
			3223 => x"03002c04",
			3224 => x"fffb32d5",
			3225 => x"001132d5",
			3226 => x"ffa932d5",
			3227 => x"0000cd04",
			3228 => x"ffd332d5",
			3229 => x"09001e04",
			3230 => x"fff032d5",
			3231 => x"004e32d5",
			3232 => x"01000708",
			3233 => x"08001c04",
			3234 => x"004032d5",
			3235 => x"ffea32d5",
			3236 => x"0a004714",
			3237 => x"0b001608",
			3238 => x"06006f04",
			3239 => x"001432d5",
			3240 => x"fff732d5",
			3241 => x"07003004",
			3242 => x"ff6432d5",
			3243 => x"0f009f04",
			3244 => x"001532d5",
			3245 => x"ffeb32d5",
			3246 => x"0a00590c",
			3247 => x"0f007204",
			3248 => x"fffb32d5",
			3249 => x"0f00a204",
			3250 => x"003d32d5",
			3251 => x"fffd32d5",
			3252 => x"ffde32d5",
			3253 => x"0000ed3c",
			3254 => x"0b00171c",
			3255 => x"05004914",
			3256 => x"07002508",
			3257 => x"05003c04",
			3258 => x"ffbe3361",
			3259 => x"00c13361",
			3260 => x"0000b404",
			3261 => x"ff1d3361",
			3262 => x"03002904",
			3263 => x"ffe63361",
			3264 => x"00983361",
			3265 => x"04003d04",
			3266 => x"01013361",
			3267 => x"ffdf3361",
			3268 => x"02009704",
			3269 => x"ff113361",
			3270 => x"0000a808",
			3271 => x"0d001704",
			3272 => x"00c53361",
			3273 => x"ffea3361",
			3274 => x"0c001908",
			3275 => x"07002b04",
			3276 => x"ff113361",
			3277 => x"005a3361",
			3278 => x"0000ad04",
			3279 => x"ff533361",
			3280 => x"03004004",
			3281 => x"00d33361",
			3282 => x"ffce3361",
			3283 => x"05005004",
			3284 => x"ff303361",
			3285 => x"0a004f04",
			3286 => x"004c3361",
			3287 => x"ffcc3361",
			3288 => x"0d001530",
			3289 => x"03003e24",
			3290 => x"0000df20",
			3291 => x"0000b414",
			3292 => x"07002508",
			3293 => x"05003c04",
			3294 => x"ffad3405",
			3295 => x"00e13405",
			3296 => x"01000504",
			3297 => x"004f3405",
			3298 => x"0c001b04",
			3299 => x"ff203405",
			3300 => x"00583405",
			3301 => x"0d001408",
			3302 => x"04002d04",
			3303 => x"ffef3405",
			3304 => x"012d3405",
			3305 => x"00093405",
			3306 => x"fef63405",
			3307 => x"04003e04",
			3308 => x"010a3405",
			3309 => x"0c001a04",
			3310 => x"ff6c3405",
			3311 => x"00a53405",
			3312 => x"0200b90c",
			3313 => x"01000704",
			3314 => x"00503405",
			3315 => x"0c001604",
			3316 => x"fff53405",
			3317 => x"fea13405",
			3318 => x"0b001904",
			3319 => x"ff3d3405",
			3320 => x"01000d0c",
			3321 => x"03006108",
			3322 => x"04003404",
			3323 => x"ffec3405",
			3324 => x"010a3405",
			3325 => x"ffde3405",
			3326 => x"08002004",
			3327 => x"00313405",
			3328 => x"ff4e3405",
			3329 => x"0d001530",
			3330 => x"03003920",
			3331 => x"0a003d1c",
			3332 => x"03003518",
			3333 => x"07002508",
			3334 => x"05003c04",
			3335 => x"ff9f34b1",
			3336 => x"00e634b1",
			3337 => x"07002a08",
			3338 => x"09002004",
			3339 => x"fef134b1",
			3340 => x"001a34b1",
			3341 => x"06008004",
			3342 => x"00a734b1",
			3343 => x"ff8334b1",
			3344 => x"00dd34b1",
			3345 => x"ff4634b1",
			3346 => x"0d001408",
			3347 => x"0000cf04",
			3348 => x"011d34b1",
			3349 => x"001034b1",
			3350 => x"0200c404",
			3351 => x"ff6134b1",
			3352 => x"007534b1",
			3353 => x"0b001910",
			3354 => x"0b001608",
			3355 => x"01000b04",
			3356 => x"006e34b1",
			3357 => x"ffb434b1",
			3358 => x"07002e04",
			3359 => x"fec534b1",
			3360 => x"ffbb34b1",
			3361 => x"0a003b04",
			3362 => x"fefe34b1",
			3363 => x"05005308",
			3364 => x"01000e04",
			3365 => x"013034b1",
			3366 => x"ff9834b1",
			3367 => x"0a004704",
			3368 => x"ff4b34b1",
			3369 => x"0a005904",
			3370 => x"00a334b1",
			3371 => x"ff8834b1",
			3372 => x"05003c04",
			3373 => x"fe783525",
			3374 => x"09001e0c",
			3375 => x"05004708",
			3376 => x"07002504",
			3377 => x"01833525",
			3378 => x"ff0c3525",
			3379 => x"01cb3525",
			3380 => x"0000c010",
			3381 => x"0e005b0c",
			3382 => x"0000ae08",
			3383 => x"05004b04",
			3384 => x"fe5e3525",
			3385 => x"00943525",
			3386 => x"01453525",
			3387 => x"fe6d3525",
			3388 => x"0e006508",
			3389 => x"0d001904",
			3390 => x"017b3525",
			3391 => x"ff113525",
			3392 => x"03003308",
			3393 => x"0f00c404",
			3394 => x"018e3525",
			3395 => x"ffcc3525",
			3396 => x"09002004",
			3397 => x"fec63525",
			3398 => x"04004704",
			3399 => x"00d83525",
			3400 => x"ff5f3525",
			3401 => x"01000938",
			3402 => x"08001b1c",
			3403 => x"05004818",
			3404 => x"07002910",
			3405 => x"07002308",
			3406 => x"09001a04",
			3407 => x"fff035d9",
			3408 => x"002635d9",
			3409 => x"06005f04",
			3410 => x"ff9d35d9",
			3411 => x"fffb35d9",
			3412 => x"0000f204",
			3413 => x"004b35d9",
			3414 => x"ffe535d9",
			3415 => x"00c535d9",
			3416 => x"05004d14",
			3417 => x"0f00640c",
			3418 => x"01000808",
			3419 => x"08001c04",
			3420 => x"000b35d9",
			3421 => x"ffb435d9",
			3422 => x"002835d9",
			3423 => x"05004204",
			3424 => x"fff535d9",
			3425 => x"008135d9",
			3426 => x"0c001b04",
			3427 => x"ff8235d9",
			3428 => x"002b35d9",
			3429 => x"09001e08",
			3430 => x"05003f04",
			3431 => x"ffd635d9",
			3432 => x"007235d9",
			3433 => x"04004314",
			3434 => x"0000c704",
			3435 => x"ff2b35d9",
			3436 => x"0201030c",
			3437 => x"03003a08",
			3438 => x"0000dd04",
			3439 => x"000535d9",
			3440 => x"ffe835d9",
			3441 => x"004835d9",
			3442 => x"ffcc35d9",
			3443 => x"0a005904",
			3444 => x"005235d9",
			3445 => x"ffd335d9",
			3446 => x"01000930",
			3447 => x"08001d20",
			3448 => x"04003818",
			3449 => x"04003614",
			3450 => x"0000e008",
			3451 => x"04002b04",
			3452 => x"ffe9369d",
			3453 => x"0066369d",
			3454 => x"07002c04",
			3455 => x"ffc0369d",
			3456 => x"07002f04",
			3457 => x"0023369d",
			3458 => x"fff9369d",
			3459 => x"ffc6369d",
			3460 => x"0c001b04",
			3461 => x"00a5369d",
			3462 => x"fffc369d",
			3463 => x"07002704",
			3464 => x"0017369d",
			3465 => x"0a003d08",
			3466 => x"09002204",
			3467 => x"000c369d",
			3468 => x"fffc369d",
			3469 => x"ffac369d",
			3470 => x"04004320",
			3471 => x"0200be10",
			3472 => x"09001e0c",
			3473 => x"00008804",
			3474 => x"fff4369d",
			3475 => x"06005604",
			3476 => x"003c369d",
			3477 => x"fffe369d",
			3478 => x"ff5f369d",
			3479 => x"0201010c",
			3480 => x"0a003b04",
			3481 => x"ffed369d",
			3482 => x"06006a04",
			3483 => x"fffe369d",
			3484 => x"0054369d",
			3485 => x"ffd4369d",
			3486 => x"04004b08",
			3487 => x"07003204",
			3488 => x"0056369d",
			3489 => x"fffb369d",
			3490 => x"0e007104",
			3491 => x"ffbd369d",
			3492 => x"07003e04",
			3493 => x"001c369d",
			3494 => x"fffa369d",
			3495 => x"08001d4c",
			3496 => x"0e005f2c",
			3497 => x"0c001918",
			3498 => x"09001f10",
			3499 => x"0500460c",
			3500 => x"07002508",
			3501 => x"05003e04",
			3502 => x"ffa73759",
			3503 => x"00db3759",
			3504 => x"ff783759",
			3505 => x"010a3759",
			3506 => x"0000b504",
			3507 => x"ff053759",
			3508 => x"00e73759",
			3509 => x"0400370c",
			3510 => x"03003208",
			3511 => x"00009b04",
			3512 => x"ffec3759",
			3513 => x"00703759",
			3514 => x"ff653759",
			3515 => x"0c001a04",
			3516 => x"00733759",
			3517 => x"013f3759",
			3518 => x"0000d00c",
			3519 => x"04003c08",
			3520 => x"0000c504",
			3521 => x"ff9d3759",
			3522 => x"00943759",
			3523 => x"fee43759",
			3524 => x"09002010",
			3525 => x"01000508",
			3526 => x"05003404",
			3527 => x"ffe13759",
			3528 => x"00bc3759",
			3529 => x"0000dd04",
			3530 => x"002e3759",
			3531 => x"fef53759",
			3532 => x"01403759",
			3533 => x"0d001408",
			3534 => x"01000c04",
			3535 => x"ffd53759",
			3536 => x"00b43759",
			3537 => x"05005e04",
			3538 => x"fee03759",
			3539 => x"03005304",
			3540 => x"00693759",
			3541 => x"ff803759",
			3542 => x"04002b04",
			3543 => x"fea637d5",
			3544 => x"08001d20",
			3545 => x"0a004518",
			3546 => x"0a004210",
			3547 => x"0000e10c",
			3548 => x"0000c008",
			3549 => x"06006404",
			3550 => x"00a737d5",
			3551 => x"fea737d5",
			3552 => x"016f37d5",
			3553 => x"ff4d37d5",
			3554 => x"0b001804",
			3555 => x"009037d5",
			3556 => x"fece37d5",
			3557 => x"09002504",
			3558 => x"016137d5",
			3559 => x"002c37d5",
			3560 => x"0c001a04",
			3561 => x"002437d5",
			3562 => x"05005e0c",
			3563 => x"07003304",
			3564 => x"fea337d5",
			3565 => x"00011204",
			3566 => x"008137d5",
			3567 => x"ff5337d5",
			3568 => x"0a005904",
			3569 => x"00b237d5",
			3570 => x"0d001b04",
			3571 => x"fff537d5",
			3572 => x"ff4237d5",
			3573 => x"05005248",
			3574 => x"0e005b20",
			3575 => x"0f006818",
			3576 => x"09001d08",
			3577 => x"05003c04",
			3578 => x"ffe13891",
			3579 => x"00723891",
			3580 => x"05004b0c",
			3581 => x"06005d08",
			3582 => x"07002304",
			3583 => x"00143891",
			3584 => x"ff3b3891",
			3585 => x"00133891",
			3586 => x"00313891",
			3587 => x"01000804",
			3588 => x"ffed3891",
			3589 => x"00873891",
			3590 => x"0200bb0c",
			3591 => x"0d001204",
			3592 => x"00043891",
			3593 => x"05004704",
			3594 => x"00003891",
			3595 => x"ff5e3891",
			3596 => x"0200ee10",
			3597 => x"05004d0c",
			3598 => x"03003508",
			3599 => x"0000df04",
			3600 => x"00293891",
			3601 => x"ffc23891",
			3602 => x"006e3891",
			3603 => x"ffe73891",
			3604 => x"0c001c04",
			3605 => x"ffa03891",
			3606 => x"03003a04",
			3607 => x"fff53891",
			3608 => x"00113891",
			3609 => x"08001c08",
			3610 => x"06007504",
			3611 => x"009a3891",
			3612 => x"fffd3891",
			3613 => x"07002f04",
			3614 => x"ffb03891",
			3615 => x"0a005904",
			3616 => x"00523891",
			3617 => x"01000b04",
			3618 => x"00013891",
			3619 => x"ffd63891",
			3620 => x"0d001544",
			3621 => x"05004930",
			3622 => x"0d00131c",
			3623 => x"07002308",
			3624 => x"05003e04",
			3625 => x"ffb73975",
			3626 => x"00993975",
			3627 => x"07002c0c",
			3628 => x"05003d08",
			3629 => x"03002f04",
			3630 => x"ffb03975",
			3631 => x"004a3975",
			3632 => x"fede3975",
			3633 => x"06009104",
			3634 => x"004d3975",
			3635 => x"ffcf3975",
			3636 => x"0200970c",
			3637 => x"07002408",
			3638 => x"00007804",
			3639 => x"fff13975",
			3640 => x"00713975",
			3641 => x"ff293975",
			3642 => x"04002d04",
			3643 => x"ff683975",
			3644 => x"01113975",
			3645 => x"04003c08",
			3646 => x"0000b804",
			3647 => x"009a3975",
			3648 => x"013e3975",
			3649 => x"0e006108",
			3650 => x"0b001804",
			3651 => x"00d13975",
			3652 => x"ffaf3975",
			3653 => x"ff323975",
			3654 => x"0c001a10",
			3655 => x"0b001608",
			3656 => x"0a003204",
			3657 => x"ffbb3975",
			3658 => x"006d3975",
			3659 => x"09002104",
			3660 => x"feba3975",
			3661 => x"ffa83975",
			3662 => x"08001d10",
			3663 => x"0a003b08",
			3664 => x"01000704",
			3665 => x"00203975",
			3666 => x"ff1a3975",
			3667 => x"04004904",
			3668 => x"011f3975",
			3669 => x"ff823975",
			3670 => x"04004804",
			3671 => x"ff183975",
			3672 => x"0f007204",
			3673 => x"ff8d3975",
			3674 => x"0a005904",
			3675 => x"00b43975",
			3676 => x"ffa43975",
			3677 => x"0d00142c",
			3678 => x"05004924",
			3679 => x"07002510",
			3680 => x"05003e0c",
			3681 => x"01000704",
			3682 => x"ffe53a41",
			3683 => x"01000804",
			3684 => x"000a3a41",
			3685 => x"fff93a41",
			3686 => x"003a3a41",
			3687 => x"06005e04",
			3688 => x"ff983a41",
			3689 => x"0b001608",
			3690 => x"0d001304",
			3691 => x"ffd83a41",
			3692 => x"00033a41",
			3693 => x"06008104",
			3694 => x"00413a41",
			3695 => x"fff53a41",
			3696 => x"09002104",
			3697 => x"00803a41",
			3698 => x"00033a41",
			3699 => x"0000ca18",
			3700 => x"07002608",
			3701 => x"00008f04",
			3702 => x"fff33a41",
			3703 => x"00373a41",
			3704 => x"03003308",
			3705 => x"09001f04",
			3706 => x"ffd93a41",
			3707 => x"00323a41",
			3708 => x"0a004704",
			3709 => x"ff563a41",
			3710 => x"000d3a41",
			3711 => x"0e006908",
			3712 => x"0f007304",
			3713 => x"ffe73a41",
			3714 => x"00683a41",
			3715 => x"0c001b0c",
			3716 => x"0a003908",
			3717 => x"0a003604",
			3718 => x"fff53a41",
			3719 => x"000a3a41",
			3720 => x"ffb13a41",
			3721 => x"0201020c",
			3722 => x"03005c08",
			3723 => x"0a003d04",
			3724 => x"fffe3a41",
			3725 => x"00493a41",
			3726 => x"fff13a41",
			3727 => x"ffe63a41",
			3728 => x"05003c04",
			3729 => x"fe653aad",
			3730 => x"0800232c",
			3731 => x"0a00451c",
			3732 => x"07002504",
			3733 => x"01a33aad",
			3734 => x"0000a608",
			3735 => x"0c001904",
			3736 => x"ffc43aad",
			3737 => x"fe3d3aad",
			3738 => x"0e005b08",
			3739 => x"0f006804",
			3740 => x"00173aad",
			3741 => x"025c3aad",
			3742 => x"0200bb04",
			3743 => x"fea53aad",
			3744 => x"00a03aad",
			3745 => x"03005c0c",
			3746 => x"08001d04",
			3747 => x"01b73aad",
			3748 => x"09002504",
			3749 => x"ff943aad",
			3750 => x"01df3aad",
			3751 => x"fe883aad",
			3752 => x"01001004",
			3753 => x"ffd13aad",
			3754 => x"fe693aad",
			3755 => x"0d001538",
			3756 => x"0200d82c",
			3757 => x"0000b418",
			3758 => x"0e005710",
			3759 => x"0500460c",
			3760 => x"07002508",
			3761 => x"05003c04",
			3762 => x"ffe63b81",
			3763 => x"00413b81",
			3764 => x"ffa33b81",
			3765 => x"00633b81",
			3766 => x"0d001204",
			3767 => x"00043b81",
			3768 => x"ff9b3b81",
			3769 => x"0e00680c",
			3770 => x"01000404",
			3771 => x"fffb3b81",
			3772 => x"04002d04",
			3773 => x"fffb3b81",
			3774 => x"00b23b81",
			3775 => x"01000604",
			3776 => x"ffe43b81",
			3777 => x"00013b81",
			3778 => x"07002b04",
			3779 => x"ffa83b81",
			3780 => x"03003304",
			3781 => x"fff03b81",
			3782 => x"001e3b81",
			3783 => x"0c001a0c",
			3784 => x"0b001608",
			3785 => x"06006f04",
			3786 => x"001b3b81",
			3787 => x"fff23b81",
			3788 => x"ff723b81",
			3789 => x"01000b18",
			3790 => x"0a003b08",
			3791 => x"08001b04",
			3792 => x"00093b81",
			3793 => x"ffc23b81",
			3794 => x"05005904",
			3795 => x"008f3b81",
			3796 => x"03004904",
			3797 => x"ffce3b81",
			3798 => x"05009a04",
			3799 => x"00273b81",
			3800 => x"fff93b81",
			3801 => x"0d001808",
			3802 => x"0000ce04",
			3803 => x"fff03b81",
			3804 => x"00253b81",
			3805 => x"0000c404",
			3806 => x"00123b81",
			3807 => x"ffa13b81",
			3808 => x"05003c04",
			3809 => x"fe8c3c0d",
			3810 => x"0d001520",
			3811 => x"0300350c",
			3812 => x"07002504",
			3813 => x"01603c0d",
			3814 => x"0000b504",
			3815 => x"feb23c0d",
			3816 => x"00053c0d",
			3817 => x"0100090c",
			3818 => x"0f006404",
			3819 => x"00773c0d",
			3820 => x"0b001604",
			3821 => x"00af3c0d",
			3822 => x"01963c0d",
			3823 => x"0000b904",
			3824 => x"ffed3c0d",
			3825 => x"013c3c0d",
			3826 => x"04003c0c",
			3827 => x"07002e04",
			3828 => x"fe803c0d",
			3829 => x"00010f04",
			3830 => x"00ab3c0d",
			3831 => x"feeb3c0d",
			3832 => x"03003e04",
			3833 => x"012c3c0d",
			3834 => x"0200b904",
			3835 => x"fe853c0d",
			3836 => x"0e006908",
			3837 => x"08001f04",
			3838 => x"01103c0d",
			3839 => x"ff4e3c0d",
			3840 => x"0f008104",
			3841 => x"fe863c0d",
			3842 => x"00a63c0d",
			3843 => x"0400310c",
			3844 => x"05003c04",
			3845 => x"fe463c81",
			3846 => x"0000f204",
			3847 => x"02df3c81",
			3848 => x"fe443c81",
			3849 => x"0d001b2c",
			3850 => x"04006128",
			3851 => x"0a004318",
			3852 => x"0d00150c",
			3853 => x"07002504",
			3854 => x"052a3c81",
			3855 => x"0000a604",
			3856 => x"00683c81",
			3857 => x"04383c81",
			3858 => x"0000cd08",
			3859 => x"0e005a04",
			3860 => x"00923c81",
			3861 => x"fe353c81",
			3862 => x"02f33c81",
			3863 => x"0700360c",
			3864 => x"07002a04",
			3865 => x"05223c81",
			3866 => x"0000c704",
			3867 => x"03233c81",
			3868 => x"046c3c81",
			3869 => x"05e73c81",
			3870 => x"fe483c81",
			3871 => x"fe473c81",
			3872 => x"0e006b40",
			3873 => x"0f007c38",
			3874 => x"09001e10",
			3875 => x"0500450c",
			3876 => x"04003108",
			3877 => x"03002c04",
			3878 => x"ff8d3d35",
			3879 => x"00e33d35",
			3880 => x"ff4e3d35",
			3881 => x"01553d35",
			3882 => x"0a003b0c",
			3883 => x"0000b704",
			3884 => x"fea23d35",
			3885 => x"0d001504",
			3886 => x"00763d35",
			3887 => x"ff7e3d35",
			3888 => x"0e006310",
			3889 => x"0000ad08",
			3890 => x"05004b04",
			3891 => x"feeb3d35",
			3892 => x"00623d35",
			3893 => x"0c001904",
			3894 => x"ff923d35",
			3895 => x"00d23d35",
			3896 => x"0000d004",
			3897 => x"fee43d35",
			3898 => x"07003204",
			3899 => x"00ea3d35",
			3900 => x"ffbe3d35",
			3901 => x"04002d04",
			3902 => x"ffbd3d35",
			3903 => x"01553d35",
			3904 => x"0c001b0c",
			3905 => x"08001908",
			3906 => x"08001804",
			3907 => x"ffa63d35",
			3908 => x"003a3d35",
			3909 => x"feb13d35",
			3910 => x"0201030c",
			3911 => x"03006108",
			3912 => x"04003604",
			3913 => x"ffe03d35",
			3914 => x"00eb3d35",
			3915 => x"ffbb3d35",
			3916 => x"ff423d35",
			3917 => x"0500410c",
			3918 => x"05003c04",
			3919 => x"fe523dc1",
			3920 => x"0b001704",
			3921 => x"01773dc1",
			3922 => x"fe4e3dc1",
			3923 => x"0d001b30",
			3924 => x"03005c2c",
			3925 => x"05004f18",
			3926 => x"0b00170c",
			3927 => x"05004908",
			3928 => x"07002504",
			3929 => x"032b3dc1",
			3930 => x"00fb3dc1",
			3931 => x"03593dc1",
			3932 => x"0f006404",
			3933 => x"fe1a3dc1",
			3934 => x"0e005b04",
			3935 => x"02c53dc1",
			3936 => x"00ae3dc1",
			3937 => x"0000c708",
			3938 => x"09002104",
			3939 => x"03203dc1",
			3940 => x"00193dc1",
			3941 => x"03004104",
			3942 => x"031b3dc1",
			3943 => x"03004504",
			3944 => x"023e3dc1",
			3945 => x"02dd3dc1",
			3946 => x"fe663dc1",
			3947 => x"01000d08",
			3948 => x"0500b604",
			3949 => x"01993dc1",
			3950 => x"fe643dc1",
			3951 => x"fe523dc1",
			3952 => x"0e006530",
			3953 => x"0000b920",
			3954 => x"0600641c",
			3955 => x"08001d14",
			3956 => x"0000ad10",
			3957 => x"09001e08",
			3958 => x"00008104",
			3959 => x"ff3a3e95",
			3960 => x"011e3e95",
			3961 => x"05004b04",
			3962 => x"fed93e95",
			3963 => x"006a3e95",
			3964 => x"00cc3e95",
			3965 => x"09001d04",
			3966 => x"000e3e95",
			3967 => x"fed23e95",
			3968 => x"fed63e95",
			3969 => x"07002704",
			3970 => x"ff683e95",
			3971 => x"0d001908",
			3972 => x"0000c004",
			3973 => x"00513e95",
			3974 => x"01523e95",
			3975 => x"ff8a3e95",
			3976 => x"0a00482c",
			3977 => x"08001b1c",
			3978 => x"0000e108",
			3979 => x"0000d004",
			3980 => x"ff8c3e95",
			3981 => x"01183e95",
			3982 => x"01000508",
			3983 => x"07002b04",
			3984 => x"ffe43e95",
			3985 => x"005e3e95",
			3986 => x"0d001304",
			3987 => x"fed53e95",
			3988 => x"07002c04",
			3989 => x"00313e95",
			3990 => x"ff9a3e95",
			3991 => x"0c001b08",
			3992 => x"0b001904",
			3993 => x"fe933e95",
			3994 => x"ffc73e95",
			3995 => x"00010c04",
			3996 => x"00653e95",
			3997 => x"ff5b3e95",
			3998 => x"0a005908",
			3999 => x"00010304",
			4000 => x"00d83e95",
			4001 => x"00133e95",
			4002 => x"0d001b04",
			4003 => x"001f3e95",
			4004 => x"ff723e95",
			4005 => x"05004934",
			4006 => x"0d001314",
			4007 => x"07002508",
			4008 => x"05003e04",
			4009 => x"ffbe3f61",
			4010 => x"006c3f61",
			4011 => x"05003d08",
			4012 => x"05003604",
			4013 => x"ffd23f61",
			4014 => x"00353f61",
			4015 => x"ff0b3f61",
			4016 => x"0a003b18",
			4017 => x"0700260c",
			4018 => x"09001e08",
			4019 => x"00008b04",
			4020 => x"ffe93f61",
			4021 => x"00a33f61",
			4022 => x"ffc03f61",
			4023 => x"01000608",
			4024 => x"0000c304",
			4025 => x"fff03f61",
			4026 => x"00433f61",
			4027 => x"ff143f61",
			4028 => x"0000dd04",
			4029 => x"00af3f61",
			4030 => x"ffa43f61",
			4031 => x"0d00140c",
			4032 => x"04003f08",
			4033 => x"01000704",
			4034 => x"00f43f61",
			4035 => x"00603f61",
			4036 => x"000a3f61",
			4037 => x"03003904",
			4038 => x"00783f61",
			4039 => x"0200ba08",
			4040 => x"03004004",
			4041 => x"ff093f61",
			4042 => x"ffd63f61",
			4043 => x"0e006a10",
			4044 => x"08001f08",
			4045 => x"04004904",
			4046 => x"008f3f61",
			4047 => x"00153f61",
			4048 => x"01000b04",
			4049 => x"000d3f61",
			4050 => x"ffbe3f61",
			4051 => x"0e007004",
			4052 => x"ff7b3f61",
			4053 => x"01001004",
			4054 => x"006e3f61",
			4055 => x"ffcd3f61",
			4056 => x"0b001720",
			4057 => x"05004918",
			4058 => x"07002508",
			4059 => x"05003c04",
			4060 => x"ffd44005",
			4061 => x"008c4005",
			4062 => x"0000b404",
			4063 => x"ff534005",
			4064 => x"0200e208",
			4065 => x"03002904",
			4066 => x"fff14005",
			4067 => x"00744005",
			4068 => x"ffb34005",
			4069 => x"05005004",
			4070 => x"00b64005",
			4071 => x"000d4005",
			4072 => x"02009704",
			4073 => x"ff5e4005",
			4074 => x"0000a808",
			4075 => x"0d001604",
			4076 => x"008f4005",
			4077 => x"ffe74005",
			4078 => x"0c00190c",
			4079 => x"07002b04",
			4080 => x"ff554005",
			4081 => x"0b001804",
			4082 => x"ffdb4005",
			4083 => x"005b4005",
			4084 => x"0100090c",
			4085 => x"0e006808",
			4086 => x"04003704",
			4087 => x"fff64005",
			4088 => x"00b14005",
			4089 => x"ff9a4005",
			4090 => x"0200b908",
			4091 => x"01000e04",
			4092 => x"ff554005",
			4093 => x"00104005",
			4094 => x"0d001b04",
			4095 => x"00574005",
			4096 => x"ffba4005",
			4097 => x"05003c04",
			4098 => x"fe6a4079",
			4099 => x"02010130",
			4100 => x"0b001710",
			4101 => x"05004908",
			4102 => x"07002304",
			4103 => x"01b44079",
			4104 => x"ffd04079",
			4105 => x"05004f04",
			4106 => x"01cb4079",
			4107 => x"006e4079",
			4108 => x"02009204",
			4109 => x"fe5c4079",
			4110 => x"0c001a0c",
			4111 => x"0d001508",
			4112 => x"0e005c04",
			4113 => x"016d4079",
			4114 => x"ffc54079",
			4115 => x"fe1f4079",
			4116 => x"0d001608",
			4117 => x"0b001904",
			4118 => x"00884079",
			4119 => x"01be4079",
			4120 => x"07002f04",
			4121 => x"ff0b4079",
			4122 => x"00f74079",
			4123 => x"05005204",
			4124 => x"fe6c4079",
			4125 => x"00414079",
			4126 => x"08001f4c",
			4127 => x"0a003614",
			4128 => x"07002508",
			4129 => x"05003b04",
			4130 => x"ffad4125",
			4131 => x"008c4125",
			4132 => x"09002004",
			4133 => x"ff1a4125",
			4134 => x"09002104",
			4135 => x"000b4125",
			4136 => x"fffb4125",
			4137 => x"0400472c",
			4138 => x"05004914",
			4139 => x"0d001308",
			4140 => x"07002a04",
			4141 => x"ff3a4125",
			4142 => x"00664125",
			4143 => x"0000ae04",
			4144 => x"fff94125",
			4145 => x"06007e04",
			4146 => x"00d84125",
			4147 => x"ffd64125",
			4148 => x"07002908",
			4149 => x"01000804",
			4150 => x"00544125",
			4151 => x"01154125",
			4152 => x"0000c708",
			4153 => x"01000904",
			4154 => x"00714125",
			4155 => x"ff364125",
			4156 => x"04004304",
			4157 => x"011d4125",
			4158 => x"ffba4125",
			4159 => x"07003004",
			4160 => x"ff684125",
			4161 => x"0b001d04",
			4162 => x"006c4125",
			4163 => x"fff34125",
			4164 => x"04004a04",
			4165 => x"ff274125",
			4166 => x"05008104",
			4167 => x"003f4125",
			4168 => x"ffbe4125",
			4169 => x"0b001710",
			4170 => x"05003c04",
			4171 => x"ffbb41c9",
			4172 => x"05004908",
			4173 => x"05004504",
			4174 => x"005641c9",
			4175 => x"ffc741c9",
			4176 => x"008541c9",
			4177 => x"05004f24",
			4178 => x"09001d04",
			4179 => x"002341c9",
			4180 => x"0000ae08",
			4181 => x"01000504",
			4182 => x"001b41c9",
			4183 => x"ff5341c9",
			4184 => x"06006508",
			4185 => x"0200b704",
			4186 => x"007041c9",
			4187 => x"ffe441c9",
			4188 => x"01000c08",
			4189 => x"07002c04",
			4190 => x"ff9341c9",
			4191 => x"000c41c9",
			4192 => x"01001004",
			4193 => x"001c41c9",
			4194 => x"ffe441c9",
			4195 => x"09002104",
			4196 => x"005c41c9",
			4197 => x"0000d008",
			4198 => x"0a004704",
			4199 => x"ff8c41c9",
			4200 => x"001c41c9",
			4201 => x"0a005908",
			4202 => x"00010704",
			4203 => x"004f41c9",
			4204 => x"fffc41c9",
			4205 => x"01000b04",
			4206 => x"000241c9",
			4207 => x"0200ce04",
			4208 => x"000041c9",
			4209 => x"ffdb41c9",
			4210 => x"04002b04",
			4211 => x"fe704255",
			4212 => x"0b001714",
			4213 => x"0000f210",
			4214 => x"0f006608",
			4215 => x"07002504",
			4216 => x"01734255",
			4217 => x"ffa34255",
			4218 => x"0a004204",
			4219 => x"01a94255",
			4220 => x"00fc4255",
			4221 => x"fefd4255",
			4222 => x"05004f18",
			4223 => x"0000ae04",
			4224 => x"fe554255",
			4225 => x"0a004210",
			4226 => x"0000dd08",
			4227 => x"03003a04",
			4228 => x"01b44255",
			4229 => x"fff74255",
			4230 => x"03003a04",
			4231 => x"fde64255",
			4232 => x"010a4255",
			4233 => x"fe3c4255",
			4234 => x"0d001408",
			4235 => x"0e006004",
			4236 => x"01a24255",
			4237 => x"00dc4255",
			4238 => x"0b001904",
			4239 => x"ff104255",
			4240 => x"03003e04",
			4241 => x"01ad4255",
			4242 => x"0200b904",
			4243 => x"fe774255",
			4244 => x"00ab4255",
			4245 => x"05003c04",
			4246 => x"fe6c42d9",
			4247 => x"08001d24",
			4248 => x"0200e720",
			4249 => x"0000d014",
			4250 => x"0e006110",
			4251 => x"0000b408",
			4252 => x"0e005a04",
			4253 => x"00a842d9",
			4254 => x"feac42d9",
			4255 => x"07002904",
			4256 => x"006242d9",
			4257 => x"01ae42d9",
			4258 => x"fe9b42d9",
			4259 => x"01000704",
			4260 => x"01c242d9",
			4261 => x"0000dd04",
			4262 => x"018442d9",
			4263 => x"ffc042d9",
			4264 => x"ff0542d9",
			4265 => x"0f007208",
			4266 => x"0f006004",
			4267 => x"002d42d9",
			4268 => x"fe4d42d9",
			4269 => x"0e006704",
			4270 => x"017042d9",
			4271 => x"0c001c04",
			4272 => x"fde542d9",
			4273 => x"0d001c08",
			4274 => x"03006104",
			4275 => x"016a42d9",
			4276 => x"ff1c42d9",
			4277 => x"fea242d9",
			4278 => x"0d001530",
			4279 => x"03003e28",
			4280 => x"0000df24",
			4281 => x"0b001814",
			4282 => x"0000b40c",
			4283 => x"0e005408",
			4284 => x"05004604",
			4285 => x"ffba4385",
			4286 => x"00fb4385",
			4287 => x"ff064385",
			4288 => x"04002d04",
			4289 => x"fff14385",
			4290 => x"00f84385",
			4291 => x"0c001b08",
			4292 => x"03003304",
			4293 => x"003f4385",
			4294 => x"ff384385",
			4295 => x"07002904",
			4296 => x"ffec4385",
			4297 => x"008b4385",
			4298 => x"ff0d4385",
			4299 => x"01000404",
			4300 => x"ffbf4385",
			4301 => x"00eb4385",
			4302 => x"06006208",
			4303 => x"0b001604",
			4304 => x"00434385",
			4305 => x"fedd4385",
			4306 => x"0b001904",
			4307 => x"ff394385",
			4308 => x"01000904",
			4309 => x"01084385",
			4310 => x"0a00470c",
			4311 => x"0c001b04",
			4312 => x"ff6c4385",
			4313 => x"05004404",
			4314 => x"ffbd4385",
			4315 => x"00274385",
			4316 => x"0a005908",
			4317 => x"04004304",
			4318 => x"fff54385",
			4319 => x"00824385",
			4320 => x"ffa74385",
			4321 => x"0000ed54",
			4322 => x"0000c72c",
			4323 => x"06006a24",
			4324 => x"09001d08",
			4325 => x"05003c04",
			4326 => x"ff3b4449",
			4327 => x"018e4449",
			4328 => x"0000b410",
			4329 => x"0a003b08",
			4330 => x"07002504",
			4331 => x"007c4449",
			4332 => x"fe824449",
			4333 => x"07002904",
			4334 => x"005d4449",
			4335 => x"ff294449",
			4336 => x"06005e04",
			4337 => x"ff144449",
			4338 => x"06006504",
			4339 => x"01734449",
			4340 => x"00624449",
			4341 => x"0d001304",
			4342 => x"ffeb4449",
			4343 => x"fe7e4449",
			4344 => x"0000dd14",
			4345 => x"0d001808",
			4346 => x"04002d04",
			4347 => x"ffa64449",
			4348 => x"01924449",
			4349 => x"01000b04",
			4350 => x"00a44449",
			4351 => x"07003204",
			4352 => x"ff0f4449",
			4353 => x"00004449",
			4354 => x"0e006804",
			4355 => x"fe8b4449",
			4356 => x"0d001504",
			4357 => x"013e4449",
			4358 => x"0200d604",
			4359 => x"ff654449",
			4360 => x"03006504",
			4361 => x"00ae4449",
			4362 => x"ffbf4449",
			4363 => x"03003d04",
			4364 => x"fe8f4449",
			4365 => x"01001008",
			4366 => x"0f008e04",
			4367 => x"ffa24449",
			4368 => x"01154449",
			4369 => x"ff214449",
			4370 => x"0d001538",
			4371 => x"03003928",
			4372 => x"07002508",
			4373 => x"05003e04",
			4374 => x"ffdb452d",
			4375 => x"0075452d",
			4376 => x"0700280c",
			4377 => x"09001d08",
			4378 => x"0d001204",
			4379 => x"fffb452d",
			4380 => x"0033452d",
			4381 => x"ff45452d",
			4382 => x"0000df10",
			4383 => x"01000908",
			4384 => x"0b001904",
			4385 => x"009c452d",
			4386 => x"fff3452d",
			4387 => x"0000b504",
			4388 => x"ffa5452d",
			4389 => x"0025452d",
			4390 => x"ffaa452d",
			4391 => x"04003c04",
			4392 => x"00a9452d",
			4393 => x"08001b08",
			4394 => x"09002004",
			4395 => x"0002452d",
			4396 => x"0082452d",
			4397 => x"ffb0452d",
			4398 => x"0b001914",
			4399 => x"0b001608",
			4400 => x"06006f04",
			4401 => x"0017452d",
			4402 => x"fff1452d",
			4403 => x"04002f08",
			4404 => x"0a003604",
			4405 => x"fff7452d",
			4406 => x"0015452d",
			4407 => x"ff41452d",
			4408 => x"0a003b04",
			4409 => x"ff95452d",
			4410 => x"04004614",
			4411 => x"01000e08",
			4412 => x"05005304",
			4413 => x"00b5452d",
			4414 => x"0012452d",
			4415 => x"06007004",
			4416 => x"ffda452d",
			4417 => x"0600a104",
			4418 => x"000c452d",
			4419 => x"fff4452d",
			4420 => x"0f007204",
			4421 => x"ffac452d",
			4422 => x"0e006804",
			4423 => x"003d452d",
			4424 => x"0e007104",
			4425 => x"ffc9452d",
			4426 => x"001d452d",
			4427 => x"0e006530",
			4428 => x"0200b924",
			4429 => x"0e005c20",
			4430 => x"08001d14",
			4431 => x"0c001a0c",
			4432 => x"03003908",
			4433 => x"09001d04",
			4434 => x"012d4601",
			4435 => x"ff0f4601",
			4436 => x"00db4601",
			4437 => x"0000a204",
			4438 => x"ff134601",
			4439 => x"01494601",
			4440 => x"09001e08",
			4441 => x"0c001704",
			4442 => x"ffdc4601",
			4443 => x"00b74601",
			4444 => x"fea64601",
			4445 => x"fed54601",
			4446 => x"0f006c04",
			4447 => x"ff034601",
			4448 => x"0200d004",
			4449 => x"016b4601",
			4450 => x"ffc74601",
			4451 => x"0100040c",
			4452 => x"0000e504",
			4453 => x"fe724601",
			4454 => x"00012804",
			4455 => x"00104601",
			4456 => x"ffd94601",
			4457 => x"03003e18",
			4458 => x"08001b14",
			4459 => x"0000e108",
			4460 => x"05002504",
			4461 => x"ffe94601",
			4462 => x"012f4601",
			4463 => x"07002b04",
			4464 => x"feb74601",
			4465 => x"07002c04",
			4466 => x"00494601",
			4467 => x"ffa34601",
			4468 => x"fe9f4601",
			4469 => x"06007004",
			4470 => x"ff444601",
			4471 => x"01000b04",
			4472 => x"014c4601",
			4473 => x"0f008508",
			4474 => x"06007204",
			4475 => x"00414601",
			4476 => x"ff394601",
			4477 => x"01001004",
			4478 => x"00e04601",
			4479 => x"ff6e4601",
			4480 => x"05003c04",
			4481 => x"fe66467d",
			4482 => x"08002334",
			4483 => x"07002508",
			4484 => x"03003304",
			4485 => x"01d8467d",
			4486 => x"0134467d",
			4487 => x"05004910",
			4488 => x"0d001304",
			4489 => x"fe83467d",
			4490 => x"0a003704",
			4491 => x"fed3467d",
			4492 => x"0d001504",
			4493 => x"0143467d",
			4494 => x"ffdb467d",
			4495 => x"0d00140c",
			4496 => x"09001f04",
			4497 => x"022b467d",
			4498 => x"08001b04",
			4499 => x"0179467d",
			4500 => x"0072467d",
			4501 => x"0b001908",
			4502 => x"08001b04",
			4503 => x"0094467d",
			4504 => x"fe8b467d",
			4505 => x"03005c04",
			4506 => x"0114467d",
			4507 => x"fe9a467d",
			4508 => x"01001004",
			4509 => x"ff60467d",
			4510 => x"fe77467d",
			4511 => x"05003c04",
			4512 => x"fe6b4709",
			4513 => x"0200e734",
			4514 => x"09001d04",
			4515 => x"01d74709",
			4516 => x"0000b414",
			4517 => x"04003b0c",
			4518 => x"0e005508",
			4519 => x"06005704",
			4520 => x"fea44709",
			4521 => x"00464709",
			4522 => x"fe344709",
			4523 => x"09002104",
			4524 => x"01334709",
			4525 => x"fe6f4709",
			4526 => x"04003c0c",
			4527 => x"0d001508",
			4528 => x"07002904",
			4529 => x"01044709",
			4530 => x"01d34709",
			4531 => x"ffd84709",
			4532 => x"06006b08",
			4533 => x"09002604",
			4534 => x"01544709",
			4535 => x"feec4709",
			4536 => x"0000d004",
			4537 => x"fe6a4709",
			4538 => x"00c74709",
			4539 => x"05005008",
			4540 => x"03003d04",
			4541 => x"fe464709",
			4542 => x"001a4709",
			4543 => x"0d001b04",
			4544 => x"01584709",
			4545 => x"fec74709",
			4546 => x"0000ed68",
			4547 => x"01000938",
			4548 => x"01000830",
			4549 => x"08001b1c",
			4550 => x"0700270c",
			4551 => x"07002508",
			4552 => x"05003704",
			4553 => x"ffeb47f7",
			4554 => x"003447f7",
			4555 => x"ffac47f7",
			4556 => x"0d001208",
			4557 => x"0f008804",
			4558 => x"001047f7",
			4559 => x"ffd947f7",
			4560 => x"06005904",
			4561 => x"fff547f7",
			4562 => x"00ce47f7",
			4563 => x"0d00140c",
			4564 => x"0000a608",
			4565 => x"0c001804",
			4566 => x"000b47f7",
			4567 => x"ffc047f7",
			4568 => x"005147f7",
			4569 => x"0c001b04",
			4570 => x"ff7347f7",
			4571 => x"000447f7",
			4572 => x"0a003b04",
			4573 => x"000f47f7",
			4574 => x"00bc47f7",
			4575 => x"0200b918",
			4576 => x"0e005a14",
			4577 => x"08001c08",
			4578 => x"05003f04",
			4579 => x"fff047f7",
			4580 => x"007647f7",
			4581 => x"0200a808",
			4582 => x"09001e04",
			4583 => x"000847f7",
			4584 => x"ffb347f7",
			4585 => x"001247f7",
			4586 => x"ff5747f7",
			4587 => x"04004c10",
			4588 => x"08001f08",
			4589 => x"04003404",
			4590 => x"fff947f7",
			4591 => x"008747f7",
			4592 => x"07003004",
			4593 => x"ffe247f7",
			4594 => x"000b47f7",
			4595 => x"0e006d04",
			4596 => x"ffcd47f7",
			4597 => x"001c47f7",
			4598 => x"05005008",
			4599 => x"03003d04",
			4600 => x"ff8447f7",
			4601 => x"000447f7",
			4602 => x"03005304",
			4603 => x"002c47f7",
			4604 => x"ffdf47f7",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1473, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2995, initial_addr_3'length));
	end generate gen_rom_8;

	gen_rom_9: if SELECT_ROM = 9 generate
		bank <= (
			0 => x"0f005814",
			1 => x"02006b0c",
			2 => x"03001a08",
			3 => x"02004604",
			4 => x"ffe8004d",
			5 => x"0038004d",
			6 => x"ffcc004d",
			7 => x"03002d04",
			8 => x"0071004d",
			9 => x"ffec004d",
			10 => x"0200bb08",
			11 => x"0200b904",
			12 => x"ffaa004d",
			13 => x"ffff004d",
			14 => x"0200f308",
			15 => x"04005004",
			16 => x"0049004d",
			17 => x"fff7004d",
			18 => x"ffe0004d",
			19 => x"05002118",
			20 => x"0f005610",
			21 => x"02004604",
			22 => x"ffe600a9",
			23 => x"08002008",
			24 => x"03001f04",
			25 => x"007100a9",
			26 => x"000400a9",
			27 => x"fffb00a9",
			28 => x"0000a404",
			29 => x"ffe100a9",
			30 => x"000500a9",
			31 => x"0000a90c",
			32 => x"04001804",
			33 => x"000600a9",
			34 => x"0c001e04",
			35 => x"ffa200a9",
			36 => x"000200a9",
			37 => x"0f006c04",
			38 => x"005200a9",
			39 => x"07002704",
			40 => x"000900a9",
			41 => x"ffc100a9",
			42 => x"0f00501c",
			43 => x"02006b14",
			44 => x"03001a10",
			45 => x"01000708",
			46 => x"02003a04",
			47 => x"fff60105",
			48 => x"00410105",
			49 => x"04000704",
			50 => x"000c0105",
			51 => x"ffd40105",
			52 => x"ffc90105",
			53 => x"03002304",
			54 => x"00710105",
			55 => x"fffd0105",
			56 => x"0200b908",
			57 => x"0a001c04",
			58 => x"00040105",
			59 => x"ff910105",
			60 => x"0f007308",
			61 => x"04006104",
			62 => x"00630105",
			63 => x"fff60105",
			64 => x"ffd10105",
			65 => x"0f006624",
			66 => x"02006b10",
			67 => x"03001a0c",
			68 => x"09001504",
			69 => x"ffd60169",
			70 => x"00004804",
			71 => x"ffec0169",
			72 => x"00510169",
			73 => x"ffb40169",
			74 => x"0f005008",
			75 => x"03002304",
			76 => x"00970169",
			77 => x"00030169",
			78 => x"0200a108",
			79 => x"0b001804",
			80 => x"ffa00169",
			81 => x"fffa0169",
			82 => x"006f0169",
			83 => x"0b002308",
			84 => x"08001504",
			85 => x"001b0169",
			86 => x"ff870169",
			87 => x"09003004",
			88 => x"002b0169",
			89 => x"fffb0169",
			90 => x"06006820",
			91 => x"02004604",
			92 => x"ffe601b5",
			93 => x"05003f08",
			94 => x"0d002004",
			95 => x"005c01b5",
			96 => x"fff801b5",
			97 => x"04003608",
			98 => x"03003904",
			99 => x"ffe001b5",
			100 => x"000201b5",
			101 => x"0a003b04",
			102 => x"fff301b5",
			103 => x"04005104",
			104 => x"002b01b5",
			105 => x"fff901b5",
			106 => x"0d002504",
			107 => x"ffd301b5",
			108 => x"000801b5",
			109 => x"0f00662c",
			110 => x"02008018",
			111 => x"06003e10",
			112 => x"02005908",
			113 => x"0b001104",
			114 => x"00140231",
			115 => x"ffc20231",
			116 => x"03002104",
			117 => x"00790231",
			118 => x"ffe30231",
			119 => x"01001004",
			120 => x"ff8f0231",
			121 => x"00040231",
			122 => x"0500480c",
			123 => x"0b001b04",
			124 => x"00800231",
			125 => x"03002d04",
			126 => x"00100231",
			127 => x"fff10231",
			128 => x"09002104",
			129 => x"ffe70231",
			130 => x"000c0231",
			131 => x"0c002008",
			132 => x"01000304",
			133 => x"000c0231",
			134 => x"ff8d0231",
			135 => x"07003908",
			136 => x"0200d504",
			137 => x"fff90231",
			138 => x"00390231",
			139 => x"fff50231",
			140 => x"0600682c",
			141 => x"0200991c",
			142 => x"0f00420c",
			143 => x"02004604",
			144 => x"ffe00295",
			145 => x"03002104",
			146 => x"006a0295",
			147 => x"ffe20295",
			148 => x"0b001808",
			149 => x"01001004",
			150 => x"ffa60295",
			151 => x"00090295",
			152 => x"0a002f04",
			153 => x"00300295",
			154 => x"ffda0295",
			155 => x"05004804",
			156 => x"00620295",
			157 => x"05005304",
			158 => x"ffeb0295",
			159 => x"04005104",
			160 => x"001a0295",
			161 => x"fffa0295",
			162 => x"0d002504",
			163 => x"ffc60295",
			164 => x"000a0295",
			165 => x"0f007328",
			166 => x"02009c1c",
			167 => x"0f004b14",
			168 => x"0300230c",
			169 => x"02004604",
			170 => x"ffc402e9",
			171 => x"03001f04",
			172 => x"00ac02e9",
			173 => x"001d02e9",
			174 => x"07002404",
			175 => x"ffb002e9",
			176 => x"000b02e9",
			177 => x"05001b04",
			178 => x"fffa02e9",
			179 => x"ff6802e9",
			180 => x"05004804",
			181 => x"00b002e9",
			182 => x"0200d004",
			183 => x"ffaa02e9",
			184 => x"004902e9",
			185 => x"ff8202e9",
			186 => x"0f006628",
			187 => x"00008314",
			188 => x"0f004010",
			189 => x"06002804",
			190 => x"ffea0355",
			191 => x"09001b04",
			192 => x"00440355",
			193 => x"03001704",
			194 => x"00080355",
			195 => x"fff10355",
			196 => x"ffb20355",
			197 => x"0d001e10",
			198 => x"0f006108",
			199 => x"05004804",
			200 => x"00560355",
			201 => x"00010355",
			202 => x"0f006404",
			203 => x"fff90355",
			204 => x"00060355",
			205 => x"fffe0355",
			206 => x"0d001004",
			207 => x"000f0355",
			208 => x"0c002004",
			209 => x"ffbe0355",
			210 => x"07003904",
			211 => x"00110355",
			212 => x"fffa0355",
			213 => x"0f00732c",
			214 => x"0200991c",
			215 => x"0f00420c",
			216 => x"03002108",
			217 => x"02004604",
			218 => x"ffe203b1",
			219 => x"006d03b1",
			220 => x"ffdf03b1",
			221 => x"0b001808",
			222 => x"01001004",
			223 => x"ffa203b1",
			224 => x"000803b1",
			225 => x"0a002f04",
			226 => x"003003b1",
			227 => x"ffd903b1",
			228 => x"05004804",
			229 => x"006403b1",
			230 => x"0a004704",
			231 => x"ffe603b1",
			232 => x"04005104",
			233 => x"002003b1",
			234 => x"fff803b1",
			235 => x"ffcc03b1",
			236 => x"08001508",
			237 => x"0d001004",
			238 => x"00570425",
			239 => x"fff20425",
			240 => x"0b00181c",
			241 => x"0f00400c",
			242 => x"0f003608",
			243 => x"05000c04",
			244 => x"ffff0425",
			245 => x"ffd50425",
			246 => x"00340425",
			247 => x"01000304",
			248 => x"00040425",
			249 => x"04003c04",
			250 => x"ff760425",
			251 => x"04003e04",
			252 => x"000a0425",
			253 => x"fff90425",
			254 => x"02008b08",
			255 => x"07001f04",
			256 => x"00020425",
			257 => x"ffd60425",
			258 => x"0f006c08",
			259 => x"0a006504",
			260 => x"00670425",
			261 => x"fff90425",
			262 => x"0d002504",
			263 => x"ffda0425",
			264 => x"000b0425",
			265 => x"06006730",
			266 => x"02006b10",
			267 => x"0600370c",
			268 => x"02004604",
			269 => x"ffc10491",
			270 => x"0a001e04",
			271 => x"008c0491",
			272 => x"ffd70491",
			273 => x"ff890491",
			274 => x"0f005008",
			275 => x"05002d04",
			276 => x"00ba0491",
			277 => x"fff60491",
			278 => x"0200a10c",
			279 => x"0d001404",
			280 => x"ff6f0491",
			281 => x"04001f04",
			282 => x"00360491",
			283 => x"ffba0491",
			284 => x"05004804",
			285 => x"00910491",
			286 => x"0000cb04",
			287 => x"ffc30491",
			288 => x"003f0491",
			289 => x"0d002504",
			290 => x"ff710491",
			291 => x"00140491",
			292 => x"06006734",
			293 => x"02008220",
			294 => x"0f004218",
			295 => x"0c00180c",
			296 => x"02004604",
			297 => x"ffd60505",
			298 => x"0d001304",
			299 => x"00bc0505",
			300 => x"fffe0505",
			301 => x"04000d08",
			302 => x"07002304",
			303 => x"00120505",
			304 => x"fff70505",
			305 => x"ffb00505",
			306 => x"01001004",
			307 => x"ff720505",
			308 => x"00040505",
			309 => x"05004508",
			310 => x"0f006604",
			311 => x"00b40505",
			312 => x"00120505",
			313 => x"0b001d08",
			314 => x"0f005c04",
			315 => x"fffc0505",
			316 => x"ff980505",
			317 => x"003c0505",
			318 => x"0d002504",
			319 => x"ff6b0505",
			320 => x"00140505",
			321 => x"08001508",
			322 => x"0d001004",
			323 => x"00550581",
			324 => x"fff20581",
			325 => x"0b00181c",
			326 => x"0f00400c",
			327 => x"0f003608",
			328 => x"05000c04",
			329 => x"ffff0581",
			330 => x"ffd60581",
			331 => x"00340581",
			332 => x"01000304",
			333 => x"00040581",
			334 => x"04003c04",
			335 => x"ff7c0581",
			336 => x"04003e04",
			337 => x"000a0581",
			338 => x"fff90581",
			339 => x"02008b0c",
			340 => x"07002308",
			341 => x"07001f04",
			342 => x"00020581",
			343 => x"ffff0581",
			344 => x"ffd70581",
			345 => x"0f006c08",
			346 => x"0a006504",
			347 => x"00640581",
			348 => x"fff90581",
			349 => x"0d002504",
			350 => x"ffdb0581",
			351 => x"000b0581",
			352 => x"0f006e30",
			353 => x"0200a124",
			354 => x"05002d1c",
			355 => x"02006b10",
			356 => x"0600370c",
			357 => x"02004604",
			358 => x"ff8205f5",
			359 => x"0a001c04",
			360 => x"00ea05f5",
			361 => x"ffb105f5",
			362 => x"ff0905f5",
			363 => x"0f005408",
			364 => x"01000904",
			365 => x"013105f5",
			366 => x"004a05f5",
			367 => x"ffb105f5",
			368 => x"04002204",
			369 => x"ffef05f5",
			370 => x"fef105f5",
			371 => x"0f006604",
			372 => x"012605f5",
			373 => x"0200d204",
			374 => x"ff5005f5",
			375 => x"00c605f5",
			376 => x"0d002504",
			377 => x"fee505f5",
			378 => x"04002e04",
			379 => x"fffa05f5",
			380 => x"003805f5",
			381 => x"0f007330",
			382 => x"00007514",
			383 => x"0f004010",
			384 => x"02004604",
			385 => x"ff970659",
			386 => x"09001b04",
			387 => x"00dd0659",
			388 => x"07002204",
			389 => x"ffc90659",
			390 => x"fffe0659",
			391 => x"ff240659",
			392 => x"06004c08",
			393 => x"05002e04",
			394 => x"010f0659",
			395 => x"00030659",
			396 => x"0200a508",
			397 => x"04001804",
			398 => x"00140659",
			399 => x"ff290659",
			400 => x"05004804",
			401 => x"00e00659",
			402 => x"0200d004",
			403 => x"ff870659",
			404 => x"006f0659",
			405 => x"ff330659",
			406 => x"06006834",
			407 => x"02008220",
			408 => x"06003f18",
			409 => x"0c00180c",
			410 => x"02004604",
			411 => x"ffe106cd",
			412 => x"0d001304",
			413 => x"009006cd",
			414 => x"000006cd",
			415 => x"05001208",
			416 => x"07002204",
			417 => x"000a06cd",
			418 => x"fff906cd",
			419 => x"ffca06cd",
			420 => x"01001004",
			421 => x"ff9306cd",
			422 => x"fffd06cd",
			423 => x"05004504",
			424 => x"008f06cd",
			425 => x"0200bc0c",
			426 => x"07002708",
			427 => x"07002604",
			428 => x"fff706cd",
			429 => x"000606cd",
			430 => x"ffb406cd",
			431 => x"004206cd",
			432 => x"0d002504",
			433 => x"ff9f06cd",
			434 => x"000e06cd",
			435 => x"0f007334",
			436 => x"02006b0c",
			437 => x"08001604",
			438 => x"00c60739",
			439 => x"04000704",
			440 => x"00400739",
			441 => x"fe760739",
			442 => x"05003214",
			443 => x"0600510c",
			444 => x"02008008",
			445 => x"07001f04",
			446 => x"01300739",
			447 => x"007b0739",
			448 => x"01830739",
			449 => x"0000af04",
			450 => x"ff0b0739",
			451 => x"01290739",
			452 => x"0200ca0c",
			453 => x"0f005808",
			454 => x"00008b04",
			455 => x"ff0d0739",
			456 => x"00780739",
			457 => x"fe9b0739",
			458 => x"04006104",
			459 => x"01660739",
			460 => x"ff730739",
			461 => x"fe840739",
			462 => x"0f007334",
			463 => x"02007114",
			464 => x"0f004010",
			465 => x"02004604",
			466 => x"ff9c07a5",
			467 => x"09001b04",
			468 => x"00d807a5",
			469 => x"07002204",
			470 => x"ffcd07a5",
			471 => x"ffff07a5",
			472 => x"ff3407a5",
			473 => x"06004c0c",
			474 => x"05002e08",
			475 => x"08002004",
			476 => x"010c07a5",
			477 => x"001207a5",
			478 => x"000c07a5",
			479 => x"0200a108",
			480 => x"04001804",
			481 => x"000407a5",
			482 => x"ff3907a5",
			483 => x"0f006604",
			484 => x"00ec07a5",
			485 => x"0200d504",
			486 => x"ff6907a5",
			487 => x"00a807a5",
			488 => x"ff3c07a5",
			489 => x"0600682c",
			490 => x"0200b928",
			491 => x"0600501c",
			492 => x"02006b10",
			493 => x"0600370c",
			494 => x"02004604",
			495 => x"ffc80809",
			496 => x"0a001e04",
			497 => x"00780809",
			498 => x"ffdc0809",
			499 => x"ff8e0809",
			500 => x"04002208",
			501 => x"08002004",
			502 => x"00ba0809",
			503 => x"fff80809",
			504 => x"ffda0809",
			505 => x"0200ac04",
			506 => x"ff760809",
			507 => x"0d001304",
			508 => x"002f0809",
			509 => x"ffde0809",
			510 => x"009e0809",
			511 => x"0d002504",
			512 => x"ff870809",
			513 => x"00110809",
			514 => x"0f007324",
			515 => x"02005004",
			516 => x"fe6d0855",
			517 => x"0700391c",
			518 => x"0000c614",
			519 => x"06005a0c",
			520 => x"0a001b04",
			521 => x"01b20855",
			522 => x"00008304",
			523 => x"feeb0855",
			524 => x"01350855",
			525 => x"0200b904",
			526 => x"fe690855",
			527 => x"ffdc0855",
			528 => x"04006104",
			529 => x"01d20855",
			530 => x"feab0855",
			531 => x"fe810855",
			532 => x"fe670855",
			533 => x"0f007330",
			534 => x"0200bb28",
			535 => x"0f00551c",
			536 => x"00007510",
			537 => x"0f003c0c",
			538 => x"02004604",
			539 => x"ffd508b9",
			540 => x"09001b04",
			541 => x"006808b9",
			542 => x"ffea08b9",
			543 => x"ff9908b9",
			544 => x"03002d08",
			545 => x"08002004",
			546 => x"008e08b9",
			547 => x"fffd08b9",
			548 => x"ffdc08b9",
			549 => x"0200ac04",
			550 => x"ff9408b9",
			551 => x"0000b904",
			552 => x"000408b9",
			553 => x"fff708b9",
			554 => x"04006104",
			555 => x"008708b9",
			556 => x"fff308b9",
			557 => x"ffb308b9",
			558 => x"01000518",
			559 => x"0400140c",
			560 => x"0a001608",
			561 => x"0f001e04",
			562 => x"fffb094d",
			563 => x"0036094d",
			564 => x"ffaa094d",
			565 => x"0d001308",
			566 => x"07002704",
			567 => x"00a9094d",
			568 => x"fff1094d",
			569 => x"ffe3094d",
			570 => x"08001504",
			571 => x"004d094d",
			572 => x"0b001814",
			573 => x"05000f08",
			574 => x"0f002404",
			575 => x"fff7094d",
			576 => x"0029094d",
			577 => x"04003c04",
			578 => x"ff4b094d",
			579 => x"04003f04",
			580 => x"0013094d",
			581 => x"fff9094d",
			582 => x"0a002f0c",
			583 => x"00007804",
			584 => x"ffd9094d",
			585 => x"07003004",
			586 => x"0082094d",
			587 => x"fff9094d",
			588 => x"0200c404",
			589 => x"ff9e094d",
			590 => x"06006c08",
			591 => x"03005c04",
			592 => x"005c094d",
			593 => x"fff3094d",
			594 => x"ffdb094d",
			595 => x"0f007338",
			596 => x"02009c24",
			597 => x"0f004b18",
			598 => x"02004604",
			599 => x"fec709c1",
			600 => x"0300220c",
			601 => x"03001a04",
			602 => x"017a09c1",
			603 => x"0a002004",
			604 => x"ff5c09c1",
			605 => x"011b09c1",
			606 => x"07002404",
			607 => x"fed909c1",
			608 => x"006409c1",
			609 => x"00008304",
			610 => x"fe6209c1",
			611 => x"0f005404",
			612 => x"00ed09c1",
			613 => x"feac09c1",
			614 => x"0f006104",
			615 => x"017a09c1",
			616 => x"0000cc08",
			617 => x"0200ba04",
			618 => x"feab09c1",
			619 => x"ff9b09c1",
			620 => x"04006104",
			621 => x"017609c1",
			622 => x"ff4609c1",
			623 => x"fe7e09c1",
			624 => x"06006834",
			625 => x"02005008",
			626 => x"0d001004",
			627 => x"fffe0a3d",
			628 => x"fe5b0a3d",
			629 => x"05004824",
			630 => x"0200a518",
			631 => x"06004e10",
			632 => x"05002d08",
			633 => x"02006b04",
			634 => x"01160a3d",
			635 => x"02b00a3d",
			636 => x"04002504",
			637 => x"00ac0a3d",
			638 => x"fe510a3d",
			639 => x"05001f04",
			640 => x"00410a3d",
			641 => x"fe500a3d",
			642 => x"0d001304",
			643 => x"02f60a3d",
			644 => x"09002004",
			645 => x"02120a3d",
			646 => x"02780a3d",
			647 => x"01001004",
			648 => x"fe560a3d",
			649 => x"01d20a3d",
			650 => x"0f007308",
			651 => x"05006304",
			652 => x"01090a3d",
			653 => x"fe6b0a3d",
			654 => x"fe590a3d",
			655 => x"0f007334",
			656 => x"02006b0c",
			657 => x"08001604",
			658 => x"00b80aa9",
			659 => x"04000704",
			660 => x"00d60aa9",
			661 => x"fe460aa9",
			662 => x"05004820",
			663 => x"0000a918",
			664 => x"06004c0c",
			665 => x"05002d08",
			666 => x"01000904",
			667 => x"01cb0aa9",
			668 => x"01150aa9",
			669 => x"000e0aa9",
			670 => x"02008e04",
			671 => x"fe740aa9",
			672 => x"0e004e04",
			673 => x"01070aa9",
			674 => x"fe970aa9",
			675 => x"0f006604",
			676 => x"01b80aa9",
			677 => x"00ba0aa9",
			678 => x"0000df04",
			679 => x"fe770aa9",
			680 => x"01b10aa9",
			681 => x"fe6b0aa9",
			682 => x"0600673c",
			683 => x"02005008",
			684 => x"0d001004",
			685 => x"000c0b35",
			686 => x"fe580b35",
			687 => x"05004024",
			688 => x"02008b10",
			689 => x"05001b08",
			690 => x"06003e04",
			691 => x"02d40b35",
			692 => x"01880b35",
			693 => x"01000704",
			694 => x"01040b35",
			695 => x"fe4f0b35",
			696 => x"0600590c",
			697 => x"0f005a08",
			698 => x"01000c04",
			699 => x"03010b35",
			700 => x"02a70b35",
			701 => x"02660b35",
			702 => x"0000ba04",
			703 => x"fe470b35",
			704 => x"03030b35",
			705 => x"0000c60c",
			706 => x"01000608",
			707 => x"06005d04",
			708 => x"00bd0b35",
			709 => x"fe630b35",
			710 => x"fe580b35",
			711 => x"030d0b35",
			712 => x"0d002504",
			713 => x"fe570b35",
			714 => x"0600b204",
			715 => x"00750b35",
			716 => x"fe680b35",
			717 => x"0f007328",
			718 => x"02005004",
			719 => x"fe8e0b89",
			720 => x"0a001604",
			721 => x"01940b89",
			722 => x"0200bb14",
			723 => x"0f006110",
			724 => x"02009808",
			725 => x"0f005004",
			726 => x"00870b89",
			727 => x"fe9f0b89",
			728 => x"0f005804",
			729 => x"01970b89",
			730 => x"00ea0b89",
			731 => x"fe880b89",
			732 => x"03005c08",
			733 => x"0000cc04",
			734 => x"00ee0b89",
			735 => x"019c0b89",
			736 => x"feef0b89",
			737 => x"fe700b89",
			738 => x"0f00733c",
			739 => x"02006b10",
			740 => x"0b001208",
			741 => x"0c001104",
			742 => x"ffb80c05",
			743 => x"01070c05",
			744 => x"04000504",
			745 => x"00320c05",
			746 => x"fea60c05",
			747 => x"01000508",
			748 => x"0f006104",
			749 => x"01620c05",
			750 => x"00290c05",
			751 => x"0b001810",
			752 => x"05001b04",
			753 => x"00dc0c05",
			754 => x"02009c04",
			755 => x"fec30c05",
			756 => x"06005f04",
			757 => x"00d70c05",
			758 => x"ff610c05",
			759 => x"0a002f08",
			760 => x"0e004f04",
			761 => x"01510c05",
			762 => x"00280c05",
			763 => x"0200c404",
			764 => x"fef90c05",
			765 => x"04006104",
			766 => x"01360c05",
			767 => x"ff9e0c05",
			768 => x"fea70c05",
			769 => x"0f006e3c",
			770 => x"02004604",
			771 => x"fe600c91",
			772 => x"05002f20",
			773 => x"0000750c",
			774 => x"03001a04",
			775 => x"01df0c91",
			776 => x"04001f04",
			777 => x"fe540c91",
			778 => x"ffff0c91",
			779 => x"0f00580c",
			780 => x"08001b04",
			781 => x"025b0c91",
			782 => x"0b001804",
			783 => x"01990c91",
			784 => x"021b0c91",
			785 => x"0000af04",
			786 => x"fe4d0c91",
			787 => x"021f0c91",
			788 => x"0200bc0c",
			789 => x"0000a904",
			790 => x"fe560c91",
			791 => x"0f006704",
			792 => x"018b0c91",
			793 => x"fe660c91",
			794 => x"03006108",
			795 => x"04003104",
			796 => x"020e0c91",
			797 => x"02c30c91",
			798 => x"fe4c0c91",
			799 => x"0d002504",
			800 => x"fe5e0c91",
			801 => x"0d002704",
			802 => x"01020c91",
			803 => x"fe7c0c91",
			804 => x"0f007348",
			805 => x"02008224",
			806 => x"06003e1c",
			807 => x"0c00180c",
			808 => x"02004604",
			809 => x"ff8d0d25",
			810 => x"05002304",
			811 => x"01360d25",
			812 => x"ffb40d25",
			813 => x"04000d0c",
			814 => x"07002208",
			815 => x"07001d04",
			816 => x"fff70d25",
			817 => x"00490d25",
			818 => x"ffd00d25",
			819 => x"ff2f0d25",
			820 => x"01001004",
			821 => x"fee70d25",
			822 => x"00180d25",
			823 => x"0f006114",
			824 => x"05004810",
			825 => x"0b001508",
			826 => x"02008f04",
			827 => x"ff990d25",
			828 => x"007e0d25",
			829 => x"01001004",
			830 => x"014f0d25",
			831 => x"00160d25",
			832 => x"ffc40d25",
			833 => x"0000cc08",
			834 => x"01000e04",
			835 => x"fee30d25",
			836 => x"ffe90d25",
			837 => x"04006104",
			838 => x"012b0d25",
			839 => x"ffb00d25",
			840 => x"feb70d25",
			841 => x"0f007330",
			842 => x"02005004",
			843 => x"fe690d89",
			844 => x"05004824",
			845 => x"0200a518",
			846 => x"0f005510",
			847 => x"05002c08",
			848 => x"00007504",
			849 => x"005c0d89",
			850 => x"01dc0d89",
			851 => x"04002204",
			852 => x"00a40d89",
			853 => x"fe6f0d89",
			854 => x"08001d04",
			855 => x"fe5a0d89",
			856 => x"ff2e0d89",
			857 => x"0f006608",
			858 => x"01000604",
			859 => x"021c0d89",
			860 => x"01b80d89",
			861 => x"012d0d89",
			862 => x"01001104",
			863 => x"fe670d89",
			864 => x"01ee0d89",
			865 => x"fe640d89",
			866 => x"0f00732c",
			867 => x"02005004",
			868 => x"fe630de5",
			869 => x"0200d924",
			870 => x"06005e18",
			871 => x"02009810",
			872 => x"0a001b08",
			873 => x"08001c04",
			874 => x"02030de5",
			875 => x"01ab0de5",
			876 => x"00008304",
			877 => x"feab0de5",
			878 => x"00790de5",
			879 => x"05004804",
			880 => x"01f00de5",
			881 => x"ffa60de5",
			882 => x"0000cc04",
			883 => x"fe580de5",
			884 => x"04009004",
			885 => x"00cc0de5",
			886 => x"fe700de5",
			887 => x"02900de5",
			888 => x"fe600de5",
			889 => x"0f007334",
			890 => x"02004604",
			891 => x"fe6d0e51",
			892 => x"0200bb24",
			893 => x"0f005818",
			894 => x"00008b0c",
			895 => x"03002108",
			896 => x"0f004304",
			897 => x"01c30e51",
			898 => x"ff4e0e51",
			899 => x"fe6a0e51",
			900 => x"0b001b08",
			901 => x"0c001804",
			902 => x"01460e51",
			903 => x"01ee0e51",
			904 => x"01620e51",
			905 => x"0200a704",
			906 => x"fe640e51",
			907 => x"03003a04",
			908 => x"015f0e51",
			909 => x"fe800e51",
			910 => x"04006108",
			911 => x"0200d904",
			912 => x"01a10e51",
			913 => x"020c0e51",
			914 => x"fe970e51",
			915 => x"fe660e51",
			916 => x"0f00733c",
			917 => x"0000c634",
			918 => x"0f005828",
			919 => x"02007118",
			920 => x"0100070c",
			921 => x"03001a08",
			922 => x"00004304",
			923 => x"ffa40ecd",
			924 => x"01520ecd",
			925 => x"ffe60ecd",
			926 => x"04000704",
			927 => x"00580ecd",
			928 => x"0a000b04",
			929 => x"fff90ecd",
			930 => x"febc0ecd",
			931 => x"0500360c",
			932 => x"08002008",
			933 => x"0b001504",
			934 => x"00a10ecd",
			935 => x"017b0ecd",
			936 => x"004f0ecd",
			937 => x"ffe90ecd",
			938 => x"0200b304",
			939 => x"feb00ecd",
			940 => x"0000c304",
			941 => x"fffa0ecd",
			942 => x"ffd80ecd",
			943 => x"04006104",
			944 => x"015a0ecd",
			945 => x"ff8f0ecd",
			946 => x"fe9a0ecd",
			947 => x"0f007330",
			948 => x"02004604",
			949 => x"fe650f31",
			950 => x"0a006528",
			951 => x"0000c51c",
			952 => x"05003210",
			953 => x"0f005408",
			954 => x"02006b04",
			955 => x"00370f31",
			956 => x"01ec0f31",
			957 => x"02009004",
			958 => x"fe4a0f31",
			959 => x"01480f31",
			960 => x"0200a504",
			961 => x"fe5c0f31",
			962 => x"05004904",
			963 => x"011c0f31",
			964 => x"fe6f0f31",
			965 => x"0000e608",
			966 => x"0e005a04",
			967 => x"01f40f31",
			968 => x"01010f31",
			969 => x"02890f31",
			970 => x"fe630f31",
			971 => x"fe610f31",
			972 => x"0f00733c",
			973 => x"08001504",
			974 => x"017c0fad",
			975 => x"00008b10",
			976 => x"06003d0c",
			977 => x"02005c08",
			978 => x"05000a04",
			979 => x"00640fad",
			980 => x"fe9b0fad",
			981 => x"01450fad",
			982 => x"fe4c0fad",
			983 => x"06005a14",
			984 => x"05004810",
			985 => x"0b001608",
			986 => x"00009904",
			987 => x"ff7a0fad",
			988 => x"00d60fad",
			989 => x"01001104",
			990 => x"01920fad",
			991 => x"00340fad",
			992 => x"ff920fad",
			993 => x"0200cf0c",
			994 => x"0200ba04",
			995 => x"fe8b0fad",
			996 => x"04004304",
			997 => x"007a0fad",
			998 => x"ff090fad",
			999 => x"04006104",
			1000 => x"01860fad",
			1001 => x"ff550fad",
			1002 => x"fe760fad",
			1003 => x"0f007340",
			1004 => x"0d000e04",
			1005 => x"01ae1031",
			1006 => x"02006b10",
			1007 => x"03000c08",
			1008 => x"00002c04",
			1009 => x"ff851031",
			1010 => x"010d1031",
			1011 => x"08001804",
			1012 => x"ff461031",
			1013 => x"fe211031",
			1014 => x"0f005514",
			1015 => x"00008b0c",
			1016 => x"06004608",
			1017 => x"01000904",
			1018 => x"01ac1031",
			1019 => x"ffe01031",
			1020 => x"fe971031",
			1021 => x"0b001b04",
			1022 => x"01a01031",
			1023 => x"00de1031",
			1024 => x"0200be10",
			1025 => x"08001d08",
			1026 => x"0200b504",
			1027 => x"fe791031",
			1028 => x"ff7e1031",
			1029 => x"03002d04",
			1030 => x"00d51031",
			1031 => x"fed81031",
			1032 => x"04006104",
			1033 => x"018d1031",
			1034 => x"fefa1031",
			1035 => x"fe721031",
			1036 => x"0f007334",
			1037 => x"02004604",
			1038 => x"fe6b109f",
			1039 => x"0a001604",
			1040 => x"01c7109f",
			1041 => x"00008b10",
			1042 => x"06003f0c",
			1043 => x"03002108",
			1044 => x"01000904",
			1045 => x"025d109f",
			1046 => x"ff58109f",
			1047 => x"fe72109f",
			1048 => x"fe4d109f",
			1049 => x"0f005f0c",
			1050 => x"05004808",
			1051 => x"04002804",
			1052 => x"01c5109f",
			1053 => x"0100109f",
			1054 => x"feb8109f",
			1055 => x"0000c708",
			1056 => x"0f006104",
			1057 => x"0039109f",
			1058 => x"fe90109f",
			1059 => x"04006104",
			1060 => x"01f6109f",
			1061 => x"fe8e109f",
			1062 => x"fe65109f",
			1063 => x"0f005818",
			1064 => x"02006b0c",
			1065 => x"03001a08",
			1066 => x"02004604",
			1067 => x"ffe810f1",
			1068 => x"003610f1",
			1069 => x"ffcd10f1",
			1070 => x"05003608",
			1071 => x"08002004",
			1072 => x"007110f1",
			1073 => x"000110f1",
			1074 => x"ffed10f1",
			1075 => x"0200bb08",
			1076 => x"0200b904",
			1077 => x"ffac10f1",
			1078 => x"ffff10f1",
			1079 => x"0200f308",
			1080 => x"04005004",
			1081 => x"004710f1",
			1082 => x"fff710f1",
			1083 => x"ffe110f1",
			1084 => x"0f00551c",
			1085 => x"00007510",
			1086 => x"0e00360c",
			1087 => x"09001b08",
			1088 => x"00004904",
			1089 => x"fff4114d",
			1090 => x"0049114d",
			1091 => x"ffe6114d",
			1092 => x"ffb4114d",
			1093 => x"0a003108",
			1094 => x"08002004",
			1095 => x"007a114d",
			1096 => x"0000114d",
			1097 => x"ffeb114d",
			1098 => x"0200c308",
			1099 => x"0d001104",
			1100 => x"ffff114d",
			1101 => x"ffb5114d",
			1102 => x"06006c08",
			1103 => x"03005c04",
			1104 => x"0055114d",
			1105 => x"fff8114d",
			1106 => x"ffd7114d",
			1107 => x"0f00501c",
			1108 => x"02006b14",
			1109 => x"03001a10",
			1110 => x"01000708",
			1111 => x"02003a04",
			1112 => x"fff611a9",
			1113 => x"004011a9",
			1114 => x"04000704",
			1115 => x"000c11a9",
			1116 => x"ffd411a9",
			1117 => x"ffcb11a9",
			1118 => x"03002304",
			1119 => x"006e11a9",
			1120 => x"fffe11a9",
			1121 => x"0200b908",
			1122 => x"0a001c04",
			1123 => x"000411a9",
			1124 => x"ff9511a9",
			1125 => x"0f007308",
			1126 => x"04006104",
			1127 => x"006111a9",
			1128 => x"fff611a9",
			1129 => x"ffd211a9",
			1130 => x"0f006120",
			1131 => x"02006b0c",
			1132 => x"01000304",
			1133 => x"00441215",
			1134 => x"04000704",
			1135 => x"00291215",
			1136 => x"ff591215",
			1137 => x"0f005008",
			1138 => x"05002d04",
			1139 => x"00dc1215",
			1140 => x"fff41215",
			1141 => x"00009e08",
			1142 => x"02008f04",
			1143 => x"ff5d1215",
			1144 => x"00011215",
			1145 => x"00b31215",
			1146 => x"0c00200c",
			1147 => x"08001608",
			1148 => x"07002804",
			1149 => x"003a1215",
			1150 => x"ffea1215",
			1151 => x"ff2e1215",
			1152 => x"07003908",
			1153 => x"04005104",
			1154 => x"00711215",
			1155 => x"fff51215",
			1156 => x"ffe21215",
			1157 => x"06005a24",
			1158 => x"02006b0c",
			1159 => x"01000304",
			1160 => x"00411289",
			1161 => x"04000704",
			1162 => x"00281289",
			1163 => x"ff5f1289",
			1164 => x"0f005008",
			1165 => x"05002d04",
			1166 => x"00d51289",
			1167 => x"fff51289",
			1168 => x"02008f04",
			1169 => x"ff621289",
			1170 => x"0200a108",
			1171 => x"05004404",
			1172 => x"00521289",
			1173 => x"ffb31289",
			1174 => x"00be1289",
			1175 => x"0c00200c",
			1176 => x"08001608",
			1177 => x"07002804",
			1178 => x"003e1289",
			1179 => x"ffeb1289",
			1180 => x"ff381289",
			1181 => x"07003908",
			1182 => x"04005104",
			1183 => x"006e1289",
			1184 => x"fff41289",
			1185 => x"ffe01289",
			1186 => x"0f006b2c",
			1187 => x"0200921c",
			1188 => x"06003d10",
			1189 => x"02004604",
			1190 => x"ff7f12fd",
			1191 => x"03002108",
			1192 => x"08001904",
			1193 => x"00fa12fd",
			1194 => x"003112fd",
			1195 => x"ffcd12fd",
			1196 => x"00008304",
			1197 => x"fef012fd",
			1198 => x"0f005204",
			1199 => x"00cd12fd",
			1200 => x"ff2e12fd",
			1201 => x"0f006108",
			1202 => x"05004804",
			1203 => x"012512fd",
			1204 => x"ffe612fd",
			1205 => x"0200ba04",
			1206 => x"ff4e12fd",
			1207 => x"00a412fd",
			1208 => x"0b002508",
			1209 => x"0c001204",
			1210 => x"002a12fd",
			1211 => x"fee912fd",
			1212 => x"09003104",
			1213 => x"004112fd",
			1214 => x"fff212fd",
			1215 => x"02006b10",
			1216 => x"07001908",
			1217 => x"0f002504",
			1218 => x"fff21361",
			1219 => x"001e1361",
			1220 => x"04000504",
			1221 => x"00041361",
			1222 => x"ffc01361",
			1223 => x"0f006e1c",
			1224 => x"05004814",
			1225 => x"04000804",
			1226 => x"fffe1361",
			1227 => x"0200820c",
			1228 => x"02007404",
			1229 => x"00221361",
			1230 => x"00008304",
			1231 => x"ffea1361",
			1232 => x"00001361",
			1233 => x"005d1361",
			1234 => x"0d001b04",
			1235 => x"ffe41361",
			1236 => x"00121361",
			1237 => x"0d002504",
			1238 => x"ffcc1361",
			1239 => x"00091361",
			1240 => x"06006c28",
			1241 => x"00008b14",
			1242 => x"0f004210",
			1243 => x"0500210c",
			1244 => x"02004604",
			1245 => x"ffd013b5",
			1246 => x"0b001a04",
			1247 => x"009813b5",
			1248 => x"fff913b5",
			1249 => x"ffbb13b5",
			1250 => x"ff7113b5",
			1251 => x"0500480c",
			1252 => x"0f006604",
			1253 => x"00a113b5",
			1254 => x"06006404",
			1255 => x"ffe913b5",
			1256 => x"002f13b5",
			1257 => x"0200d004",
			1258 => x"ffa413b5",
			1259 => x"004713b5",
			1260 => x"ff9a13b5",
			1261 => x"00008b14",
			1262 => x"0f004210",
			1263 => x"0500210c",
			1264 => x"02004604",
			1265 => x"ffcf1431",
			1266 => x"0b001a04",
			1267 => x"009b1431",
			1268 => x"fff91431",
			1269 => x"ffb71431",
			1270 => x"ff691431",
			1271 => x"0f006614",
			1272 => x"0500480c",
			1273 => x"0b001b04",
			1274 => x"00b01431",
			1275 => x"0b001c04",
			1276 => x"fff51431",
			1277 => x"001c1431",
			1278 => x"05005104",
			1279 => x"ffdb1431",
			1280 => x"000d1431",
			1281 => x"0c00200c",
			1282 => x"08001608",
			1283 => x"07002804",
			1284 => x"00301431",
			1285 => x"fff11431",
			1286 => x"ff631431",
			1287 => x"07003908",
			1288 => x"0200d504",
			1289 => x"fff71431",
			1290 => x"005b1431",
			1291 => x"ffee1431",
			1292 => x"0f006630",
			1293 => x"02008018",
			1294 => x"0f004214",
			1295 => x"01000708",
			1296 => x"00004904",
			1297 => x"ffec14b5",
			1298 => x"008c14b5",
			1299 => x"05001208",
			1300 => x"00004104",
			1301 => x"fff014b5",
			1302 => x"002d14b5",
			1303 => x"ffad14b5",
			1304 => x"ff8314b5",
			1305 => x"05004810",
			1306 => x"0b001508",
			1307 => x"0b001404",
			1308 => x"001314b5",
			1309 => x"fff114b5",
			1310 => x"0d001d04",
			1311 => x"009214b5",
			1312 => x"000114b5",
			1313 => x"09002104",
			1314 => x"ffe114b5",
			1315 => x"001214b5",
			1316 => x"08001608",
			1317 => x"07002804",
			1318 => x"002e14b5",
			1319 => x"fff614b5",
			1320 => x"0b002004",
			1321 => x"ff6f14b5",
			1322 => x"07003904",
			1323 => x"002514b5",
			1324 => x"fff314b5",
			1325 => x"06006828",
			1326 => x"02004604",
			1327 => x"ffe71511",
			1328 => x"05003f10",
			1329 => x"0d00200c",
			1330 => x"06004e04",
			1331 => x"00601511",
			1332 => x"06005004",
			1333 => x"ffe81511",
			1334 => x"00221511",
			1335 => x"fff81511",
			1336 => x"04003608",
			1337 => x"03003904",
			1338 => x"ffe11511",
			1339 => x"00021511",
			1340 => x"0a003b04",
			1341 => x"fff41511",
			1342 => x"04005104",
			1343 => x"002a1511",
			1344 => x"fff91511",
			1345 => x"0d002504",
			1346 => x"ffd41511",
			1347 => x"00081511",
			1348 => x"0f006e30",
			1349 => x"00006e10",
			1350 => x"0d001004",
			1351 => x"002a157d",
			1352 => x"07001908",
			1353 => x"06002104",
			1354 => x"fffc157d",
			1355 => x"001e157d",
			1356 => x"ffa0157d",
			1357 => x"0f005008",
			1358 => x"05002d04",
			1359 => x"00ad157d",
			1360 => x"fff5157d",
			1361 => x"0b001810",
			1362 => x"0d001108",
			1363 => x"0a002804",
			1364 => x"ffe7157d",
			1365 => x"0045157d",
			1366 => x"04003c04",
			1367 => x"ff96157d",
			1368 => x"0006157d",
			1369 => x"07003904",
			1370 => x"0067157d",
			1371 => x"ffee157d",
			1372 => x"0d002504",
			1373 => x"ff97157d",
			1374 => x"0010157d",
			1375 => x"06006c30",
			1376 => x"02006b10",
			1377 => x"0600370c",
			1378 => x"02004604",
			1379 => x"ffdc15e1",
			1380 => x"0a001c04",
			1381 => x"005115e1",
			1382 => x"ffe915e1",
			1383 => x"ffb815e1",
			1384 => x"05003f0c",
			1385 => x"06004e04",
			1386 => x"008715e1",
			1387 => x"02009004",
			1388 => x"ffb315e1",
			1389 => x"005615e1",
			1390 => x"0000c60c",
			1391 => x"08001908",
			1392 => x"0d001304",
			1393 => x"001815e1",
			1394 => x"fff215e1",
			1395 => x"ffad15e1",
			1396 => x"04006104",
			1397 => x"004915e1",
			1398 => x"fff715e1",
			1399 => x"ffbe15e1",
			1400 => x"07002728",
			1401 => x"02005808",
			1402 => x"0d001004",
			1403 => x"da341675",
			1404 => x"d55c1675",
			1405 => x"0a001b08",
			1406 => x"09001904",
			1407 => x"e5da1675",
			1408 => x"eb6c1675",
			1409 => x"0200a10c",
			1410 => x"06004808",
			1411 => x"02006b04",
			1412 => x"d5671675",
			1413 => x"e30b1675",
			1414 => x"d55e1675",
			1415 => x"06005a04",
			1416 => x"eb451675",
			1417 => x"06006a04",
			1418 => x"dda81675",
			1419 => x"d5681675",
			1420 => x"0f006c18",
			1421 => x"0200b510",
			1422 => x"02009c08",
			1423 => x"02009004",
			1424 => x"d55c1675",
			1425 => x"d7bc1675",
			1426 => x"03003104",
			1427 => x"e9a51675",
			1428 => x"d5611675",
			1429 => x"04003b04",
			1430 => x"eb4f1675",
			1431 => x"d9ef1675",
			1432 => x"06006c08",
			1433 => x"0200d004",
			1434 => x"d55f1675",
			1435 => x"d81b1675",
			1436 => x"d55b1675",
			1437 => x"0f006c30",
			1438 => x"02009c20",
			1439 => x"0d000e04",
			1440 => x"00c316e9",
			1441 => x"0f00420c",
			1442 => x"02005904",
			1443 => x"ff8716e9",
			1444 => x"03002104",
			1445 => x"00dd16e9",
			1446 => x"ffb316e9",
			1447 => x"00008b04",
			1448 => x"ff0916e9",
			1449 => x"0d001304",
			1450 => x"ffa616e9",
			1451 => x"0b001804",
			1452 => x"ffe216e9",
			1453 => x"008616e9",
			1454 => x"0f006608",
			1455 => x"05004a04",
			1456 => x"00ee16e9",
			1457 => x"fff916e9",
			1458 => x"0f006a04",
			1459 => x"ffb816e9",
			1460 => x"004816e9",
			1461 => x"01000304",
			1462 => x"001d16e9",
			1463 => x"0d002504",
			1464 => x"ff2b16e9",
			1465 => x"001d16e9",
			1466 => x"0600682c",
			1467 => x"0200ac20",
			1468 => x"0600501c",
			1469 => x"02006b10",
			1470 => x"0600370c",
			1471 => x"02004604",
			1472 => x"ffc6174d",
			1473 => x"0a001e04",
			1474 => x"007d174d",
			1475 => x"ffdb174d",
			1476 => x"ff89174d",
			1477 => x"04002208",
			1478 => x"08001f04",
			1479 => x"00c1174d",
			1480 => x"fffc174d",
			1481 => x"ffd8174d",
			1482 => x"ff6f174d",
			1483 => x"03003d04",
			1484 => x"00a7174d",
			1485 => x"03004404",
			1486 => x"ffef174d",
			1487 => x"001d174d",
			1488 => x"0d002504",
			1489 => x"ff81174d",
			1490 => x"0012174d",
			1491 => x"0600682c",
			1492 => x"0200b928",
			1493 => x"0f004b14",
			1494 => x"0300230c",
			1495 => x"02004604",
			1496 => x"ffdc17b1",
			1497 => x"0d001804",
			1498 => x"007e17b1",
			1499 => x"000217b1",
			1500 => x"0a002d04",
			1501 => x"ffd717b1",
			1502 => x"000217b1",
			1503 => x"02008b04",
			1504 => x"ffa317b1",
			1505 => x"0f005808",
			1506 => x"0b001904",
			1507 => x"005717b1",
			1508 => x"fff617b1",
			1509 => x"0d001204",
			1510 => x"000217b1",
			1511 => x"ffb117b1",
			1512 => x"007517b1",
			1513 => x"0d002504",
			1514 => x"ffbb17b1",
			1515 => x"000b17b1",
			1516 => x"06006c34",
			1517 => x"0200a524",
			1518 => x"0f004b18",
			1519 => x"03002310",
			1520 => x"02004604",
			1521 => x"ff68181d",
			1522 => x"02006b08",
			1523 => x"06003104",
			1524 => x"00e3181d",
			1525 => x"ff8a181d",
			1526 => x"012a181d",
			1527 => x"07002404",
			1528 => x"ff4d181d",
			1529 => x"0018181d",
			1530 => x"02008b04",
			1531 => x"fee0181d",
			1532 => x"0f005804",
			1533 => x"00b0181d",
			1534 => x"ff0d181d",
			1535 => x"05004808",
			1536 => x"0f006604",
			1537 => x"0142181d",
			1538 => x"0050181d",
			1539 => x"0200d004",
			1540 => x"ff48181d",
			1541 => x"00a6181d",
			1542 => x"fee0181d",
			1543 => x"06006c38",
			1544 => x"02006b14",
			1545 => x"0e002e0c",
			1546 => x"02004604",
			1547 => x"ff901891",
			1548 => x"0d001304",
			1549 => x"00b31891",
			1550 => x"ffed1891",
			1551 => x"07002004",
			1552 => x"ff2b1891",
			1553 => x"fff21891",
			1554 => x"0f00500c",
			1555 => x"05002d08",
			1556 => x"08002004",
			1557 => x"01321891",
			1558 => x"001a1891",
			1559 => x"ffed1891",
			1560 => x"0200a508",
			1561 => x"04001804",
			1562 => x"ffef1891",
			1563 => x"ff101891",
			1564 => x"05004808",
			1565 => x"0f006604",
			1566 => x"010b1891",
			1567 => x"003e1891",
			1568 => x"0200d004",
			1569 => x"ff6f1891",
			1570 => x"008d1891",
			1571 => x"ff161891",
			1572 => x"0f007330",
			1573 => x"02008218",
			1574 => x"0a001408",
			1575 => x"00005204",
			1576 => x"fff018f5",
			1577 => x"004918f5",
			1578 => x"0b001204",
			1579 => x"001018f5",
			1580 => x"06003e08",
			1581 => x"06003804",
			1582 => x"ffe618f5",
			1583 => x"001418f5",
			1584 => x"ffaf18f5",
			1585 => x"04005114",
			1586 => x"09001a04",
			1587 => x"000118f5",
			1588 => x"05004504",
			1589 => x"005518f5",
			1590 => x"05005308",
			1591 => x"05004804",
			1592 => x"000418f5",
			1593 => x"ffed18f5",
			1594 => x"001818f5",
			1595 => x"fff718f5",
			1596 => x"ffdd18f5",
			1597 => x"0f00733c",
			1598 => x"0200a528",
			1599 => x"0f004b14",
			1600 => x"0300230c",
			1601 => x"02004604",
			1602 => x"ff5f1971",
			1603 => x"0f004304",
			1604 => x"011d1971",
			1605 => x"005a1971",
			1606 => x"07002404",
			1607 => x"ff461971",
			1608 => x"001c1971",
			1609 => x"0b00180c",
			1610 => x"02009908",
			1611 => x"01000e04",
			1612 => x"fecf1971",
			1613 => x"ffce1971",
			1614 => x"ffd81971",
			1615 => x"03002b04",
			1616 => x"00d91971",
			1617 => x"ff1e1971",
			1618 => x"05004808",
			1619 => x"0f006604",
			1620 => x"014d1971",
			1621 => x"005c1971",
			1622 => x"0200d004",
			1623 => x"ff3f1971",
			1624 => x"03008404",
			1625 => x"00b61971",
			1626 => x"fff41971",
			1627 => x"fed71971",
			1628 => x"0f007334",
			1629 => x"0200ac24",
			1630 => x"0f00581c",
			1631 => x"02007110",
			1632 => x"06003c0c",
			1633 => x"02004604",
			1634 => x"ff0a19dd",
			1635 => x"09001b04",
			1636 => x"014b19dd",
			1637 => x"ff7919dd",
			1638 => x"feb719dd",
			1639 => x"04002508",
			1640 => x"0b001604",
			1641 => x"006019dd",
			1642 => x"017419dd",
			1643 => x"ffba19dd",
			1644 => x"0b001a04",
			1645 => x"feab19dd",
			1646 => x"ffe619dd",
			1647 => x"05004804",
			1648 => x"015619dd",
			1649 => x"0200d004",
			1650 => x"ff1919dd",
			1651 => x"0500bf04",
			1652 => x"00f119dd",
			1653 => x"ffe619dd",
			1654 => x"fe9619dd",
			1655 => x"0f007328",
			1656 => x"02005004",
			1657 => x"fe871a31",
			1658 => x"0500481c",
			1659 => x"0200aa14",
			1660 => x"0f005810",
			1661 => x"02008008",
			1662 => x"03002104",
			1663 => x"00d61a31",
			1664 => x"fe8b1a31",
			1665 => x"04002804",
			1666 => x"01a11a31",
			1667 => x"00271a31",
			1668 => x"fe9a1a31",
			1669 => x"0200ba04",
			1670 => x"00ff1a31",
			1671 => x"01a11a31",
			1672 => x"0200d004",
			1673 => x"fe821a31",
			1674 => x"01381a31",
			1675 => x"fe6f1a31",
			1676 => x"0f007338",
			1677 => x"02007110",
			1678 => x"0f003c0c",
			1679 => x"02004604",
			1680 => x"ff901aa5",
			1681 => x"09001b04",
			1682 => x"00d61aa5",
			1683 => x"ffc21aa5",
			1684 => x"ff211aa5",
			1685 => x"06004c0c",
			1686 => x"05002d08",
			1687 => x"08002004",
			1688 => x"01201aa5",
			1689 => x"00171aa5",
			1690 => x"00191aa5",
			1691 => x"0200ac0c",
			1692 => x"0f005808",
			1693 => x"02008c04",
			1694 => x"ff6a1aa5",
			1695 => x"00861aa5",
			1696 => x"ff231aa5",
			1697 => x"0400610c",
			1698 => x"0200bc08",
			1699 => x"0f006604",
			1700 => x"00a21aa5",
			1701 => x"ff8d1aa5",
			1702 => x"00fc1aa5",
			1703 => x"ffdc1aa5",
			1704 => x"ff211aa5",
			1705 => x"0f006c34",
			1706 => x"0200a128",
			1707 => x"05002d20",
			1708 => x"0d000e04",
			1709 => x"00c91b21",
			1710 => x"02006b0c",
			1711 => x"03000c08",
			1712 => x"0c001804",
			1713 => x"00481b21",
			1714 => x"fff81b21",
			1715 => x"ff4c1b21",
			1716 => x"09001d08",
			1717 => x"06004704",
			1718 => x"005d1b21",
			1719 => x"ff691b21",
			1720 => x"01000d04",
			1721 => x"00ce1b21",
			1722 => x"00061b21",
			1723 => x"04002204",
			1724 => x"00001b21",
			1725 => x"ff381b21",
			1726 => x"0f006604",
			1727 => x"00e91b21",
			1728 => x"0f006a04",
			1729 => x"ffbb1b21",
			1730 => x"004e1b21",
			1731 => x"01000304",
			1732 => x"001e1b21",
			1733 => x"0d002504",
			1734 => x"ff221b21",
			1735 => x"001e1b21",
			1736 => x"0f00733c",
			1737 => x"02006b10",
			1738 => x"08001604",
			1739 => x"00cc1b9d",
			1740 => x"04000704",
			1741 => x"00e91b9d",
			1742 => x"09001604",
			1743 => x"fdb21b9d",
			1744 => x"fe731b9d",
			1745 => x"0f005510",
			1746 => x"02008008",
			1747 => x"06004404",
			1748 => x"01631b9d",
			1749 => x"fe821b9d",
			1750 => x"04002104",
			1751 => x"01af1b9d",
			1752 => x"01261b9d",
			1753 => x"0200b90c",
			1754 => x"06005a08",
			1755 => x"02009804",
			1756 => x"fe791b9d",
			1757 => x"012b1b9d",
			1758 => x"fe6e1b9d",
			1759 => x"0400610c",
			1760 => x"0200c308",
			1761 => x"0f006c04",
			1762 => x"01901b9d",
			1763 => x"fed11b9d",
			1764 => x"01c61b9d",
			1765 => x"fead1b9d",
			1766 => x"fe6a1b9d",
			1767 => x"0f007338",
			1768 => x"02009c24",
			1769 => x"0d000e04",
			1770 => x"016b1c11",
			1771 => x"0f004b14",
			1772 => x"02006b0c",
			1773 => x"03001308",
			1774 => x"00003b04",
			1775 => x"ff0a1c11",
			1776 => x"01061c11",
			1777 => x"fe951c11",
			1778 => x"01000904",
			1779 => x"01801c11",
			1780 => x"00621c11",
			1781 => x"02009204",
			1782 => x"fe671c11",
			1783 => x"04002d04",
			1784 => x"00a41c11",
			1785 => x"ff0b1c11",
			1786 => x"0f006104",
			1787 => x"01861c11",
			1788 => x"0000cc08",
			1789 => x"08001d04",
			1790 => x"fea41c11",
			1791 => x"ff8f1c11",
			1792 => x"04006104",
			1793 => x"017e1c11",
			1794 => x"ff3a1c11",
			1795 => x"fe7b1c11",
			1796 => x"0600683c",
			1797 => x"02005008",
			1798 => x"0d001004",
			1799 => x"ffb91c9d",
			1800 => x"fe4e1c9d",
			1801 => x"05003e24",
			1802 => x"02008b14",
			1803 => x"05001b0c",
			1804 => x"0f004008",
			1805 => x"09001b04",
			1806 => x"05d01c9d",
			1807 => x"048a1c9d",
			1808 => x"02bf1c9d",
			1809 => x"01000704",
			1810 => x"01f11c9d",
			1811 => x"fe481c9d",
			1812 => x"06005e0c",
			1813 => x"06005108",
			1814 => x"09002004",
			1815 => x"04a41c9d",
			1816 => x"054a1c9d",
			1817 => x"04531c9d",
			1818 => x"032d1c9d",
			1819 => x"0200ca0c",
			1820 => x"01000608",
			1821 => x"05004904",
			1822 => x"01cb1c9d",
			1823 => x"fe571c9d",
			1824 => x"fe4c1c9d",
			1825 => x"048b1c9d",
			1826 => x"0d002504",
			1827 => x"fe4e1c9d",
			1828 => x"0e009d04",
			1829 => x"000d1c9d",
			1830 => x"fe5e1c9d",
			1831 => x"0f007334",
			1832 => x"02004604",
			1833 => x"fe821d09",
			1834 => x"0500321c",
			1835 => x"0f005410",
			1836 => x"0200710c",
			1837 => x"03001a04",
			1838 => x"01b41d09",
			1839 => x"05002c04",
			1840 => x"fe7b1d09",
			1841 => x"00811d09",
			1842 => x"01a11d09",
			1843 => x"02009004",
			1844 => x"fe811d09",
			1845 => x"08001b04",
			1846 => x"00781d09",
			1847 => x"01911d09",
			1848 => x"0000c60c",
			1849 => x"0e005208",
			1850 => x"00009e04",
			1851 => x"fe841d09",
			1852 => x"01311d09",
			1853 => x"fe751d09",
			1854 => x"04006104",
			1855 => x"01a21d09",
			1856 => x"fec31d09",
			1857 => x"fe6c1d09",
			1858 => x"06006840",
			1859 => x"02005008",
			1860 => x"01000404",
			1861 => x"ff8d1d9d",
			1862 => x"fe4a1d9d",
			1863 => x"05004028",
			1864 => x"00009414",
			1865 => x"0a001908",
			1866 => x"06003504",
			1867 => x"086a1d9d",
			1868 => x"06121d9d",
			1869 => x"01000704",
			1870 => x"02791d9d",
			1871 => x"03001f04",
			1872 => x"ffa41d9d",
			1873 => x"fe461d9d",
			1874 => x"0200a50c",
			1875 => x"0f005908",
			1876 => x"04001304",
			1877 => x"06ce1d9d",
			1878 => x"08751d9d",
			1879 => x"fe441d9d",
			1880 => x"0f006204",
			1881 => x"06961d9d",
			1882 => x"087a1d9d",
			1883 => x"0000d50c",
			1884 => x"0e005208",
			1885 => x"08001904",
			1886 => x"00af1d9d",
			1887 => x"fe541d9d",
			1888 => x"fe481d9d",
			1889 => x"06c81d9d",
			1890 => x"0d002504",
			1891 => x"fe4a1d9d",
			1892 => x"03003804",
			1893 => x"fe561d9d",
			1894 => x"ffeb1d9d",
			1895 => x"0f006e3c",
			1896 => x"02004604",
			1897 => x"fe5f1e29",
			1898 => x"05002f20",
			1899 => x"02006b08",
			1900 => x"03001a04",
			1901 => x"02521e29",
			1902 => x"fe551e29",
			1903 => x"0600510c",
			1904 => x"01000804",
			1905 => x"028a1e29",
			1906 => x"00008104",
			1907 => x"01371e29",
			1908 => x"02331e29",
			1909 => x"02009904",
			1910 => x"fe461e29",
			1911 => x"01000a04",
			1912 => x"01b51e29",
			1913 => x"024e1e29",
			1914 => x"0200bc0c",
			1915 => x"0000a904",
			1916 => x"fe531e29",
			1917 => x"0f006704",
			1918 => x"01b91e29",
			1919 => x"fe621e29",
			1920 => x"03006108",
			1921 => x"04003104",
			1922 => x"022b1e29",
			1923 => x"030c1e29",
			1924 => x"fe3f1e29",
			1925 => x"0d002504",
			1926 => x"fe5c1e29",
			1927 => x"0600b604",
			1928 => x"00e81e29",
			1929 => x"fe781e29",
			1930 => x"0f007340",
			1931 => x"01000510",
			1932 => x"03003a0c",
			1933 => x"04001408",
			1934 => x"07002104",
			1935 => x"00901ead",
			1936 => x"ff641ead",
			1937 => x"01391ead",
			1938 => x"ff9a1ead",
			1939 => x"00008b14",
			1940 => x"05001b10",
			1941 => x"08001804",
			1942 => x"00c01ead",
			1943 => x"0c001404",
			1944 => x"ff101ead",
			1945 => x"09002004",
			1946 => x"009f1ead",
			1947 => x"ff961ead",
			1948 => x"fed01ead",
			1949 => x"05003208",
			1950 => x"0b001504",
			1951 => x"00031ead",
			1952 => x"01341ead",
			1953 => x"0000cc0c",
			1954 => x"08001804",
			1955 => x"004b1ead",
			1956 => x"0d001a04",
			1957 => x"fedb1ead",
			1958 => x"ffe71ead",
			1959 => x"04006104",
			1960 => x"010a1ead",
			1961 => x"ffb41ead",
			1962 => x"fec31ead",
			1963 => x"0f00733c",
			1964 => x"0200ac2c",
			1965 => x"0f005524",
			1966 => x"02007114",
			1967 => x"0f004010",
			1968 => x"09001b08",
			1969 => x"00004904",
			1970 => x"ff971f29",
			1971 => x"01061f29",
			1972 => x"08001904",
			1973 => x"00051f29",
			1974 => x"ff501f29",
			1975 => x"fecf1f29",
			1976 => x"0800200c",
			1977 => x"04002508",
			1978 => x"0f005004",
			1979 => x"015c1f29",
			1980 => x"00631f29",
			1981 => x"00491f29",
			1982 => x"ffed1f29",
			1983 => x"0d001904",
			1984 => x"feda1f29",
			1985 => x"ffe01f29",
			1986 => x"0400610c",
			1987 => x"0f006c04",
			1988 => x"013c1f29",
			1989 => x"0f007004",
			1990 => x"ffcb1f29",
			1991 => x"003f1f29",
			1992 => x"ffb01f29",
			1993 => x"febf1f29",
			1994 => x"0f007338",
			1995 => x"02005004",
			1996 => x"fe621f9d",
			1997 => x"05003e24",
			1998 => x"00008b10",
			1999 => x"0a001908",
			2000 => x"07001e04",
			2001 => x"02321f9d",
			2002 => x"01931f9d",
			2003 => x"0d001204",
			2004 => x"00281f9d",
			2005 => x"fe551f9d",
			2006 => x"0f005a08",
			2007 => x"0000a104",
			2008 => x"02581f9d",
			2009 => x"01f61f9d",
			2010 => x"0000bc04",
			2011 => x"fe5a1f9d",
			2012 => x"06005d04",
			2013 => x"01e71f9d",
			2014 => x"024c1f9d",
			2015 => x"0000e10c",
			2016 => x"0f006608",
			2017 => x"0200a504",
			2018 => x"fe641f9d",
			2019 => x"02201f9d",
			2020 => x"fe5a1f9d",
			2021 => x"02d81f9d",
			2022 => x"fe5f1f9d",
			2023 => x"0f00733c",
			2024 => x"0000c634",
			2025 => x"0f005828",
			2026 => x"02007118",
			2027 => x"0100070c",
			2028 => x"03001a08",
			2029 => x"00004304",
			2030 => x"ffa92019",
			2031 => x"01482019",
			2032 => x"ffeb2019",
			2033 => x"04000704",
			2034 => x"00572019",
			2035 => x"0a000b04",
			2036 => x"fffa2019",
			2037 => x"fec92019",
			2038 => x"0500360c",
			2039 => x"0b001504",
			2040 => x"00762019",
			2041 => x"08002004",
			2042 => x"01732019",
			2043 => x"006c2019",
			2044 => x"fff22019",
			2045 => x"0200b504",
			2046 => x"febc2019",
			2047 => x"0000c304",
			2048 => x"00082019",
			2049 => x"ffdc2019",
			2050 => x"04006104",
			2051 => x"01522019",
			2052 => x"ff972019",
			2053 => x"fea02019",
			2054 => x"0f007330",
			2055 => x"02004604",
			2056 => x"fe76207d",
			2057 => x"0d000e04",
			2058 => x"020d207d",
			2059 => x"02006b0c",
			2060 => x"06003308",
			2061 => x"05001c04",
			2062 => x"00e2207d",
			2063 => x"febd207d",
			2064 => x"fded207d",
			2065 => x"06004c0c",
			2066 => x"00008308",
			2067 => x"03002104",
			2068 => x"0190207d",
			2069 => x"fe8c207d",
			2070 => x"01bc207d",
			2071 => x"0200a508",
			2072 => x"04001804",
			2073 => x"ffe1207d",
			2074 => x"fe6e207d",
			2075 => x"0f006604",
			2076 => x"019d207d",
			2077 => x"0041207d",
			2078 => x"fe69207d",
			2079 => x"0f00733c",
			2080 => x"08001404",
			2081 => x"019c20f9",
			2082 => x"02008214",
			2083 => x"0f003f10",
			2084 => x"02005004",
			2085 => x"fead20f9",
			2086 => x"03002108",
			2087 => x"08001904",
			2088 => x"017520f9",
			2089 => x"007120f9",
			2090 => x"ff4520f9",
			2091 => x"fe5520f9",
			2092 => x"06005a14",
			2093 => x"05004810",
			2094 => x"0b001508",
			2095 => x"02008f04",
			2096 => x"ff4920f9",
			2097 => x"00d120f9",
			2098 => x"01001104",
			2099 => x"017620f9",
			2100 => x"003420f9",
			2101 => x"ff9920f9",
			2102 => x"0000cc08",
			2103 => x"0200ba04",
			2104 => x"fe9120f9",
			2105 => x"ff9920f9",
			2106 => x"04006104",
			2107 => x"018020f9",
			2108 => x"ff2120f9",
			2109 => x"fe7920f9",
			2110 => x"0f007340",
			2111 => x"08001504",
			2112 => x"0162217f",
			2113 => x"00006e10",
			2114 => x"04000708",
			2115 => x"0e002004",
			2116 => x"ff97217f",
			2117 => x"00b1217f",
			2118 => x"08001804",
			2119 => x"ffd4217f",
			2120 => x"fe2d217f",
			2121 => x"0f005514",
			2122 => x"00008b0c",
			2123 => x"06003f08",
			2124 => x"0c001704",
			2125 => x"019b217f",
			2126 => x"008e217f",
			2127 => x"fe95217f",
			2128 => x"0b001b04",
			2129 => x"019e217f",
			2130 => x"00cb217f",
			2131 => x"0200c010",
			2132 => x"08001d08",
			2133 => x"0200b504",
			2134 => x"fe7c217f",
			2135 => x"ff6f217f",
			2136 => x"05003304",
			2137 => x"00cd217f",
			2138 => x"fee2217f",
			2139 => x"04006104",
			2140 => x"018b217f",
			2141 => x"ff0a217f",
			2142 => x"fe74217f",
			2143 => x"05002118",
			2144 => x"0f005610",
			2145 => x"02004604",
			2146 => x"ffe621d9",
			2147 => x"08002008",
			2148 => x"03001f04",
			2149 => x"007421d9",
			2150 => x"000321d9",
			2151 => x"fffb21d9",
			2152 => x"0000a404",
			2153 => x"ffe021d9",
			2154 => x"000521d9",
			2155 => x"0000a90c",
			2156 => x"09002004",
			2157 => x"ff9e21d9",
			2158 => x"04002204",
			2159 => x"002921d9",
			2160 => x"ffd521d9",
			2161 => x"0f006c04",
			2162 => x"005521d9",
			2163 => x"07002704",
			2164 => x"000921d9",
			2165 => x"ffc021d9",
			2166 => x"02006b10",
			2167 => x"07001908",
			2168 => x"06002404",
			2169 => x"fff3222d",
			2170 => x"001f222d",
			2171 => x"04000504",
			2172 => x"0005222d",
			2173 => x"ffc7222d",
			2174 => x"0f005008",
			2175 => x"03002304",
			2176 => x"0066222d",
			2177 => x"fffc222d",
			2178 => x"0200a504",
			2179 => x"ffbf222d",
			2180 => x"0f006c04",
			2181 => x"0048222d",
			2182 => x"0d002508",
			2183 => x"07002604",
			2184 => x"0007222d",
			2185 => x"ffcd222d",
			2186 => x"0008222d",
			2187 => x"0f006624",
			2188 => x"02006b10",
			2189 => x"03001a0c",
			2190 => x"09001504",
			2191 => x"ffd52291",
			2192 => x"00004804",
			2193 => x"ffeb2291",
			2194 => x"00542291",
			2195 => x"ffb12291",
			2196 => x"0f005008",
			2197 => x"03002304",
			2198 => x"009c2291",
			2199 => x"00022291",
			2200 => x"0200a108",
			2201 => x"0b001804",
			2202 => x"ff9c2291",
			2203 => x"fffa2291",
			2204 => x"00732291",
			2205 => x"0b002308",
			2206 => x"08001504",
			2207 => x"001b2291",
			2208 => x"ff812291",
			2209 => x"09003004",
			2210 => x"002c2291",
			2211 => x"fffb2291",
			2212 => x"0f004b1c",
			2213 => x"03002310",
			2214 => x"02004604",
			2215 => x"ffe922f5",
			2216 => x"08001d04",
			2217 => x"006922f5",
			2218 => x"08001f04",
			2219 => x"fff622f5",
			2220 => x"000422f5",
			2221 => x"08001d04",
			2222 => x"ffe322f5",
			2223 => x"08002004",
			2224 => x"000622f5",
			2225 => x"fffc22f5",
			2226 => x"02008b04",
			2227 => x"ffb522f5",
			2228 => x"06006c10",
			2229 => x"05004508",
			2230 => x"04001504",
			2231 => x"ffff22f5",
			2232 => x"005a22f5",
			2233 => x"0200d004",
			2234 => x"ffcf22f5",
			2235 => x"001a22f5",
			2236 => x"ffd522f5",
			2237 => x"01000514",
			2238 => x"04001408",
			2239 => x"0a001404",
			2240 => x"00172369",
			2241 => x"ffd52369",
			2242 => x"0d001308",
			2243 => x"07002704",
			2244 => x"00602369",
			2245 => x"fffa2369",
			2246 => x"fff42369",
			2247 => x"05001b10",
			2248 => x"00006b08",
			2249 => x"01000c04",
			2250 => x"ffde2369",
			2251 => x"000a2369",
			2252 => x"06004b04",
			2253 => x"00402369",
			2254 => x"00002369",
			2255 => x"0c001c08",
			2256 => x"08001504",
			2257 => x"00002369",
			2258 => x"ffab2369",
			2259 => x"0700390c",
			2260 => x"04005008",
			2261 => x"00009704",
			2262 => x"fffb2369",
			2263 => x"003e2369",
			2264 => x"fff92369",
			2265 => x"fff32369",
			2266 => x"06006c20",
			2267 => x"02004604",
			2268 => x"ffde23ad",
			2269 => x"05003f08",
			2270 => x"0d001f04",
			2271 => x"006723ad",
			2272 => x"fff823ad",
			2273 => x"0d001a0c",
			2274 => x"01000504",
			2275 => x"001823ad",
			2276 => x"08001804",
			2277 => x"000023ad",
			2278 => x"ffbf23ad",
			2279 => x"04005104",
			2280 => x"003223ad",
			2281 => x"fffa23ad",
			2282 => x"ffc923ad",
			2283 => x"02006b10",
			2284 => x"07001908",
			2285 => x"0f002504",
			2286 => x"fff32411",
			2287 => x"001e2411",
			2288 => x"04000504",
			2289 => x"00052411",
			2290 => x"ffc32411",
			2291 => x"0f006e1c",
			2292 => x"05004814",
			2293 => x"04000804",
			2294 => x"fffe2411",
			2295 => x"0200820c",
			2296 => x"02007404",
			2297 => x"00222411",
			2298 => x"02007e04",
			2299 => x"ffea2411",
			2300 => x"00002411",
			2301 => x"00592411",
			2302 => x"0d001b04",
			2303 => x"ffe42411",
			2304 => x"00122411",
			2305 => x"0d002504",
			2306 => x"ffce2411",
			2307 => x"00092411",
			2308 => x"0600662c",
			2309 => x"02006b10",
			2310 => x"0600370c",
			2311 => x"02004604",
			2312 => x"feeb247d",
			2313 => x"0a001c04",
			2314 => x"0176247d",
			2315 => x"ff5c247d",
			2316 => x"fe7c247d",
			2317 => x"0f005008",
			2318 => x"05002d04",
			2319 => x"018b247d",
			2320 => x"ffff247d",
			2321 => x"0200a508",
			2322 => x"0f005504",
			2323 => x"0018247d",
			2324 => x"febb247d",
			2325 => x"05004804",
			2326 => x"0171247d",
			2327 => x"0200b904",
			2328 => x"ff35247d",
			2329 => x"00e5247d",
			2330 => x"0d002504",
			2331 => x"fe86247d",
			2332 => x"0c002904",
			2333 => x"0097247d",
			2334 => x"ffd6247d",
			2335 => x"0600682c",
			2336 => x"02006b10",
			2337 => x"07001908",
			2338 => x"0f002604",
			2339 => x"ffec24d9",
			2340 => x"003224d9",
			2341 => x"04000504",
			2342 => x"000824d9",
			2343 => x"ffad24d9",
			2344 => x"05003b0c",
			2345 => x"06004e04",
			2346 => x"007f24d9",
			2347 => x"02009004",
			2348 => x"ffb824d9",
			2349 => x"004a24d9",
			2350 => x"0000c60c",
			2351 => x"0c001708",
			2352 => x"04003404",
			2353 => x"fff624d9",
			2354 => x"001724d9",
			2355 => x"ffa424d9",
			2356 => x"004c24d9",
			2357 => x"ffb424d9",
			2358 => x"0f00732c",
			2359 => x"02006b0c",
			2360 => x"07001a08",
			2361 => x"01000504",
			2362 => x"00fe2535",
			2363 => x"ff962535",
			2364 => x"feb82535",
			2365 => x"0f006114",
			2366 => x"0200900c",
			2367 => x"0f005008",
			2368 => x"03002304",
			2369 => x"013e2535",
			2370 => x"ffb02535",
			2371 => x"fef42535",
			2372 => x"05004804",
			2373 => x"01692535",
			2374 => x"ffda2535",
			2375 => x"0000cc04",
			2376 => x"fed42535",
			2377 => x"04006104",
			2378 => x"013f2535",
			2379 => x"ffa52535",
			2380 => x"feaf2535",
			2381 => x"0f00732c",
			2382 => x"02008218",
			2383 => x"0a001408",
			2384 => x"00005204",
			2385 => x"fff02591",
			2386 => x"00472591",
			2387 => x"0b001204",
			2388 => x"00102591",
			2389 => x"06003e08",
			2390 => x"06003804",
			2391 => x"ffe72591",
			2392 => x"00152591",
			2393 => x"ffb22591",
			2394 => x"04005110",
			2395 => x"0200a50c",
			2396 => x"05003508",
			2397 => x"0b001504",
			2398 => x"fff02591",
			2399 => x"003e2591",
			2400 => x"ffd72591",
			2401 => x"00552591",
			2402 => x"fff72591",
			2403 => x"ffdd2591",
			2404 => x"06006634",
			2405 => x"02006b14",
			2406 => x"07001a08",
			2407 => x"00004504",
			2408 => x"ff5d260d",
			2409 => x"0160260d",
			2410 => x"06003708",
			2411 => x"0f003304",
			2412 => x"ff04260d",
			2413 => x"00bc260d",
			2414 => x"fe8b260d",
			2415 => x"0f005008",
			2416 => x"05002d04",
			2417 => x"0182260d",
			2418 => x"fffb260d",
			2419 => x"0200a508",
			2420 => x"04001804",
			2421 => x"fff7260d",
			2422 => x"feac260d",
			2423 => x"05004808",
			2424 => x"06005f04",
			2425 => x"0189260d",
			2426 => x"00ad260d",
			2427 => x"0200b904",
			2428 => x"ff3f260d",
			2429 => x"00d9260d",
			2430 => x"0d002504",
			2431 => x"fe8a260d",
			2432 => x"0c002904",
			2433 => x"0090260d",
			2434 => x"ffd9260d",
			2435 => x"06006c30",
			2436 => x"02006b10",
			2437 => x"0600370c",
			2438 => x"02004604",
			2439 => x"ffdd2671",
			2440 => x"0a001c04",
			2441 => x"00502671",
			2442 => x"ffea2671",
			2443 => x"ffba2671",
			2444 => x"05003f0c",
			2445 => x"06004e04",
			2446 => x"00822671",
			2447 => x"02009004",
			2448 => x"ffb62671",
			2449 => x"00532671",
			2450 => x"0000c60c",
			2451 => x"08001908",
			2452 => x"0d001304",
			2453 => x"00192671",
			2454 => x"fff32671",
			2455 => x"ffaf2671",
			2456 => x"04006104",
			2457 => x"00472671",
			2458 => x"fff72671",
			2459 => x"ffc02671",
			2460 => x"0f006624",
			2461 => x"0200991c",
			2462 => x"06003d10",
			2463 => x"02004604",
			2464 => x"ff7726f5",
			2465 => x"08001904",
			2466 => x"010326f5",
			2467 => x"03001704",
			2468 => x"008626f5",
			2469 => x"ff8b26f5",
			2470 => x"00008304",
			2471 => x"fee426f5",
			2472 => x"0f005204",
			2473 => x"00e626f5",
			2474 => x"ff2f26f5",
			2475 => x"05004804",
			2476 => x"012326f5",
			2477 => x"ffef26f5",
			2478 => x"08001504",
			2479 => x"006326f5",
			2480 => x"0b002314",
			2481 => x"0c00230c",
			2482 => x"08001608",
			2483 => x"0c001404",
			2484 => x"000b26f5",
			2485 => x"ffe726f5",
			2486 => x"fed526f5",
			2487 => x"09002c04",
			2488 => x"001026f5",
			2489 => x"fff026f5",
			2490 => x"07003b04",
			2491 => x"005a26f5",
			2492 => x"ffe426f5",
			2493 => x"0f007330",
			2494 => x"02006b10",
			2495 => x"0600370c",
			2496 => x"02004604",
			2497 => x"ff892759",
			2498 => x"0a001c04",
			2499 => x"00b92759",
			2500 => x"ffc32759",
			2501 => x"ff222759",
			2502 => x"0f005008",
			2503 => x"05002d04",
			2504 => x"01342759",
			2505 => x"ffeb2759",
			2506 => x"0200a508",
			2507 => x"04001804",
			2508 => x"ffee2759",
			2509 => x"ff062759",
			2510 => x"05004808",
			2511 => x"0f006604",
			2512 => x"01122759",
			2513 => x"00442759",
			2514 => x"0200d004",
			2515 => x"ff682759",
			2516 => x"00932759",
			2517 => x"ff0c2759",
			2518 => x"0f007334",
			2519 => x"02006b10",
			2520 => x"0600370c",
			2521 => x"08001604",
			2522 => x"003d27c5",
			2523 => x"04000704",
			2524 => x"001527c5",
			2525 => x"ffca27c5",
			2526 => x"ffbc27c5",
			2527 => x"05003e10",
			2528 => x"02008208",
			2529 => x"06004804",
			2530 => x"003f27c5",
			2531 => x"ffc627c5",
			2532 => x"04000d04",
			2533 => x"000227c5",
			2534 => x"007927c5",
			2535 => x"0000c60c",
			2536 => x"0c001708",
			2537 => x"04003404",
			2538 => x"fff927c5",
			2539 => x"001627c5",
			2540 => x"ffb127c5",
			2541 => x"04006104",
			2542 => x"004a27c5",
			2543 => x"fff927c5",
			2544 => x"ffc527c5",
			2545 => x"0f007334",
			2546 => x"02006b0c",
			2547 => x"08001604",
			2548 => x"00d72831",
			2549 => x"04000704",
			2550 => x"00402831",
			2551 => x"fe6c2831",
			2552 => x"05003214",
			2553 => x"0600510c",
			2554 => x"01000904",
			2555 => x"01922831",
			2556 => x"00008604",
			2557 => x"ffa52831",
			2558 => x"01602831",
			2559 => x"0000a404",
			2560 => x"fed42831",
			2561 => x"010a2831",
			2562 => x"0200ca0c",
			2563 => x"0f005808",
			2564 => x"00008b04",
			2565 => x"ff032831",
			2566 => x"00852831",
			2567 => x"fe952831",
			2568 => x"04006104",
			2569 => x"016e2831",
			2570 => x"ff672831",
			2571 => x"fe812831",
			2572 => x"0f006e2c",
			2573 => x"0200ac24",
			2574 => x"0f005520",
			2575 => x"02006b10",
			2576 => x"0600370c",
			2577 => x"09001b08",
			2578 => x"00004904",
			2579 => x"ffb1289d",
			2580 => x"00e8289d",
			2581 => x"ff76289d",
			2582 => x"fefa289d",
			2583 => x"05002d08",
			2584 => x"05002304",
			2585 => x"0136289d",
			2586 => x"0068289d",
			2587 => x"00008804",
			2588 => x"ff73289d",
			2589 => x"002c289d",
			2590 => x"ff0b289d",
			2591 => x"04006604",
			2592 => x"010b289d",
			2593 => x"ffd2289d",
			2594 => x"0d002504",
			2595 => x"fedc289d",
			2596 => x"04002e04",
			2597 => x"fffa289d",
			2598 => x"0039289d",
			2599 => x"0f006e34",
			2600 => x"00006e10",
			2601 => x"0d001004",
			2602 => x"00282911",
			2603 => x"07001908",
			2604 => x"06002104",
			2605 => x"fffc2911",
			2606 => x"001e2911",
			2607 => x"ffa32911",
			2608 => x"0f005008",
			2609 => x"05002d04",
			2610 => x"00a52911",
			2611 => x"fff52911",
			2612 => x"0200ac0c",
			2613 => x"0f005508",
			2614 => x"00009404",
			2615 => x"ffc12911",
			2616 => x"004f2911",
			2617 => x"ff862911",
			2618 => x"0400660c",
			2619 => x"0200b908",
			2620 => x"0000b804",
			2621 => x"000d2911",
			2622 => x"fffb2911",
			2623 => x"00912911",
			2624 => x"fff82911",
			2625 => x"0d002504",
			2626 => x"ff9b2911",
			2627 => x"000f2911",
			2628 => x"0f007334",
			2629 => x"00006e0c",
			2630 => x"08001604",
			2631 => x"006a297d",
			2632 => x"04000704",
			2633 => x"001a297d",
			2634 => x"ff4d297d",
			2635 => x"05004518",
			2636 => x"0f006610",
			2637 => x"01000904",
			2638 => x"00e6297d",
			2639 => x"00009408",
			2640 => x"05001804",
			2641 => x"0068297d",
			2642 => x"ff64297d",
			2643 => x"0093297d",
			2644 => x"06006304",
			2645 => x"ffe2297d",
			2646 => x"003a297d",
			2647 => x"0200d008",
			2648 => x"08001804",
			2649 => x"fffe297d",
			2650 => x"ff6b297d",
			2651 => x"01001004",
			2652 => x"fff8297d",
			2653 => x"0069297d",
			2654 => x"ff59297d",
			2655 => x"06006c30",
			2656 => x"0200bb28",
			2657 => x"0f00551c",
			2658 => x"00007510",
			2659 => x"0f003c0c",
			2660 => x"02004604",
			2661 => x"ffd429e1",
			2662 => x"09001b04",
			2663 => x"006c29e1",
			2664 => x"ffe929e1",
			2665 => x"ff9429e1",
			2666 => x"03002d08",
			2667 => x"08002004",
			2668 => x"009129e1",
			2669 => x"fffd29e1",
			2670 => x"ffdb29e1",
			2671 => x"0200ac04",
			2672 => x"ff8f29e1",
			2673 => x"0d001304",
			2674 => x"001a29e1",
			2675 => x"ffe129e1",
			2676 => x"04006104",
			2677 => x"008b29e1",
			2678 => x"fff429e1",
			2679 => x"ffb029e1",
			2680 => x"0f007334",
			2681 => x"02006b0c",
			2682 => x"08001604",
			2683 => x"002b2a4d",
			2684 => x"04000504",
			2685 => x"00092a4d",
			2686 => x"ff6a2a4d",
			2687 => x"0400220c",
			2688 => x"06005304",
			2689 => x"00b32a4d",
			2690 => x"0200b504",
			2691 => x"ffb62a4d",
			2692 => x"004b2a4d",
			2693 => x"0200ac0c",
			2694 => x"04003c04",
			2695 => x"ff642a4d",
			2696 => x"0200a404",
			2697 => x"ffea2a4d",
			2698 => x"00142a4d",
			2699 => x"0400610c",
			2700 => x"0000c608",
			2701 => x"0f006a04",
			2702 => x"002a2a4d",
			2703 => x"ffdd2a4d",
			2704 => x"00b12a4d",
			2705 => x"ffe92a4d",
			2706 => x"ff702a4d",
			2707 => x"06006c34",
			2708 => x"02006b10",
			2709 => x"03001a0c",
			2710 => x"09001504",
			2711 => x"ffd32ab9",
			2712 => x"02004504",
			2713 => x"ffea2ab9",
			2714 => x"00602ab9",
			2715 => x"ffaa2ab9",
			2716 => x"0f005008",
			2717 => x"03002304",
			2718 => x"009f2ab9",
			2719 => x"fffb2ab9",
			2720 => x"0200a408",
			2721 => x"04001804",
			2722 => x"fff82ab9",
			2723 => x"ff8d2ab9",
			2724 => x"04005110",
			2725 => x"0200ac08",
			2726 => x"06005f04",
			2727 => x"00172ab9",
			2728 => x"ffec2ab9",
			2729 => x"06006804",
			2730 => x"008c2ab9",
			2731 => x"00032ab9",
			2732 => x"fff22ab9",
			2733 => x"ffac2ab9",
			2734 => x"0f007338",
			2735 => x"00007510",
			2736 => x"0f003c0c",
			2737 => x"02004604",
			2738 => x"ff952b2d",
			2739 => x"09001b04",
			2740 => x"00ce2b2d",
			2741 => x"ffc32b2d",
			2742 => x"ff252b2d",
			2743 => x"06004c0c",
			2744 => x"05002d08",
			2745 => x"08002004",
			2746 => x"011a2b2d",
			2747 => x"00162b2d",
			2748 => x"000f2b2d",
			2749 => x"0200ac0c",
			2750 => x"0f005808",
			2751 => x"02008c04",
			2752 => x"ff722b2d",
			2753 => x"007f2b2d",
			2754 => x"ff2d2b2d",
			2755 => x"0400610c",
			2756 => x"0200bc08",
			2757 => x"0f006604",
			2758 => x"009c2b2d",
			2759 => x"ff942b2d",
			2760 => x"00f62b2d",
			2761 => x"ffde2b2d",
			2762 => x"ff2a2b2d",
			2763 => x"06006c30",
			2764 => x"02004604",
			2765 => x"ffdf2b91",
			2766 => x"05002f14",
			2767 => x"06004e0c",
			2768 => x"00006e08",
			2769 => x"0b001504",
			2770 => x"001d2b91",
			2771 => x"ffef2b91",
			2772 => x"00802b91",
			2773 => x"00009504",
			2774 => x"ffc92b91",
			2775 => x"00342b91",
			2776 => x"0000c610",
			2777 => x"0800190c",
			2778 => x"0000ab04",
			2779 => x"ffee2b91",
			2780 => x"01000604",
			2781 => x"001c2b91",
			2782 => x"fff92b91",
			2783 => x"ffa72b91",
			2784 => x"04006104",
			2785 => x"00602b91",
			2786 => x"fff72b91",
			2787 => x"ffca2b91",
			2788 => x"0600673c",
			2789 => x"02005008",
			2790 => x"01000404",
			2791 => x"ffeb2c1d",
			2792 => x"fe552c1d",
			2793 => x"05004024",
			2794 => x"02008b10",
			2795 => x"05001b08",
			2796 => x"06003e04",
			2797 => x"033e2c1d",
			2798 => x"01d62c1d",
			2799 => x"01000704",
			2800 => x"01402c1d",
			2801 => x"fe4c2c1d",
			2802 => x"0f005a08",
			2803 => x"0200a004",
			2804 => x"03822c1d",
			2805 => x"030d2c1d",
			2806 => x"0000ba04",
			2807 => x"fe412c1d",
			2808 => x"0f006204",
			2809 => x"03072c1d",
			2810 => x"03c92c1d",
			2811 => x"0000c60c",
			2812 => x"01000608",
			2813 => x"06005d04",
			2814 => x"00d02c1d",
			2815 => x"fe5d2c1d",
			2816 => x"fe552c1d",
			2817 => x"03aa2c1d",
			2818 => x"0d002504",
			2819 => x"fe542c1d",
			2820 => x"09003304",
			2821 => x"00562c1d",
			2822 => x"fe642c1d",
			2823 => x"0f007338",
			2824 => x"0200bb30",
			2825 => x"0500211c",
			2826 => x"02006e14",
			2827 => x"07001908",
			2828 => x"02003804",
			2829 => x"ffde2c91",
			2830 => x"005a2c91",
			2831 => x"0a001408",
			2832 => x"05001504",
			2833 => x"ffc62c91",
			2834 => x"00482c91",
			2835 => x"ff982c91",
			2836 => x"06004e04",
			2837 => x"00bc2c91",
			2838 => x"ffe22c91",
			2839 => x"0100080c",
			2840 => x"0f006108",
			2841 => x"00008b04",
			2842 => x"ffc92c91",
			2843 => x"006a2c91",
			2844 => x"ffb72c91",
			2845 => x"0200b704",
			2846 => x"ff6a2c91",
			2847 => x"fffe2c91",
			2848 => x"04006104",
			2849 => x"00b52c91",
			2850 => x"ffef2c91",
			2851 => x"ff872c91",
			2852 => x"06006c40",
			2853 => x"02007114",
			2854 => x"0f004010",
			2855 => x"08001908",
			2856 => x"02004604",
			2857 => x"ffd52d15",
			2858 => x"00ac2d15",
			2859 => x"02005904",
			2860 => x"ffa62d15",
			2861 => x"00192d15",
			2862 => x"ff592d15",
			2863 => x"04002310",
			2864 => x"0f005404",
			2865 => x"00e12d15",
			2866 => x"0b001808",
			2867 => x"0b001404",
			2868 => x"000a2d15",
			2869 => x"ffba2d15",
			2870 => x"00682d15",
			2871 => x"0200ac0c",
			2872 => x"04003c04",
			2873 => x"ff5b2d15",
			2874 => x"0200a404",
			2875 => x"ffe92d15",
			2876 => x"00162d15",
			2877 => x"0400610c",
			2878 => x"0000c608",
			2879 => x"0f006a04",
			2880 => x"002d2d15",
			2881 => x"ffdc2d15",
			2882 => x"00b62d15",
			2883 => x"ffea2d15",
			2884 => x"ff6a2d15",
			2885 => x"0f007334",
			2886 => x"02004604",
			2887 => x"fe872d81",
			2888 => x"0500321c",
			2889 => x"06004e10",
			2890 => x"0200710c",
			2891 => x"03001a04",
			2892 => x"019f2d81",
			2893 => x"05002c04",
			2894 => x"fe822d81",
			2895 => x"007a2d81",
			2896 => x"019e2d81",
			2897 => x"02009004",
			2898 => x"fe882d81",
			2899 => x"01000604",
			2900 => x"00022d81",
			2901 => x"01732d81",
			2902 => x"0000c60c",
			2903 => x"0e005208",
			2904 => x"00009e04",
			2905 => x"fe8a2d81",
			2906 => x"011b2d81",
			2907 => x"fe792d81",
			2908 => x"04006104",
			2909 => x"01922d81",
			2910 => x"fed02d81",
			2911 => x"fe6e2d81",
			2912 => x"06006840",
			2913 => x"02005008",
			2914 => x"01000404",
			2915 => x"ffcc2e15",
			2916 => x"fe522e15",
			2917 => x"05003e28",
			2918 => x"02008210",
			2919 => x"03001708",
			2920 => x"01000704",
			2921 => x"046c2e15",
			2922 => x"031b2e15",
			2923 => x"08001b04",
			2924 => x"00df2e15",
			2925 => x"fe4c2e15",
			2926 => x"0f00570c",
			2927 => x"0000a108",
			2928 => x"04001204",
			2929 => x"03c62e15",
			2930 => x"055d2e15",
			2931 => x"03a82e15",
			2932 => x"0000b804",
			2933 => x"fe3e2e15",
			2934 => x"0b001504",
			2935 => x"04a82e15",
			2936 => x"03a72e15",
			2937 => x"0200ca0c",
			2938 => x"01000404",
			2939 => x"00942e15",
			2940 => x"0f005704",
			2941 => x"ffdf2e15",
			2942 => x"fe4f2e15",
			2943 => x"03872e15",
			2944 => x"0d002504",
			2945 => x"fe522e15",
			2946 => x"0d002704",
			2947 => x"00382e15",
			2948 => x"fe622e15",
			2949 => x"0f007330",
			2950 => x"02005004",
			2951 => x"fe672e79",
			2952 => x"05004824",
			2953 => x"0200820c",
			2954 => x"05002108",
			2955 => x"0a001604",
			2956 => x"01912e79",
			2957 => x"005f2e79",
			2958 => x"fe592e79",
			2959 => x"0f005508",
			2960 => x"07002604",
			2961 => x"01ad2e79",
			2962 => x"020e2e79",
			2963 => x"0000af08",
			2964 => x"06005304",
			2965 => x"ffaf2e79",
			2966 => x"fe652e79",
			2967 => x"0200bb04",
			2968 => x"01542e79",
			2969 => x"01de2e79",
			2970 => x"01001104",
			2971 => x"fe642e79",
			2972 => x"021a2e79",
			2973 => x"fe632e79",
			2974 => x"0f007340",
			2975 => x"01000510",
			2976 => x"03003a0c",
			2977 => x"04001408",
			2978 => x"07002104",
			2979 => x"00882efd",
			2980 => x"ff6a2efd",
			2981 => x"01282efd",
			2982 => x"ffa12efd",
			2983 => x"00008b14",
			2984 => x"05001b10",
			2985 => x"08001804",
			2986 => x"00b52efd",
			2987 => x"0c001404",
			2988 => x"ff1b2efd",
			2989 => x"09002004",
			2990 => x"00992efd",
			2991 => x"ff9d2efd",
			2992 => x"fed82efd",
			2993 => x"05003208",
			2994 => x"0b001504",
			2995 => x"00032efd",
			2996 => x"012c2efd",
			2997 => x"0000cc0c",
			2998 => x"08001804",
			2999 => x"004e2efd",
			3000 => x"0d001a04",
			3001 => x"fee42efd",
			3002 => x"ffe82efd",
			3003 => x"04006104",
			3004 => x"01002efd",
			3005 => x"ffb92efd",
			3006 => x"fecc2efd",
			3007 => x"0f007328",
			3008 => x"02005004",
			3009 => x"fe6f2f51",
			3010 => x"0a001604",
			3011 => x"01b62f51",
			3012 => x"02006e04",
			3013 => x"fe642f51",
			3014 => x"06004c0c",
			3015 => x"05002d08",
			3016 => x"01000c04",
			3017 => x"01fa2f51",
			3018 => x"01502f51",
			3019 => x"00762f51",
			3020 => x"0200a508",
			3021 => x"0f005704",
			3022 => x"ffe42f51",
			3023 => x"fe6a2f51",
			3024 => x"04005104",
			3025 => x"01632f51",
			3026 => x"fe952f51",
			3027 => x"fe672f51",
			3028 => x"06006840",
			3029 => x"02005008",
			3030 => x"05002004",
			3031 => x"fe5d2fe5",
			3032 => x"001f2fe5",
			3033 => x"05004830",
			3034 => x"02009a1c",
			3035 => x"0500210c",
			3036 => x"06004d08",
			3037 => x"00007204",
			3038 => x"01962fe5",
			3039 => x"02862fe5",
			3040 => x"ffd12fe5",
			3041 => x"09002008",
			3042 => x"0f003f04",
			3043 => x"00032fe5",
			3044 => x"fe4c2fe5",
			3045 => x"04002704",
			3046 => x"01d62fe5",
			3047 => x"fe672fe5",
			3048 => x"0200a508",
			3049 => x"06005004",
			3050 => x"02572fe5",
			3051 => x"ffe32fe5",
			3052 => x"0d001304",
			3053 => x"02b42fe5",
			3054 => x"0200b004",
			3055 => x"01f62fe5",
			3056 => x"024e2fe5",
			3057 => x"01001004",
			3058 => x"fe5a2fe5",
			3059 => x"01942fe5",
			3060 => x"0d002504",
			3061 => x"fe5b2fe5",
			3062 => x"0d002704",
			3063 => x"00d32fe5",
			3064 => x"fe702fe5",
			3065 => x"0f007330",
			3066 => x"0200bb28",
			3067 => x"0f006124",
			3068 => x"02009820",
			3069 => x"0f004210",
			3070 => x"01000708",
			3071 => x"00004904",
			3072 => x"ff893049",
			3073 => x"01763049",
			3074 => x"05001604",
			3075 => x"00813049",
			3076 => x"fef03049",
			3077 => x"00008308",
			3078 => x"01000e04",
			3079 => x"fe9a3049",
			3080 => x"ffa53049",
			3081 => x"04002204",
			3082 => x"00de3049",
			3083 => x"fedc3049",
			3084 => x"015b3049",
			3085 => x"feba3049",
			3086 => x"03005c04",
			3087 => x"015e3049",
			3088 => x"ff7d3049",
			3089 => x"fe913049",
			3090 => x"0f00733c",
			3091 => x"08001504",
			3092 => x"00d630c5",
			3093 => x"00006e10",
			3094 => x"03000c08",
			3095 => x"05000d04",
			3096 => x"fff030c5",
			3097 => x"002a30c5",
			3098 => x"08001804",
			3099 => x"000330c5",
			3100 => x"ff4f30c5",
			3101 => x"04002214",
			3102 => x"0b001404",
			3103 => x"ffd030c5",
			3104 => x"06005308",
			3105 => x"01000f04",
			3106 => x"00db30c5",
			3107 => x"000730c5",
			3108 => x"0d001604",
			3109 => x"ffe030c5",
			3110 => x"002c30c5",
			3111 => x"0200a508",
			3112 => x"03002d04",
			3113 => x"fffc30c5",
			3114 => x"ff5b30c5",
			3115 => x"0f006604",
			3116 => x"00a130c5",
			3117 => x"0200d504",
			3118 => x"ff7a30c5",
			3119 => x"006630c5",
			3120 => x"ff5230c5",
			3121 => x"0f007334",
			3122 => x"02004604",
			3123 => x"fe743131",
			3124 => x"0d000e04",
			3125 => x"021e3131",
			3126 => x"02006b10",
			3127 => x"06003308",
			3128 => x"04001204",
			3129 => x"00e93131",
			3130 => x"feb33131",
			3131 => x"0c001504",
			3132 => x"fd9a3131",
			3133 => x"fe983131",
			3134 => x"06004c0c",
			3135 => x"05002d08",
			3136 => x"01000904",
			3137 => x"01f93131",
			3138 => x"01483131",
			3139 => x"00523131",
			3140 => x"0200a408",
			3141 => x"04001804",
			3142 => x"ffd13131",
			3143 => x"fe6b3131",
			3144 => x"0f006604",
			3145 => x"01ab3131",
			3146 => x"00383131",
			3147 => x"fe683131",
			3148 => x"0f007334",
			3149 => x"02004604",
			3150 => x"fe67319f",
			3151 => x"0a00652c",
			3152 => x"0200bb20",
			3153 => x"0f005510",
			3154 => x"02007108",
			3155 => x"08001804",
			3156 => x"01ec319f",
			3157 => x"ff1d319f",
			3158 => x"04002504",
			3159 => x"01ef319f",
			3160 => x"0005319f",
			3161 => x"0200ac08",
			3162 => x"0f005904",
			3163 => x"ff80319f",
			3164 => x"fe5a319f",
			3165 => x"0a003d04",
			3166 => x"019f319f",
			3167 => x"fe7b319f",
			3168 => x"0000e608",
			3169 => x"0e005c04",
			3170 => x"01e1319f",
			3171 => x"003f319f",
			3172 => x"0267319f",
			3173 => x"fe69319f",
			3174 => x"fe62319f",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1063, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2143, initial_addr_3'length));
	end generate gen_rom_9;

	gen_rom_10: if SELECT_ROM = 10 generate
		bank <= (
			0 => x"0b001f04",
			1 => x"ffce001d",
			2 => x"04002004",
			3 => x"ffe6001d",
			4 => x"0f009304",
			5 => x"005d001d",
			6 => x"fff9001d",
			7 => x"0a005c0c",
			8 => x"0c002504",
			9 => x"ff9e0041",
			10 => x"0a004304",
			11 => x"fff40041",
			12 => x"00210041",
			13 => x"04006104",
			14 => x"00020041",
			15 => x"004a0041",
			16 => x"03006110",
			17 => x"0f004808",
			18 => x"0a002d04",
			19 => x"ff9b0065",
			20 => x"00960065",
			21 => x"0c002a04",
			22 => x"fee70065",
			23 => x"00270065",
			24 => x"00e50065",
			25 => x"0c001f04",
			26 => x"ff550089",
			27 => x"0200da08",
			28 => x"04002004",
			29 => x"ffc30089",
			30 => x"00ba0089",
			31 => x"03006104",
			32 => x"ff840089",
			33 => x"005a0089",
			34 => x"0c001f04",
			35 => x"ff8900ad",
			36 => x"0200da08",
			37 => x"03003504",
			38 => x"ffe800ad",
			39 => x"008e00ad",
			40 => x"03006104",
			41 => x"ffa800ad",
			42 => x"004300ad",
			43 => x"03006110",
			44 => x"0f004808",
			45 => x"0a002f04",
			46 => x"ffe100d1",
			47 => x"004900d1",
			48 => x"0c002a04",
			49 => x"ff7500d1",
			50 => x"001200d1",
			51 => x"006900d1",
			52 => x"0a005c10",
			53 => x"0f004108",
			54 => x"03002c04",
			55 => x"ffe900f5",
			56 => x"003c00f5",
			57 => x"0c002a04",
			58 => x"ff8400f5",
			59 => x"000900f5",
			60 => x"005500f5",
			61 => x"03004004",
			62 => x"ff9d0119",
			63 => x"0200da08",
			64 => x"0b001d04",
			65 => x"fff90119",
			66 => x"00600119",
			67 => x"03006104",
			68 => x"ffca0119",
			69 => x"00280119",
			70 => x"03003504",
			71 => x"ffd0013d",
			72 => x"0200da08",
			73 => x"0b001d04",
			74 => x"fff4013d",
			75 => x"004d013d",
			76 => x"03006104",
			77 => x"ffd6013d",
			78 => x"001e013d",
			79 => x"05008110",
			80 => x"0f004108",
			81 => x"04002004",
			82 => x"fff40161",
			83 => x"00280161",
			84 => x"0c002a04",
			85 => x"ffb60161",
			86 => x"000c0161",
			87 => x"00370161",
			88 => x"0a005c10",
			89 => x"0f004808",
			90 => x"0a002f04",
			91 => x"ff6f018d",
			92 => x"00ca018d",
			93 => x"0c002a04",
			94 => x"febc018d",
			95 => x"0014018d",
			96 => x"0d002204",
			97 => x"0108018d",
			98 => x"001e018d",
			99 => x"0a005c10",
			100 => x"02006808",
			101 => x"0a002c04",
			102 => x"ffb601b9",
			103 => x"007401b9",
			104 => x"0c002a04",
			105 => x"ff1001b9",
			106 => x"000101b9",
			107 => x"04006104",
			108 => x"000a01b9",
			109 => x"00bb01b9",
			110 => x"0a005c10",
			111 => x"0c002504",
			112 => x"fe6b01dd",
			113 => x"0000e508",
			114 => x"04001a04",
			115 => x"ff2001dd",
			116 => x"00fa01dd",
			117 => x"feb801dd",
			118 => x"019101dd",
			119 => x"0a005c10",
			120 => x"0b002004",
			121 => x"fecf0201",
			122 => x"0000d308",
			123 => x"0a002f04",
			124 => x"ffc90201",
			125 => x"009e0201",
			126 => x"ff840201",
			127 => x"00fa0201",
			128 => x"03003504",
			129 => x"ff740225",
			130 => x"0c001f04",
			131 => x"ffcf0225",
			132 => x"0200da04",
			133 => x"008c0225",
			134 => x"03006104",
			135 => x"ffa70225",
			136 => x"00470225",
			137 => x"03003504",
			138 => x"ffa20249",
			139 => x"0c001f04",
			140 => x"ffe50249",
			141 => x"0200f204",
			142 => x"00740249",
			143 => x"01001404",
			144 => x"000f0249",
			145 => x"ffe50249",
			146 => x"03003504",
			147 => x"ffc6026d",
			148 => x"0c001f04",
			149 => x"ffed026d",
			150 => x"0200f204",
			151 => x"0057026d",
			152 => x"01001404",
			153 => x"000d026d",
			154 => x"ffed026d",
			155 => x"0a005c10",
			156 => x"0b002004",
			157 => x"fe610299",
			158 => x"03003504",
			159 => x"fe6e0299",
			160 => x"0200dc04",
			161 => x"02880299",
			162 => x"fe540299",
			163 => x"0200f204",
			164 => x"01b10299",
			165 => x"00f20299",
			166 => x"0b001f08",
			167 => x"04005004",
			168 => x"feaa02c5",
			169 => x"ffca02c5",
			170 => x"03003504",
			171 => x"ff5702c5",
			172 => x"0200e404",
			173 => x"012502c5",
			174 => x"03006104",
			175 => x"ff4802c5",
			176 => x"00b802c5",
			177 => x"0b001f08",
			178 => x"0c002204",
			179 => x"ffb102f1",
			180 => x"000302f1",
			181 => x"04002004",
			182 => x"ffdf02f1",
			183 => x"0200f204",
			184 => x"006402f1",
			185 => x"03006e04",
			186 => x"ffe302f1",
			187 => x"001402f1",
			188 => x"0a00480c",
			189 => x"03004004",
			190 => x"ff180325",
			191 => x"0a004704",
			192 => x"00070325",
			193 => x"ffef0325",
			194 => x"0200da08",
			195 => x"0b001d04",
			196 => x"ffea0325",
			197 => x"00ba0325",
			198 => x"03006104",
			199 => x"ff860325",
			200 => x"006c0325",
			201 => x"05008114",
			202 => x"0f004808",
			203 => x"0a002f04",
			204 => x"ffe20351",
			205 => x"00480351",
			206 => x"0c002a04",
			207 => x"ff710351",
			208 => x"0a004804",
			209 => x"fff60351",
			210 => x"00260351",
			211 => x"00670351",
			212 => x"03005014",
			213 => x"0b00240c",
			214 => x"0b002004",
			215 => x"fe500385",
			216 => x"0b002104",
			217 => x"fe9c0385",
			218 => x"fe540385",
			219 => x"03003504",
			220 => x"fe530385",
			221 => x"02860385",
			222 => x"03006104",
			223 => x"028c0385",
			224 => x"03980385",
			225 => x"03005014",
			226 => x"0b00240c",
			227 => x"0b002004",
			228 => x"fe5c03b9",
			229 => x"09002804",
			230 => x"014903b9",
			231 => x"fe6103b9",
			232 => x"03003804",
			233 => x"fe6203b9",
			234 => x"022303b9",
			235 => x"03006104",
			236 => x"00b703b9",
			237 => x"021e03b9",
			238 => x"03005014",
			239 => x"0b00240c",
			240 => x"0b002004",
			241 => x"fe4d03f5",
			242 => x"0b002104",
			243 => x"fe8f03f5",
			244 => x"fe5003f5",
			245 => x"0a003d04",
			246 => x"fe4f03f5",
			247 => x"02f603f5",
			248 => x"0000c504",
			249 => x"05c503f5",
			250 => x"04006104",
			251 => x"00c603f5",
			252 => x"048603f5",
			253 => x"0c001f04",
			254 => x"fe8d0421",
			255 => x"03006110",
			256 => x"0000cc08",
			257 => x"04001f04",
			258 => x"ff320421",
			259 => x"01540421",
			260 => x"0b002804",
			261 => x"fec70421",
			262 => x"fff40421",
			263 => x"01520421",
			264 => x"05008114",
			265 => x"0b002004",
			266 => x"fea3044d",
			267 => x"0000d308",
			268 => x"03003504",
			269 => x"ff9e044d",
			270 => x"00cb044d",
			271 => x"0c002a04",
			272 => x"ff39044d",
			273 => x"000b044d",
			274 => x"0124044d",
			275 => x"03003504",
			276 => x"ff490479",
			277 => x"0c001f04",
			278 => x"ffbb0479",
			279 => x"0f008508",
			280 => x"0200e404",
			281 => x"00b20479",
			282 => x"00070479",
			283 => x"03006104",
			284 => x"ffbc0479",
			285 => x"00390479",
			286 => x"0a006518",
			287 => x"0b002008",
			288 => x"04005004",
			289 => x"fe6604ad",
			290 => x"ff4e04ad",
			291 => x"0000d308",
			292 => x"04001e04",
			293 => x"fe7f04ad",
			294 => x"023604ad",
			295 => x"08002904",
			296 => x"ff9404ad",
			297 => x"fe4d04ad",
			298 => x"01a404ad",
			299 => x"0b001f08",
			300 => x"04005004",
			301 => x"fe8904e1",
			302 => x"fff404e1",
			303 => x"03003504",
			304 => x"ff1b04e1",
			305 => x"0f00930c",
			306 => x"01001104",
			307 => x"016904e1",
			308 => x"0000db04",
			309 => x"00c704e1",
			310 => x"fff604e1",
			311 => x"ff9804e1",
			312 => x"03003504",
			313 => x"ff6e0515",
			314 => x"0b001f0c",
			315 => x"06006908",
			316 => x"03004504",
			317 => x"ffec0515",
			318 => x"002d0515",
			319 => x"ffc20515",
			320 => x"0200f204",
			321 => x"00880515",
			322 => x"01001604",
			323 => x"00180515",
			324 => x"ffd60515",
			325 => x"0a005c14",
			326 => x"03005010",
			327 => x"0b00280c",
			328 => x"0a004a04",
			329 => x"d5e80541",
			330 => x"0000ca04",
			331 => x"d7440541",
			332 => x"d5ea0541",
			333 => x"d7b30541",
			334 => x"da9a0541",
			335 => x"eb810541",
			336 => x"03005018",
			337 => x"0b002814",
			338 => x"0a004a0c",
			339 => x"0b002004",
			340 => x"fe53057d",
			341 => x"07002d04",
			342 => x"002e057d",
			343 => x"fe55057d",
			344 => x"0000cb04",
			345 => x"0068057d",
			346 => x"fe5b057d",
			347 => x"003d057d",
			348 => x"0a006504",
			349 => x"01c5057d",
			350 => x"030c057d",
			351 => x"0b001f08",
			352 => x"05006804",
			353 => x"fe6b05b9",
			354 => x"000405b9",
			355 => x"03003504",
			356 => x"fe9005b9",
			357 => x"0200f20c",
			358 => x"0000c504",
			359 => x"021d05b9",
			360 => x"06006704",
			361 => x"004705b9",
			362 => x"018d05b9",
			363 => x"03007a04",
			364 => x"fe7e05b9",
			365 => x"016005b9",
			366 => x"0a004814",
			367 => x"0300400c",
			368 => x"03003504",
			369 => x"fe60060d",
			370 => x"07002604",
			371 => x"02a2060d",
			372 => x"fe62060d",
			373 => x"0e005d04",
			374 => x"014b060d",
			375 => x"fe7f060d",
			376 => x"0b001f08",
			377 => x"0f007204",
			378 => x"0070060d",
			379 => x"fe3a060d",
			380 => x"0200e408",
			381 => x"0a006e04",
			382 => x"02cc060d",
			383 => x"01da060d",
			384 => x"03007304",
			385 => x"ff81060d",
			386 => x"01df060d",
			387 => x"0300611c",
			388 => x"0b002008",
			389 => x"0c002204",
			390 => x"fe7f0649",
			391 => x"ffdb0649",
			392 => x"01001108",
			393 => x"04001a04",
			394 => x"ffb00649",
			395 => x"01660649",
			396 => x"0c002a04",
			397 => x"fec40649",
			398 => x"0a003904",
			399 => x"ffb50649",
			400 => x"00960649",
			401 => x"016c0649",
			402 => x"03003504",
			403 => x"ffb1067d",
			404 => x"0c001f04",
			405 => x"ffe6067d",
			406 => x"0200da04",
			407 => x"0060067d",
			408 => x"06007d08",
			409 => x"08002204",
			410 => x"0008067d",
			411 => x"ffe3067d",
			412 => x"0f009304",
			413 => x"0015067d",
			414 => x"fff9067d",
			415 => x"0b001e0c",
			416 => x"0b001d04",
			417 => x"fe7006c9",
			418 => x"05003a04",
			419 => x"ff6e06c9",
			420 => x"001d06c9",
			421 => x"03003504",
			422 => x"fe9e06c9",
			423 => x"0200f210",
			424 => x"01001108",
			425 => x"06007804",
			426 => x"01dc06c9",
			427 => x"00b106c9",
			428 => x"0c002a04",
			429 => x"fff506c9",
			430 => x"015e06c9",
			431 => x"03006e04",
			432 => x"fe9306c9",
			433 => x"013a06c9",
			434 => x"0c001f04",
			435 => x"fe98071f",
			436 => x"0100110c",
			437 => x"03003504",
			438 => x"ffa9071f",
			439 => x"0f008a04",
			440 => x"0155071f",
			441 => x"ffef071f",
			442 => x"0c002a14",
			443 => x"0800270c",
			444 => x"09002904",
			445 => x"ffaa071f",
			446 => x"00005c04",
			447 => x"ffe6071f",
			448 => x"0057071f",
			449 => x"09003104",
			450 => x"fef4071f",
			451 => x"fffc071f",
			452 => x"03004504",
			453 => x"ffba071f",
			454 => x"00eb071f",
			455 => x"0b001f04",
			456 => x"ffcf0739",
			457 => x"04002004",
			458 => x"ffe60739",
			459 => x"0f009304",
			460 => x"005a0739",
			461 => x"fff90739",
			462 => x"0a005c0c",
			463 => x"0c002504",
			464 => x"ffa1075d",
			465 => x"0a004304",
			466 => x"fff4075d",
			467 => x"0021075d",
			468 => x"04006104",
			469 => x"0002075d",
			470 => x"0049075d",
			471 => x"03006110",
			472 => x"02006808",
			473 => x"0a002c04",
			474 => x"ffb30781",
			475 => x"00780781",
			476 => x"0c002a04",
			477 => x"ff0d0781",
			478 => x"00170781",
			479 => x"00c60781",
			480 => x"0c001f04",
			481 => x"ff5d07a5",
			482 => x"0200da08",
			483 => x"04002004",
			484 => x"ffc507a5",
			485 => x"00b307a5",
			486 => x"03006104",
			487 => x"ff8907a5",
			488 => x"005807a5",
			489 => x"0a005c10",
			490 => x"0f004808",
			491 => x"03002c04",
			492 => x"ffdd07c9",
			493 => x"004d07c9",
			494 => x"0c002a04",
			495 => x"ff6907c9",
			496 => x"000a07c9",
			497 => x"007607c9",
			498 => x"05008110",
			499 => x"0f004808",
			500 => x"0a002d04",
			501 => x"ffe207ed",
			502 => x"004807ed",
			503 => x"0c002a04",
			504 => x"ff7807ed",
			505 => x"001107ed",
			506 => x"006607ed",
			507 => x"05008110",
			508 => x"0f004108",
			509 => x"03002c04",
			510 => x"ffe90811",
			511 => x"003b0811",
			512 => x"0c002a04",
			513 => x"ff810811",
			514 => x"00180811",
			515 => x"00580811",
			516 => x"03006110",
			517 => x"0f004808",
			518 => x"05002e04",
			519 => x"ffef0835",
			520 => x"00320835",
			521 => x"0c002a04",
			522 => x"ffaa0835",
			523 => x"000b0835",
			524 => x"00420835",
			525 => x"03003504",
			526 => x"ffd10859",
			527 => x"0200da08",
			528 => x"0b001d04",
			529 => x"fff40859",
			530 => x"004b0859",
			531 => x"03006104",
			532 => x"ffd70859",
			533 => x"001d0859",
			534 => x"05008110",
			535 => x"0f004808",
			536 => x"05002e04",
			537 => x"fff4087d",
			538 => x"002a087d",
			539 => x"0c002a04",
			540 => x"ffb9087d",
			541 => x"0008087d",
			542 => x"0037087d",
			543 => x"0a005c10",
			544 => x"02005808",
			545 => x"0a002c04",
			546 => x"ff9208a9",
			547 => x"00ab08a9",
			548 => x"0c002a04",
			549 => x"fec008a9",
			550 => x"002408a9",
			551 => x"01001404",
			552 => x"00fb08a9",
			553 => x"001608a9",
			554 => x"0a005c10",
			555 => x"02007108",
			556 => x"03002c04",
			557 => x"ffd308d5",
			558 => x"006608d5",
			559 => x"0c002a04",
			560 => x"ff4b08d5",
			561 => x"000a08d5",
			562 => x"01001604",
			563 => x"008408d5",
			564 => x"000108d5",
			565 => x"0c001f04",
			566 => x"fe7908f9",
			567 => x"03003504",
			568 => x"fec908f9",
			569 => x"0200da04",
			570 => x"018b08f9",
			571 => x"03006104",
			572 => x"fea208f9",
			573 => x"015908f9",
			574 => x"0c001f04",
			575 => x"ff07091d",
			576 => x"03003504",
			577 => x"ff98091d",
			578 => x"0200f204",
			579 => x"00c9091d",
			580 => x"03006e04",
			581 => x"ffa2091d",
			582 => x"003c091d",
			583 => x"05008110",
			584 => x"0b002004",
			585 => x"ff5f0941",
			586 => x"0000df08",
			587 => x"03003504",
			588 => x"ffe40941",
			589 => x"00610941",
			590 => x"ffcd0941",
			591 => x"00800941",
			592 => x"03003504",
			593 => x"ffa50965",
			594 => x"0c001f04",
			595 => x"ffe50965",
			596 => x"0200f204",
			597 => x"00700965",
			598 => x"01001404",
			599 => x"000f0965",
			600 => x"ffe60965",
			601 => x"0a006510",
			602 => x"0200ba0c",
			603 => x"03003504",
			604 => x"ffe70989",
			605 => x"0c001d04",
			606 => x"fff90989",
			607 => x"00300989",
			608 => x"ffba0989",
			609 => x"003a0989",
			610 => x"0a005c10",
			611 => x"0b002004",
			612 => x"fe6209b5",
			613 => x"03003504",
			614 => x"fe7009b5",
			615 => x"0200dc04",
			616 => x"025709b5",
			617 => x"fe5c09b5",
			618 => x"05008104",
			619 => x"00d709b5",
			620 => x"01ab09b5",
			621 => x"0b001f08",
			622 => x"04005004",
			623 => x"ff3609e1",
			624 => x"ffe809e1",
			625 => x"04002004",
			626 => x"ffc509e1",
			627 => x"0200f204",
			628 => x"00ba09e1",
			629 => x"03006e04",
			630 => x"ffb309e1",
			631 => x"003009e1",
			632 => x"0b001f08",
			633 => x"0c002204",
			634 => x"ffb30a0d",
			635 => x"00030a0d",
			636 => x"04002004",
			637 => x"ffe00a0d",
			638 => x"0200f204",
			639 => x"00610a0d",
			640 => x"03006e04",
			641 => x"ffe40a0d",
			642 => x"00140a0d",
			643 => x"0a00480c",
			644 => x"07002408",
			645 => x"03003304",
			646 => x"fff70a41",
			647 => x"00220a41",
			648 => x"ffb50a41",
			649 => x"0200da08",
			650 => x"0b001d04",
			651 => x"fffb0a41",
			652 => x"004a0a41",
			653 => x"03006104",
			654 => x"ffd70a41",
			655 => x"00230a41",
			656 => x"05008114",
			657 => x"0f004808",
			658 => x"05002e04",
			659 => x"fff30a6d",
			660 => x"00290a6d",
			661 => x"0c002a04",
			662 => x"ffb10a6d",
			663 => x"0c002f04",
			664 => x"00000a6d",
			665 => x"000b0a6d",
			666 => x"003b0a6d",
			667 => x"03005014",
			668 => x"0b00240c",
			669 => x"0b002004",
			670 => x"fe580aa1",
			671 => x"07002d04",
			672 => x"00890aa1",
			673 => x"fe5c0aa1",
			674 => x"0a003e04",
			675 => x"fe5d0aa1",
			676 => x"03580aa1",
			677 => x"0a006504",
			678 => x"01370aa1",
			679 => x"026f0aa1",
			680 => x"03005014",
			681 => x"0300400c",
			682 => x"03003504",
			683 => x"fe5d0ad5",
			684 => x"00009b04",
			685 => x"01c60ad5",
			686 => x"fe5e0ad5",
			687 => x"0000be04",
			688 => x"03870ad5",
			689 => x"fe630ad5",
			690 => x"03006104",
			691 => x"009e0ad5",
			692 => x"02030ad5",
			693 => x"03005014",
			694 => x"0a00480c",
			695 => x"03003504",
			696 => x"fe560b11",
			697 => x"07002604",
			698 => x"00c80b11",
			699 => x"fe570b11",
			700 => x"0f007004",
			701 => x"03130b11",
			702 => x"fe5d0b11",
			703 => x"0a005c04",
			704 => x"01190b11",
			705 => x"01001604",
			706 => x"02ae0b11",
			707 => x"025b0b11",
			708 => x"0c001f04",
			709 => x"fe920b3d",
			710 => x"03006110",
			711 => x"0000cc08",
			712 => x"04001f04",
			713 => x"ff3f0b3d",
			714 => x"01470b3d",
			715 => x"0b002804",
			716 => x"fed20b3d",
			717 => x"fff40b3d",
			718 => x"014a0b3d",
			719 => x"05008114",
			720 => x"0b002004",
			721 => x"feaa0b69",
			722 => x"0000d308",
			723 => x"03003504",
			724 => x"ffa40b69",
			725 => x"00c20b69",
			726 => x"0c002a04",
			727 => x"ff450b69",
			728 => x"000b0b69",
			729 => x"011b0b69",
			730 => x"0a005c18",
			731 => x"0c00250c",
			732 => x"0b002004",
			733 => x"fe600ba5",
			734 => x"0c002104",
			735 => x"02090ba5",
			736 => x"fe6b0ba5",
			737 => x"0000e508",
			738 => x"03001d04",
			739 => x"fe880ba5",
			740 => x"021e0ba5",
			741 => x"fe470ba5",
			742 => x"01001604",
			743 => x"01bf0ba5",
			744 => x"011e0ba5",
			745 => x"0a006518",
			746 => x"0b002008",
			747 => x"0c002204",
			748 => x"fe680bd9",
			749 => x"00250bd9",
			750 => x"0000d308",
			751 => x"04001d04",
			752 => x"feab0bd9",
			753 => x"022a0bd9",
			754 => x"0d002004",
			755 => x"ffa40bd9",
			756 => x"fe700bd9",
			757 => x"01970bd9",
			758 => x"0a005c14",
			759 => x"0b002004",
			760 => x"fec70c0d",
			761 => x"07002d04",
			762 => x"009b0c0d",
			763 => x"0c002a08",
			764 => x"0d001c04",
			765 => x"00090c0d",
			766 => x"ff620c0d",
			767 => x"001e0c0d",
			768 => x"01001404",
			769 => x"00f20c0d",
			770 => x"00160c0d",
			771 => x"03003504",
			772 => x"ffba0c41",
			773 => x"0b001f0c",
			774 => x"06006908",
			775 => x"0200b804",
			776 => x"fff80c41",
			777 => x"00180c41",
			778 => x"ffdb0c41",
			779 => x"0200f204",
			780 => x"00500c41",
			781 => x"01001704",
			782 => x"00110c41",
			783 => x"ffec0c41",
			784 => x"0a00480c",
			785 => x"0b002004",
			786 => x"fe610c85",
			787 => x"07002d04",
			788 => x"02b20c85",
			789 => x"fe670c85",
			790 => x"0b001f08",
			791 => x"06006904",
			792 => x"00b80c85",
			793 => x"fe470c85",
			794 => x"0200e408",
			795 => x"0a006e04",
			796 => x"02610c85",
			797 => x"01c30c85",
			798 => x"04007704",
			799 => x"ff690c85",
			800 => x"01c40c85",
			801 => x"0b001f08",
			802 => x"04005004",
			803 => x"fe680cc1",
			804 => x"003c0cc1",
			805 => x"03003504",
			806 => x"fe7f0cc1",
			807 => x"0200f20c",
			808 => x"0c002304",
			809 => x"02a40cc1",
			810 => x"0200e404",
			811 => x"01990cc1",
			812 => x"00aa0cc1",
			813 => x"03006e04",
			814 => x"fe550cc1",
			815 => x"017d0cc1",
			816 => x"0b001f08",
			817 => x"05006804",
			818 => x"fe720cfd",
			819 => x"fff00cfd",
			820 => x"03003504",
			821 => x"febe0cfd",
			822 => x"01001308",
			823 => x"0200ec04",
			824 => x"01bf0cfd",
			825 => x"00cc0cfd",
			826 => x"0c002a08",
			827 => x"08002904",
			828 => x"fff50cfd",
			829 => x"feb60cfd",
			830 => x"01350cfd",
			831 => x"0a004814",
			832 => x"0a00450c",
			833 => x"03003504",
			834 => x"fe610d51",
			835 => x"00009b04",
			836 => x"01c70d51",
			837 => x"fe640d51",
			838 => x"04003b04",
			839 => x"01b30d51",
			840 => x"fe7f0d51",
			841 => x"0b001f08",
			842 => x"06006904",
			843 => x"00cd0d51",
			844 => x"fe410d51",
			845 => x"0200e408",
			846 => x"0a006e04",
			847 => x"02940d51",
			848 => x"01cd0d51",
			849 => x"03007304",
			850 => x"ff5f0d51",
			851 => x"01cf0d51",
			852 => x"0300611c",
			853 => x"0b002008",
			854 => x"0c002204",
			855 => x"fe830d8d",
			856 => x"ffe20d8d",
			857 => x"01001108",
			858 => x"04001a04",
			859 => x"ffb60d8d",
			860 => x"01510d8d",
			861 => x"0c002a04",
			862 => x"fecf0d8d",
			863 => x"0a003904",
			864 => x"ffb90d8d",
			865 => x"008e0d8d",
			866 => x"01650d8d",
			867 => x"03003504",
			868 => x"ffc60dc1",
			869 => x"0c001f04",
			870 => x"ffed0dc1",
			871 => x"0200da04",
			872 => x"00560dc1",
			873 => x"06007d08",
			874 => x"08002204",
			875 => x"00070dc1",
			876 => x"ffe80dc1",
			877 => x"0f009304",
			878 => x"00120dc1",
			879 => x"fff80dc1",
			880 => x"0b001f08",
			881 => x"05006804",
			882 => x"fe710e0f",
			883 => x"ffef0e0f",
			884 => x"01001108",
			885 => x"03003504",
			886 => x"ff2c0e0f",
			887 => x"01c00e0f",
			888 => x"0c002a10",
			889 => x"08002708",
			890 => x"03004404",
			891 => x"ff2c0e0f",
			892 => x"00bf0e0f",
			893 => x"09003104",
			894 => x"fe930e0f",
			895 => x"fffb0e0f",
			896 => x"03004504",
			897 => x"ff490e0f",
			898 => x"015b0e0f",
			899 => x"03003504",
			900 => x"ffd80e29",
			901 => x"0c001f04",
			902 => x"fff40e29",
			903 => x"0f009304",
			904 => x"00410e29",
			905 => x"fffb0e29",
			906 => x"03006110",
			907 => x"0f004808",
			908 => x"0a002f04",
			909 => x"ff660e4d",
			910 => x"00d60e4d",
			911 => x"0c002a04",
			912 => x"fec30e4d",
			913 => x"002a0e4d",
			914 => x"01140e4d",
			915 => x"0a005c10",
			916 => x"0f004808",
			917 => x"0a002f04",
			918 => x"ffc80e71",
			919 => x"00760e71",
			920 => x"0c002a04",
			921 => x"ff350e71",
			922 => x"000a0e71",
			923 => x"00aa0e71",
			924 => x"0c001f04",
			925 => x"ff840e95",
			926 => x"0200da08",
			927 => x"03003504",
			928 => x"ffe70e95",
			929 => x"00930e95",
			930 => x"03006104",
			931 => x"ffa50e95",
			932 => x"00440e95",
			933 => x"0a005c10",
			934 => x"0f004808",
			935 => x"03002c04",
			936 => x"ffde0eb9",
			937 => x"004b0eb9",
			938 => x"0c002a04",
			939 => x"ff6f0eb9",
			940 => x"000a0eb9",
			941 => x"00730eb9",
			942 => x"05008110",
			943 => x"0f004808",
			944 => x"0a002d04",
			945 => x"ffe30edd",
			946 => x"00470edd",
			947 => x"0c002a04",
			948 => x"ff7d0edd",
			949 => x"00110edd",
			950 => x"00630edd",
			951 => x"0a004504",
			952 => x"ff9a0f01",
			953 => x"0200da08",
			954 => x"0b001d04",
			955 => x"fff90f01",
			956 => x"00610f01",
			957 => x"03006104",
			958 => x"ffc90f01",
			959 => x"00290f01",
			960 => x"0a006510",
			961 => x"0f004808",
			962 => x"05002e04",
			963 => x"fff10f25",
			964 => x"00280f25",
			965 => x"0c002a04",
			966 => x"ffb30f25",
			967 => x"000a0f25",
			968 => x"003b0f25",
			969 => x"05008110",
			970 => x"0f004108",
			971 => x"03002c04",
			972 => x"fff40f49",
			973 => x"00280f49",
			974 => x"0c002a04",
			975 => x"ffb40f49",
			976 => x"000c0f49",
			977 => x"00380f49",
			978 => x"05008110",
			979 => x"0f004808",
			980 => x"05002e04",
			981 => x"fff50f6d",
			982 => x"00290f6d",
			983 => x"0c002a04",
			984 => x"ffbb0f6d",
			985 => x"00080f6d",
			986 => x"00370f6d",
			987 => x"0a005c10",
			988 => x"0f004808",
			989 => x"03002c04",
			990 => x"ff9f0f99",
			991 => x"008f0f99",
			992 => x"0c002a04",
			993 => x"fee60f99",
			994 => x"000e0f99",
			995 => x"0200f204",
			996 => x"00db0f99",
			997 => x"00080f99",
			998 => x"0a005c10",
			999 => x"0c002504",
			1000 => x"fe690fbd",
			1001 => x"0000e508",
			1002 => x"04001a04",
			1003 => x"ff120fbd",
			1004 => x"010b0fbd",
			1005 => x"feac0fbd",
			1006 => x"01940fbd",
			1007 => x"0c001f04",
			1008 => x"fe7c0fe1",
			1009 => x"03003504",
			1010 => x"fed40fe1",
			1011 => x"0200da04",
			1012 => x"017e0fe1",
			1013 => x"03006104",
			1014 => x"feab0fe1",
			1015 => x"01500fe1",
			1016 => x"0c001f04",
			1017 => x"ff101005",
			1018 => x"03003504",
			1019 => x"ff9c1005",
			1020 => x"0200ec04",
			1021 => x"00c41005",
			1022 => x"03006a04",
			1023 => x"ff9e1005",
			1024 => x"00491005",
			1025 => x"03006110",
			1026 => x"0200ba0c",
			1027 => x"03003504",
			1028 => x"ffbf1029",
			1029 => x"0d001904",
			1030 => x"ffec1029",
			1031 => x"005e1029",
			1032 => x"ff691029",
			1033 => x"007c1029",
			1034 => x"03003504",
			1035 => x"ffc4104d",
			1036 => x"0c001f04",
			1037 => x"ffec104d",
			1038 => x"0200f204",
			1039 => x"005a104d",
			1040 => x"01001404",
			1041 => x"000d104d",
			1042 => x"ffed104d",
			1043 => x"0a005c10",
			1044 => x"0b002004",
			1045 => x"fe611079",
			1046 => x"03003504",
			1047 => x"fe6c1079",
			1048 => x"0000f004",
			1049 => x"02c81079",
			1050 => x"fe4a1079",
			1051 => x"01001604",
			1052 => x"01b71079",
			1053 => x"010a1079",
			1054 => x"0b001f08",
			1055 => x"04005004",
			1056 => x"fea410a5",
			1057 => x"ffc410a5",
			1058 => x"03003504",
			1059 => x"ff4c10a5",
			1060 => x"0200e404",
			1061 => x"013210a5",
			1062 => x"03006104",
			1063 => x"ff3d10a5",
			1064 => x"00c210a5",
			1065 => x"0b001f08",
			1066 => x"04005004",
			1067 => x"ff3f10d1",
			1068 => x"ffeb10d1",
			1069 => x"04002004",
			1070 => x"ffc710d1",
			1071 => x"0200f204",
			1072 => x"00b210d1",
			1073 => x"03006e04",
			1074 => x"ffb610d1",
			1075 => x"002e10d1",
			1076 => x"0a00480c",
			1077 => x"0a004504",
			1078 => x"ff0f1105",
			1079 => x"0a004704",
			1080 => x"000b1105",
			1081 => x"ffeb1105",
			1082 => x"0200da08",
			1083 => x"0b001d04",
			1084 => x"ffe91105",
			1085 => x"00c11105",
			1086 => x"03006104",
			1087 => x"ff811105",
			1088 => x"00711105",
			1089 => x"03006114",
			1090 => x"0c002508",
			1091 => x"04004d04",
			1092 => x"fe671131",
			1093 => x"ff671131",
			1094 => x"0000e508",
			1095 => x"04001e04",
			1096 => x"feaf1131",
			1097 => x"01a21131",
			1098 => x"fe4d1131",
			1099 => x"019f1131",
			1100 => x"05008114",
			1101 => x"0f004808",
			1102 => x"0a002d04",
			1103 => x"fff4115d",
			1104 => x"0028115d",
			1105 => x"0c002a04",
			1106 => x"ffb3115d",
			1107 => x"0c002f04",
			1108 => x"0000115d",
			1109 => x"000b115d",
			1110 => x"0039115d",
			1111 => x"03005014",
			1112 => x"0b00240c",
			1113 => x"0b002004",
			1114 => x"fe5a1191",
			1115 => x"07002d04",
			1116 => x"00a11191",
			1117 => x"fe5f1191",
			1118 => x"0a003e04",
			1119 => x"fe601191",
			1120 => x"028e1191",
			1121 => x"0a006504",
			1122 => x"01061191",
			1123 => x"02411191",
			1124 => x"0a005c14",
			1125 => x"0c00250c",
			1126 => x"0b002004",
			1127 => x"fe5b11c5",
			1128 => x"0c002104",
			1129 => x"012911c5",
			1130 => x"fe6011c5",
			1131 => x"0a004204",
			1132 => x"fe6411c5",
			1133 => x"025a11c5",
			1134 => x"01001604",
			1135 => x"01ee11c5",
			1136 => x"017c11c5",
			1137 => x"0b001f08",
			1138 => x"04005004",
			1139 => x"fe7611f9",
			1140 => x"ffe811f9",
			1141 => x"03003504",
			1142 => x"fed411f9",
			1143 => x"0200f208",
			1144 => x"0d002304",
			1145 => x"019211f9",
			1146 => x"00a611f9",
			1147 => x"03006e04",
			1148 => x"fed211f9",
			1149 => x"010111f9",
			1150 => x"0c001f04",
			1151 => x"fe9f1225",
			1152 => x"03003504",
			1153 => x"ff291225",
			1154 => x"01001308",
			1155 => x"0f008a04",
			1156 => x"013c1225",
			1157 => x"00121225",
			1158 => x"0000d704",
			1159 => x"00a21225",
			1160 => x"ff681225",
			1161 => x"0a005c14",
			1162 => x"0b002004",
			1163 => x"fed81251",
			1164 => x"06004a08",
			1165 => x"02002504",
			1166 => x"ffdc1251",
			1167 => x"00a21251",
			1168 => x"0c002a04",
			1169 => x"ff811251",
			1170 => x"001c1251",
			1171 => x"00f31251",
			1172 => x"0a006518",
			1173 => x"0b002008",
			1174 => x"04005004",
			1175 => x"fe651285",
			1176 => x"ff3f1285",
			1177 => x"0000d308",
			1178 => x"04001e04",
			1179 => x"fe7b1285",
			1180 => x"024a1285",
			1181 => x"0d002004",
			1182 => x"ff851285",
			1183 => x"fe431285",
			1184 => x"01a81285",
			1185 => x"0b001f08",
			1186 => x"04005004",
			1187 => x"fe8412b9",
			1188 => x"ffed12b9",
			1189 => x"03003504",
			1190 => x"ff1012b9",
			1191 => x"0f00930c",
			1192 => x"01001104",
			1193 => x"017212b9",
			1194 => x"0000db04",
			1195 => x"00d112b9",
			1196 => x"ffeb12b9",
			1197 => x"ff9212b9",
			1198 => x"03003504",
			1199 => x"ff6512ed",
			1200 => x"0b001f0c",
			1201 => x"0f006c08",
			1202 => x"0200b804",
			1203 => x"ffec12ed",
			1204 => x"002612ed",
			1205 => x"ffbe12ed",
			1206 => x"0200f204",
			1207 => x"008c12ed",
			1208 => x"01001704",
			1209 => x"001e12ed",
			1210 => x"ffd512ed",
			1211 => x"03003504",
			1212 => x"ffbc1321",
			1213 => x"0b001f0c",
			1214 => x"06006908",
			1215 => x"0200b804",
			1216 => x"fff81321",
			1217 => x"00181321",
			1218 => x"ffdc1321",
			1219 => x"0200f204",
			1220 => x"004e1321",
			1221 => x"01001704",
			1222 => x"00101321",
			1223 => x"ffed1321",
			1224 => x"03005514",
			1225 => x"0b002810",
			1226 => x"0a00510c",
			1227 => x"0a004a04",
			1228 => x"fe4c135d",
			1229 => x"08001f04",
			1230 => x"fe4f135d",
			1231 => x"ffd5135d",
			1232 => x"ff75135d",
			1233 => x"001b135d",
			1234 => x"0000cb04",
			1235 => x"074d135d",
			1236 => x"0b002004",
			1237 => x"0554135d",
			1238 => x"0650135d",
			1239 => x"0b001f08",
			1240 => x"04005004",
			1241 => x"fe691399",
			1242 => x"00351399",
			1243 => x"03003504",
			1244 => x"fe831399",
			1245 => x"0200f20c",
			1246 => x"0c002304",
			1247 => x"027a1399",
			1248 => x"0200e404",
			1249 => x"01921399",
			1250 => x"009f1399",
			1251 => x"03006e04",
			1252 => x"fe641399",
			1253 => x"01751399",
			1254 => x"0b001f08",
			1255 => x"04005004",
			1256 => x"fe7413d5",
			1257 => x"ffdf13d5",
			1258 => x"03003504",
			1259 => x"fec813d5",
			1260 => x"0200f20c",
			1261 => x"01001104",
			1262 => x"01b113d5",
			1263 => x"01001804",
			1264 => x"006e13d5",
			1265 => x"012c13d5",
			1266 => x"03006e04",
			1267 => x"fec313d5",
			1268 => x"010a13d5",
			1269 => x"0a004504",
			1270 => x"fe661411",
			1271 => x"0b001f10",
			1272 => x"0f006c04",
			1273 => x"00761411",
			1274 => x"0000f704",
			1275 => x"fe7a1411",
			1276 => x"00010604",
			1277 => x"00441411",
			1278 => x"feba1411",
			1279 => x"0200f208",
			1280 => x"0200e404",
			1281 => x"01a81411",
			1282 => x"011d1411",
			1283 => x"00361411",
			1284 => x"03003504",
			1285 => x"ffae1445",
			1286 => x"0c001f04",
			1287 => x"ffe51445",
			1288 => x"0200da04",
			1289 => x"00631445",
			1290 => x"06007d08",
			1291 => x"08002204",
			1292 => x"00081445",
			1293 => x"ffe21445",
			1294 => x"0f009304",
			1295 => x"00151445",
			1296 => x"fff91445",
			1297 => x"0b001e08",
			1298 => x"05006404",
			1299 => x"fe6e1489",
			1300 => x"ffa81489",
			1301 => x"03003504",
			1302 => x"fe961489",
			1303 => x"0200f210",
			1304 => x"01001108",
			1305 => x"07003504",
			1306 => x"025c1489",
			1307 => x"01731489",
			1308 => x"0c002a04",
			1309 => x"fff21489",
			1310 => x"01681489",
			1311 => x"03006e04",
			1312 => x"fe861489",
			1313 => x"01431489",
			1314 => x"03003504",
			1315 => x"ffc814c7",
			1316 => x"0c001f04",
			1317 => x"ffed14c7",
			1318 => x"0200da04",
			1319 => x"005314c7",
			1320 => x"0b002008",
			1321 => x"08002304",
			1322 => x"ffed14c7",
			1323 => x"000114c7",
			1324 => x"0f007704",
			1325 => x"ffee14c7",
			1326 => x"06008a04",
			1327 => x"001c14c7",
			1328 => x"ffff14c7",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(455, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(899, initial_addr_3'length));
	end generate gen_rom_10;

	gen_rom_11: if SELECT_ROM = 11 generate
		bank <= (
			0 => x"00007c18",
			1 => x"0b00150c",
			2 => x"01000404",
			3 => x"00300075",
			4 => x"0e002404",
			5 => x"00020075",
			6 => x"ffb50075",
			7 => x"06002808",
			8 => x"07002304",
			9 => x"00220075",
			10 => x"ffc40075",
			11 => x"00880075",
			12 => x"0d001314",
			13 => x"06004d04",
			14 => x"ffbe0075",
			15 => x"09001704",
			16 => x"ffd90075",
			17 => x"0f007808",
			18 => x"04003104",
			19 => x"00970075",
			20 => x"fff50075",
			21 => x"ffdf0075",
			22 => x"0c001b08",
			23 => x"01000404",
			24 => x"00020075",
			25 => x"ff7d0075",
			26 => x"02009904",
			27 => x"002f0075",
			28 => x"ffcf0075",
			29 => x"01000a24",
			30 => x"03001c10",
			31 => x"02004608",
			32 => x"0f001b04",
			33 => x"fff400f9",
			34 => x"002900f9",
			35 => x"05001b04",
			36 => x"ffb300f9",
			37 => x"000400f9",
			38 => x"0500410c",
			39 => x"06007208",
			40 => x"08001c04",
			41 => x"005400f9",
			42 => x"fffc00f9",
			43 => x"ffed00f9",
			44 => x"0c001b04",
			45 => x"ffd600f9",
			46 => x"001700f9",
			47 => x"04001c18",
			48 => x"0b001b0c",
			49 => x"06002408",
			50 => x"04000c04",
			51 => x"000a00f9",
			52 => x"ffff00f9",
			53 => x"ffe500f9",
			54 => x"0f002704",
			55 => x"fff600f9",
			56 => x"0c001e04",
			57 => x"000000f9",
			58 => x"002f00f9",
			59 => x"08001904",
			60 => x"000b00f9",
			61 => x"ffaf00f9",
			62 => x"01000414",
			63 => x"05002008",
			64 => x"09001a04",
			65 => x"005c017d",
			66 => x"ffff017d",
			67 => x"03002304",
			68 => x"ffe1017d",
			69 => x"07002804",
			70 => x"0014017d",
			71 => x"fffb017d",
			72 => x"0c00190c",
			73 => x"05000b04",
			74 => x"0011017d",
			75 => x"03003504",
			76 => x"ffac017d",
			77 => x"000d017d",
			78 => x"01000a10",
			79 => x"0a002708",
			80 => x"07002004",
			81 => x"0007017d",
			82 => x"ffeb017d",
			83 => x"04003704",
			84 => x"0059017d",
			85 => x"fff1017d",
			86 => x"04001e0c",
			87 => x"00009408",
			88 => x"00003304",
			89 => x"fff3017d",
			90 => x"003b017d",
			91 => x"fff2017d",
			92 => x"03002704",
			93 => x"0008017d",
			94 => x"ffbc017d",
			95 => x"00007c20",
			96 => x"0c001710",
			97 => x"00004608",
			98 => x"0b001204",
			99 => x"ffdb0209",
			100 => x"006f0209",
			101 => x"0f004604",
			102 => x"ff7d0209",
			103 => x"00020209",
			104 => x"06002808",
			105 => x"07002304",
			106 => x"00280209",
			107 => x"ffb60209",
			108 => x"05001504",
			109 => x"00070209",
			110 => x"00a50209",
			111 => x"08001b20",
			112 => x"06004e04",
			113 => x"ffac0209",
			114 => x"06006610",
			115 => x"05003d08",
			116 => x"07002204",
			117 => x"00000209",
			118 => x"00910209",
			119 => x"07002904",
			120 => x"ffc40209",
			121 => x"00120209",
			122 => x"0c001604",
			123 => x"ffb10209",
			124 => x"09001b04",
			125 => x"002b0209",
			126 => x"ffee0209",
			127 => x"0b002f04",
			128 => x"ff570209",
			129 => x"00250209",
			130 => x"05002b2c",
			131 => x"00007510",
			132 => x"0b001204",
			133 => x"ffe402a5",
			134 => x"02002004",
			135 => x"ffee02a5",
			136 => x"09002a04",
			137 => x"006a02a5",
			138 => x"000102a5",
			139 => x"06004e04",
			140 => x"ffa902a5",
			141 => x"0600670c",
			142 => x"08001b04",
			143 => x"005302a5",
			144 => x"0b001a04",
			145 => x"ffe402a5",
			146 => x"000f02a5",
			147 => x"0c001604",
			148 => x"ffd302a5",
			149 => x"0d001304",
			150 => x"001802a5",
			151 => x"fff802a5",
			152 => x"0c001b14",
			153 => x"08001608",
			154 => x"03002d04",
			155 => x"001102a5",
			156 => x"fffb02a5",
			157 => x"0f004304",
			158 => x"000302a5",
			159 => x"0b001904",
			160 => x"ff9f02a5",
			161 => x"ffff02a5",
			162 => x"08001d08",
			163 => x"04003704",
			164 => x"004902a5",
			165 => x"fff502a5",
			166 => x"04001f04",
			167 => x"001002a5",
			168 => x"ffc902a5",
			169 => x"04001424",
			170 => x"03001a1c",
			171 => x"04000c0c",
			172 => x"00002104",
			173 => x"fff40349",
			174 => x"04000504",
			175 => x"00000349",
			176 => x"00390349",
			177 => x"05001b0c",
			178 => x"0c001f08",
			179 => x"0e001d04",
			180 => x"00010349",
			181 => x"ffad0349",
			182 => x"00030349",
			183 => x"00130349",
			184 => x"06007b04",
			185 => x"00570349",
			186 => x"fffb0349",
			187 => x"0c001b18",
			188 => x"0e003a08",
			189 => x"01000b04",
			190 => x"002f0349",
			191 => x"ffec0349",
			192 => x"01000304",
			193 => x"000e0349",
			194 => x"0b001904",
			195 => x"ff870349",
			196 => x"0d001504",
			197 => x"00090349",
			198 => x"ffff0349",
			199 => x"0d001608",
			200 => x"04003704",
			201 => x"004e0349",
			202 => x"fff50349",
			203 => x"04001c0c",
			204 => x"0f002804",
			205 => x"fffa0349",
			206 => x"0d001a04",
			207 => x"fffc0349",
			208 => x"00260349",
			209 => x"ffb60349",
			210 => x"0e003a20",
			211 => x"01000b10",
			212 => x"0b001204",
			213 => x"ffcd03e5",
			214 => x"02006b08",
			215 => x"00002104",
			216 => x"ffe603e5",
			217 => x"00a403e5",
			218 => x"fff103e5",
			219 => x"0400140c",
			220 => x"02002904",
			221 => x"fff403e5",
			222 => x"02004c04",
			223 => x"002a03e5",
			224 => x"fffb03e5",
			225 => x"ffb703e5",
			226 => x"0c001b24",
			227 => x"0400140c",
			228 => x"09001704",
			229 => x"ffc103e5",
			230 => x"06007004",
			231 => x"007e03e5",
			232 => x"ffef03e5",
			233 => x"01000304",
			234 => x"002a03e5",
			235 => x"0b00190c",
			236 => x"0d000f04",
			237 => x"fffe03e5",
			238 => x"08001604",
			239 => x"ffe603e5",
			240 => x"ff3903e5",
			241 => x"0d001504",
			242 => x"001703e5",
			243 => x"ffdd03e5",
			244 => x"02009904",
			245 => x"008303e5",
			246 => x"01000704",
			247 => x"001903e5",
			248 => x"ffb103e5",
			249 => x"04001424",
			250 => x"0c001104",
			251 => x"ffe00489",
			252 => x"0a00160c",
			253 => x"00005208",
			254 => x"02002004",
			255 => x"fff00489",
			256 => x"00370489",
			257 => x"ffcd0489",
			258 => x"06006b0c",
			259 => x"00003704",
			260 => x"fffd0489",
			261 => x"00009f04",
			262 => x"00630489",
			263 => x"ffff0489",
			264 => x"05001e04",
			265 => x"00010489",
			266 => x"fffc0489",
			267 => x"0c001b18",
			268 => x"0e003a08",
			269 => x"0c001604",
			270 => x"ffe60489",
			271 => x"003c0489",
			272 => x"01000304",
			273 => x"000e0489",
			274 => x"0b001904",
			275 => x"ff8d0489",
			276 => x"0d001504",
			277 => x"00090489",
			278 => x"ffff0489",
			279 => x"0d001608",
			280 => x"04003704",
			281 => x"004d0489",
			282 => x"fff50489",
			283 => x"04001c0c",
			284 => x"0f002804",
			285 => x"fffa0489",
			286 => x"0d001a04",
			287 => x"fffc0489",
			288 => x"00250489",
			289 => x"ffb80489",
			290 => x"05002b34",
			291 => x"03001c1c",
			292 => x"0500150c",
			293 => x"0f001b04",
			294 => x"ffe1053d",
			295 => x"04000504",
			296 => x"fffe053d",
			297 => x"0069053d",
			298 => x"0a001e0c",
			299 => x"08002404",
			300 => x"ff67053d",
			301 => x"08002604",
			302 => x"0004053d",
			303 => x"fffa053d",
			304 => x"0000053d",
			305 => x"0f007a14",
			306 => x"01000a04",
			307 => x"00be053d",
			308 => x"0d001908",
			309 => x"02005c04",
			310 => x"000d053d",
			311 => x"ffbd053d",
			312 => x"00003d04",
			313 => x"fff8053d",
			314 => x"003d053d",
			315 => x"ffb5053d",
			316 => x"0c001b18",
			317 => x"0f004304",
			318 => x"0010053d",
			319 => x"08001608",
			320 => x"01000504",
			321 => x"fffb053d",
			322 => x"0024053d",
			323 => x"0d001104",
			324 => x"0004053d",
			325 => x"0b001904",
			326 => x"ff18053d",
			327 => x"fff2053d",
			328 => x"08001d08",
			329 => x"05004a04",
			330 => x"00a7053d",
			331 => x"fff0053d",
			332 => x"04001f04",
			333 => x"0019053d",
			334 => x"ff8d053d",
			335 => x"01000a30",
			336 => x"0e005020",
			337 => x"0b001204",
			338 => x"ff9d05e9",
			339 => x"08001d14",
			340 => x"0400220c",
			341 => x"05002608",
			342 => x"05002104",
			343 => x"001e05e9",
			344 => x"00b405e9",
			345 => x"ffb805e9",
			346 => x"0f005904",
			347 => x"00d305e9",
			348 => x"ffef05e9",
			349 => x"00004904",
			350 => x"000905e9",
			351 => x"ffcf05e9",
			352 => x"02009704",
			353 => x"ff4305e9",
			354 => x"05003c08",
			355 => x"06007204",
			356 => x"00d905e9",
			357 => x"ffa105e9",
			358 => x"ff6b05e9",
			359 => x"0e003d18",
			360 => x"0b001604",
			361 => x"ffb705e9",
			362 => x"0b00200c",
			363 => x"00007c08",
			364 => x"00003304",
			365 => x"fff405e9",
			366 => x"00a105e9",
			367 => x"ffed05e9",
			368 => x"08002304",
			369 => x"000b05e9",
			370 => x"ffb005e9",
			371 => x"09003008",
			372 => x"08001804",
			373 => x"002605e9",
			374 => x"ff0705e9",
			375 => x"0a003b04",
			376 => x"005705e9",
			377 => x"ffe805e9",
			378 => x"02009a44",
			379 => x"03001c24",
			380 => x"05001514",
			381 => x"01000404",
			382 => x"004a067d",
			383 => x"0a001108",
			384 => x"05000b04",
			385 => x"0005067d",
			386 => x"ffd1067d",
			387 => x"00002f04",
			388 => x"fffb067d",
			389 => x"0016067d",
			390 => x"0b001808",
			391 => x"05001b04",
			392 => x"ff99067d",
			393 => x"fffb067d",
			394 => x"09002704",
			395 => x"0013067d",
			396 => x"fff5067d",
			397 => x"04001c08",
			398 => x"00003504",
			399 => x"fffc067d",
			400 => x"0073067d",
			401 => x"0b00170c",
			402 => x"0e003a04",
			403 => x"0005067d",
			404 => x"0e004e04",
			405 => x"ffb0067d",
			406 => x"0006067d",
			407 => x"07002908",
			408 => x"0e004504",
			409 => x"0069067d",
			410 => x"0007067d",
			411 => x"ffd7067d",
			412 => x"08001604",
			413 => x"fffa067d",
			414 => x"ff8f067d",
			415 => x"01000a38",
			416 => x"0c001514",
			417 => x"0d000f0c",
			418 => x"0b001004",
			419 => x"ffe20721",
			420 => x"01000504",
			421 => x"00490721",
			422 => x"00030721",
			423 => x"08001604",
			424 => x"00080721",
			425 => x"ffa40721",
			426 => x"0400331c",
			427 => x"0f007918",
			428 => x"0a00180c",
			429 => x"00006b08",
			430 => x"00002504",
			431 => x"fff70721",
			432 => x"00170721",
			433 => x"ffe50721",
			434 => x"08001d08",
			435 => x"09001e04",
			436 => x"00820721",
			437 => x"001b0721",
			438 => x"fff80721",
			439 => x"ffeb0721",
			440 => x"01000904",
			441 => x"ffc90721",
			442 => x"00160721",
			443 => x"09003014",
			444 => x"08001804",
			445 => x"000f0721",
			446 => x"05000d04",
			447 => x"00050721",
			448 => x"05003f04",
			449 => x"ff9b0721",
			450 => x"05004004",
			451 => x"00180721",
			452 => x"ffe20721",
			453 => x"04001b04",
			454 => x"00290721",
			455 => x"fff30721",
			456 => x"0e005240",
			457 => x"0c001820",
			458 => x"05002b18",
			459 => x"0c001304",
			460 => x"ff3107e5",
			461 => x"08001c10",
			462 => x"0c001608",
			463 => x"0a001404",
			464 => x"001f07e5",
			465 => x"010d07e5",
			466 => x"00006e04",
			467 => x"00a407e5",
			468 => x"ff5107e5",
			469 => x"ff8107e5",
			470 => x"0f005a04",
			471 => x"ff0007e5",
			472 => x"fffb07e5",
			473 => x"08001d10",
			474 => x"0e004308",
			475 => x"00002f04",
			476 => x"ffb707e5",
			477 => x"012e07e5",
			478 => x"0c001904",
			479 => x"ffb807e5",
			480 => x"009007e5",
			481 => x"04001c0c",
			482 => x"00007c08",
			483 => x"00003504",
			484 => x"ffba07e5",
			485 => x"00cf07e5",
			486 => x"ffa207e5",
			487 => x"ff4c07e5",
			488 => x"0a002810",
			489 => x"0c001608",
			490 => x"0d001004",
			491 => x"006c07e5",
			492 => x"ff0607e5",
			493 => x"0f007d04",
			494 => x"00d007e5",
			495 => x"ffce07e5",
			496 => x"08001608",
			497 => x"05003204",
			498 => x"ffe207e5",
			499 => x"004907e5",
			500 => x"0c001b04",
			501 => x"feba07e5",
			502 => x"0000ad04",
			503 => x"005507e5",
			504 => x"ff4a07e5",
			505 => x"0e006134",
			506 => x"05002b18",
			507 => x"0c001104",
			508 => x"feaa0851",
			509 => x"02002004",
			510 => x"fec00851",
			511 => x"0e002204",
			512 => x"019d0851",
			513 => x"0c001304",
			514 => x"feaa0851",
			515 => x"0a001604",
			516 => x"ff6b0851",
			517 => x"00c80851",
			518 => x"08001d14",
			519 => x"0c001b10",
			520 => x"08001604",
			521 => x"01230851",
			522 => x"00007c04",
			523 => x"005a0851",
			524 => x"01000404",
			525 => x"00390851",
			526 => x"fe6a0851",
			527 => x"016d0851",
			528 => x"07003304",
			529 => x"fe450851",
			530 => x"00360851",
			531 => x"fe740851",
			532 => x"0700252c",
			533 => x"02006b18",
			534 => x"0b001204",
			535 => x"fe6308ed",
			536 => x"01000404",
			537 => x"032808ed",
			538 => x"0c001504",
			539 => x"ff8108ed",
			540 => x"0b001504",
			541 => x"011a08ed",
			542 => x"07002304",
			543 => x"025108ed",
			544 => x"016908ed",
			545 => x"04001304",
			546 => x"fe5508ed",
			547 => x"05002608",
			548 => x"0f005904",
			549 => x"008708ed",
			550 => x"022b08ed",
			551 => x"00008804",
			552 => x"012d08ed",
			553 => x"fe5508ed",
			554 => x"0200a21c",
			555 => x"00002f04",
			556 => x"fe5b08ed",
			557 => x"03003914",
			558 => x"0c001b0c",
			559 => x"0d001304",
			560 => x"011808ed",
			561 => x"06005504",
			562 => x"ffce08ed",
			563 => x"fe4c08ed",
			564 => x"0a002c04",
			565 => x"00eb08ed",
			566 => x"033d08ed",
			567 => x"fe1c08ed",
			568 => x"0a002004",
			569 => x"fff908ed",
			570 => x"fe5808ed",
			571 => x"0e00391c",
			572 => x"0b00150c",
			573 => x"06002204",
			574 => x"006b09a9",
			575 => x"00004604",
			576 => x"fff809a9",
			577 => x"ff4709a9",
			578 => x"07002308",
			579 => x"00007504",
			580 => x"00f509a9",
			581 => x"ffdf09a9",
			582 => x"06002904",
			583 => x"ff8409a9",
			584 => x"003709a9",
			585 => x"0c001b34",
			586 => x"08001818",
			587 => x"03001f08",
			588 => x"06008004",
			589 => x"006509a9",
			590 => x"fff909a9",
			591 => x"01000a0c",
			592 => x"0c001708",
			593 => x"0c001604",
			594 => x"ffe709a9",
			595 => x"001209a9",
			596 => x"ff8b09a9",
			597 => x"002a09a9",
			598 => x"0b001910",
			599 => x"00009b04",
			600 => x"fee209a9",
			601 => x"08001b08",
			602 => x"0000ad04",
			603 => x"006509a9",
			604 => x"ffcd09a9",
			605 => x"ff5e09a9",
			606 => x"0d001704",
			607 => x"ffd309a9",
			608 => x"0d001904",
			609 => x"002e09a9",
			610 => x"ffec09a9",
			611 => x"01000a08",
			612 => x"05004704",
			613 => x"00c509a9",
			614 => x"ffdc09a9",
			615 => x"02009204",
			616 => x"003709a9",
			617 => x"ff7009a9",
			618 => x"07002740",
			619 => x"00007c28",
			620 => x"0b001510",
			621 => x"00004608",
			622 => x"0b001204",
			623 => x"fe830a65",
			624 => x"026f0a65",
			625 => x"01000704",
			626 => x"00850a65",
			627 => x"fe350a65",
			628 => x"00002804",
			629 => x"fe060a65",
			630 => x"08001d08",
			631 => x"00005e04",
			632 => x"01f00a65",
			633 => x"02ec0a65",
			634 => x"02004e08",
			635 => x"06002804",
			636 => x"016f0a65",
			637 => x"01f70a65",
			638 => x"01200a65",
			639 => x"0100060c",
			640 => x"03002d08",
			641 => x"0200af04",
			642 => x"01a80a65",
			643 => x"fe630a65",
			644 => x"fe5a0a65",
			645 => x"0a003808",
			646 => x"0f006104",
			647 => x"fe4b0a65",
			648 => x"ff360a65",
			649 => x"008c0a65",
			650 => x"0000aa1c",
			651 => x"0600370c",
			652 => x"07002808",
			653 => x"00001204",
			654 => x"fe800a65",
			655 => x"00350a65",
			656 => x"fe580a65",
			657 => x"03003a0c",
			658 => x"07002a08",
			659 => x"01000b04",
			660 => x"00df0a65",
			661 => x"fe570a65",
			662 => x"02650a65",
			663 => x"fe3a0a65",
			664 => x"fe5d0a65",
			665 => x"02009a34",
			666 => x"0c001104",
			667 => x"ffd20af1",
			668 => x"08001d20",
			669 => x"05004118",
			670 => x"05002310",
			671 => x"0c001608",
			672 => x"05001a04",
			673 => x"004e0af1",
			674 => x"fffe0af1",
			675 => x"00006b04",
			676 => x"000d0af1",
			677 => x"ffb70af1",
			678 => x"0c001604",
			679 => x"fff60af1",
			680 => x"00870af1",
			681 => x"04003404",
			682 => x"001b0af1",
			683 => x"ffd60af1",
			684 => x"04001c0c",
			685 => x"02003804",
			686 => x"fff20af1",
			687 => x"09001e04",
			688 => x"fff90af1",
			689 => x"00440af1",
			690 => x"ffb50af1",
			691 => x"01000610",
			692 => x"0a002808",
			693 => x"0200ae04",
			694 => x"00340af1",
			695 => x"fffb0af1",
			696 => x"09002104",
			697 => x"ffd80af1",
			698 => x"00110af1",
			699 => x"ffad0af1",
			700 => x"07002538",
			701 => x"0f003318",
			702 => x"0b001204",
			703 => x"fe6f0b95",
			704 => x"07002310",
			705 => x"00003304",
			706 => x"02c00b95",
			707 => x"0f002e08",
			708 => x"01000e04",
			709 => x"02030b95",
			710 => x"01b50b95",
			711 => x"01430b95",
			712 => x"00c40b95",
			713 => x"0c001714",
			714 => x"0100060c",
			715 => x"0000af08",
			716 => x"06004e04",
			717 => x"00350b95",
			718 => x"02180b95",
			719 => x"fe730b95",
			720 => x"08001804",
			721 => x"ffe30b95",
			722 => x"fe410b95",
			723 => x"02007404",
			724 => x"02d80b95",
			725 => x"0e004404",
			726 => x"fe550b95",
			727 => x"010d0b95",
			728 => x"0200ae18",
			729 => x"00002f04",
			730 => x"fe600b95",
			731 => x"04003310",
			732 => x"0c001604",
			733 => x"fe530b95",
			734 => x"01000a04",
			735 => x"01fa0b95",
			736 => x"05003304",
			737 => x"00ff0b95",
			738 => x"fe100b95",
			739 => x"fe560b95",
			740 => x"fe5c0b95",
			741 => x"0200ae38",
			742 => x"05002b20",
			743 => x"0c001104",
			744 => x"fea20c09",
			745 => x"02002004",
			746 => x"feb40c09",
			747 => x"0200460c",
			748 => x"09002a08",
			749 => x"01000e04",
			750 => x"01a00c09",
			751 => x"00960c09",
			752 => x"ff3d0c09",
			753 => x"07001d04",
			754 => x"fec30c09",
			755 => x"00007804",
			756 => x"014f0c09",
			757 => x"00410c09",
			758 => x"08001d10",
			759 => x"0b00190c",
			760 => x"05004108",
			761 => x"0c001604",
			762 => x"feb80c09",
			763 => x"00950c09",
			764 => x"fe880c09",
			765 => x"01280c09",
			766 => x"07002c04",
			767 => x"fe300c09",
			768 => x"ffdc0c09",
			769 => x"fe720c09",
			770 => x"0e006130",
			771 => x"0500412c",
			772 => x"0800180c",
			773 => x"0b001204",
			774 => x"ffab0c6d",
			775 => x"0a002304",
			776 => x"015e0c6d",
			777 => x"00750c6d",
			778 => x"0c001608",
			779 => x"06002704",
			780 => x"00010c6d",
			781 => x"fec20c6d",
			782 => x"0700220c",
			783 => x"02006b08",
			784 => x"0a000f04",
			785 => x"00110c6d",
			786 => x"014b0c6d",
			787 => x"ff9b0c6d",
			788 => x"06002804",
			789 => x"fee80c6d",
			790 => x"0a002f04",
			791 => x"ffd80c6d",
			792 => x"00ed0c6d",
			793 => x"fec20c6d",
			794 => x"fea00c6d",
			795 => x"04001420",
			796 => x"0a00160c",
			797 => x"05000c08",
			798 => x"00004104",
			799 => x"00650d29",
			800 => x"fffa0d29",
			801 => x"ff760d29",
			802 => x"06006b0c",
			803 => x"00009f08",
			804 => x"00003504",
			805 => x"fff50d29",
			806 => x"00c80d29",
			807 => x"fff70d29",
			808 => x"0b001404",
			809 => x"ffa80d29",
			810 => x"00480d29",
			811 => x"0c00180c",
			812 => x"06003104",
			813 => x"001f0d29",
			814 => x"0b001704",
			815 => x"ff340d29",
			816 => x"00070d29",
			817 => x"0d001308",
			818 => x"04003304",
			819 => x"00bf0d29",
			820 => x"fff50d29",
			821 => x"02008b14",
			822 => x"08001d04",
			823 => x"00ac0d29",
			824 => x"07003308",
			825 => x"0a002c04",
			826 => x"00050d29",
			827 => x"ffa80d29",
			828 => x"01001404",
			829 => x"fff80d29",
			830 => x"002e0d29",
			831 => x"0900240c",
			832 => x"07002b04",
			833 => x"ff120d29",
			834 => x"07002c04",
			835 => x"002b0d29",
			836 => x"ffd10d29",
			837 => x"01000904",
			838 => x"002d0d29",
			839 => x"08003504",
			840 => x"ffcc0d29",
			841 => x"00180d29",
			842 => x"07002948",
			843 => x"00007c28",
			844 => x"00002104",
			845 => x"fe4a0de5",
			846 => x"0c001714",
			847 => x"06002408",
			848 => x"01000704",
			849 => x"024f0de5",
			850 => x"015d0de5",
			851 => x"01000a08",
			852 => x"03001804",
			853 => x"feb50de5",
			854 => x"00bc0de5",
			855 => x"fe480de5",
			856 => x"0800230c",
			857 => x"05002308",
			858 => x"0a001104",
			859 => x"01390de5",
			860 => x"01be0de5",
			861 => x"022a0de5",
			862 => x"00cc0de5",
			863 => x"0d001310",
			864 => x"0200ae0c",
			865 => x"06004d04",
			866 => x"fe370de5",
			867 => x"04003104",
			868 => x"01d30de5",
			869 => x"fe850de5",
			870 => x"fe680de5",
			871 => x"0c001b08",
			872 => x"09001b04",
			873 => x"ff9e0de5",
			874 => x"fe4e0de5",
			875 => x"04001d04",
			876 => x"fe6a0de5",
			877 => x"00ef0de5",
			878 => x"0c002c14",
			879 => x"0e005a10",
			880 => x"08001c08",
			881 => x"0c001b04",
			882 => x"fe820de5",
			883 => x"01aa0de5",
			884 => x"0d002204",
			885 => x"fe5a0de5",
			886 => x"ff3c0de5",
			887 => x"fe610de5",
			888 => x"00e60de5",
			889 => x"0200ae34",
			890 => x"05004130",
			891 => x"0800180c",
			892 => x"09001804",
			893 => x"00770e51",
			894 => x"06004504",
			895 => x"00560e51",
			896 => x"014b0e51",
			897 => x"0c00160c",
			898 => x"06002704",
			899 => x"00020e51",
			900 => x"00009604",
			901 => x"fea30e51",
			902 => x"ffde0e51",
			903 => x"0700220c",
			904 => x"02006b08",
			905 => x"0a000f04",
			906 => x"00130e51",
			907 => x"01530e51",
			908 => x"ff940e51",
			909 => x"06002804",
			910 => x"feda0e51",
			911 => x"0a002f04",
			912 => x"ffcf0e51",
			913 => x"00fd0e51",
			914 => x"fec00e51",
			915 => x"fe9a0e51",
			916 => x"0e005d3c",
			917 => x"0c001104",
			918 => x"ffbc0ed5",
			919 => x"05002b1c",
			920 => x"07002510",
			921 => x"0c001304",
			922 => x"00010ed5",
			923 => x"04000504",
			924 => x"fffe0ed5",
			925 => x"09001e04",
			926 => x"00970ed5",
			927 => x"000d0ed5",
			928 => x"06005308",
			929 => x"0a000b04",
			930 => x"00030ed5",
			931 => x"ffb00ed5",
			932 => x"00510ed5",
			933 => x"0c001b10",
			934 => x"0f004304",
			935 => x"00190ed5",
			936 => x"08001604",
			937 => x"00200ed5",
			938 => x"0b001904",
			939 => x"ff6c0ed5",
			940 => x"00090ed5",
			941 => x"0d001704",
			942 => x"00730ed5",
			943 => x"01001104",
			944 => x"ffce0ed5",
			945 => x"ffff0ed5",
			946 => x"07002704",
			947 => x"fffb0ed5",
			948 => x"ff9f0ed5",
			949 => x"0200ae44",
			950 => x"04000e10",
			951 => x"00002104",
			952 => x"ff4c0f61",
			953 => x"02005804",
			954 => x"01480f61",
			955 => x"06004504",
			956 => x"ff300f61",
			957 => x"00d10f61",
			958 => x"01000b18",
			959 => x"0c001304",
			960 => x"feb00f61",
			961 => x"0500410c",
			962 => x"0a002d08",
			963 => x"09001e04",
			964 => x"00650f61",
			965 => x"ff390f61",
			966 => x"01320f61",
			967 => x"09002104",
			968 => x"fe990f61",
			969 => x"00790f61",
			970 => x"04001c14",
			971 => x"0a00240c",
			972 => x"05001608",
			973 => x"07002804",
			974 => x"003d0f61",
			975 => x"ffe60f61",
			976 => x"fefd0f61",
			977 => x"09002404",
			978 => x"00470f61",
			979 => x"01120f61",
			980 => x"0d001504",
			981 => x"ff4e0f61",
			982 => x"fe7f0f61",
			983 => x"fe7d0f61",
			984 => x"0e006134",
			985 => x"0500412c",
			986 => x"0b001204",
			987 => x"fede0fcd",
			988 => x"0800180c",
			989 => x"06005008",
			990 => x"00005204",
			991 => x"01300fcd",
			992 => x"ffe80fcd",
			993 => x"014b0fcd",
			994 => x"0c00160c",
			995 => x"06003004",
			996 => x"00140fcd",
			997 => x"07002204",
			998 => x"feb10fcd",
			999 => x"ffd50fcd",
			1000 => x"07002208",
			1001 => x"02006b04",
			1002 => x"013b0fcd",
			1003 => x"ff8c0fcd",
			1004 => x"05003a04",
			1005 => x"ffab0fcd",
			1006 => x"00e80fcd",
			1007 => x"09002404",
			1008 => x"feaf0fcd",
			1009 => x"009f0fcd",
			1010 => x"fe940fcd",
			1011 => x"0200a548",
			1012 => x"0700252c",
			1013 => x"0c001820",
			1014 => x"01000a18",
			1015 => x"02006b0c",
			1016 => x"0b001204",
			1017 => x"fe9b1061",
			1018 => x"00004804",
			1019 => x"01e11061",
			1020 => x"01371061",
			1021 => x"06004e04",
			1022 => x"fe341061",
			1023 => x"03002e04",
			1024 => x"01141061",
			1025 => x"fef41061",
			1026 => x"04001204",
			1027 => x"ffb61061",
			1028 => x"fe5f1061",
			1029 => x"02007408",
			1030 => x"0a001204",
			1031 => x"00c31061",
			1032 => x"01bd1061",
			1033 => x"fff71061",
			1034 => x"00002f04",
			1035 => x"fe751061",
			1036 => x"0b00190c",
			1037 => x"08001904",
			1038 => x"005b1061",
			1039 => x"05002804",
			1040 => x"ff901061",
			1041 => x"fe5a1061",
			1042 => x"03003a08",
			1043 => x"02009204",
			1044 => x"01af1061",
			1045 => x"00421061",
			1046 => x"fe7c1061",
			1047 => x"fe661061",
			1048 => x"0e006140",
			1049 => x"08001d20",
			1050 => x"0500461c",
			1051 => x"0a003614",
			1052 => x"0c001104",
			1053 => x"ff2f10e5",
			1054 => x"05002b08",
			1055 => x"0f005604",
			1056 => x"004910e5",
			1057 => x"012610e5",
			1058 => x"0c001604",
			1059 => x"ff1310e5",
			1060 => x"004310e5",
			1061 => x"0b001704",
			1062 => x"ffb910e5",
			1063 => x"015d10e5",
			1064 => x"ff2a10e5",
			1065 => x"04001c1c",
			1066 => x"0b001b10",
			1067 => x"0600310c",
			1068 => x"02003608",
			1069 => x"0a000f04",
			1070 => x"000510e5",
			1071 => x"ffdb10e5",
			1072 => x"003810e5",
			1073 => x"ff7410e5",
			1074 => x"00003704",
			1075 => x"ffaf10e5",
			1076 => x"00009f04",
			1077 => x"010510e5",
			1078 => x"ffd510e5",
			1079 => x"fed410e5",
			1080 => x"fec210e5",
			1081 => x"01000414",
			1082 => x"05002008",
			1083 => x"09001a04",
			1084 => x"005f11a9",
			1085 => x"ffff11a9",
			1086 => x"03002304",
			1087 => x"ffdf11a9",
			1088 => x"07002804",
			1089 => x"001411a9",
			1090 => x"fffb11a9",
			1091 => x"0c001710",
			1092 => x"05000d04",
			1093 => x"000b11a9",
			1094 => x"0b001708",
			1095 => x"09001e04",
			1096 => x"ffa111a9",
			1097 => x"000211a9",
			1098 => x"000511a9",
			1099 => x"05004134",
			1100 => x"0a00271c",
			1101 => x"07002510",
			1102 => x"00006e08",
			1103 => x"0e002004",
			1104 => x"fffd11a9",
			1105 => x"002011a9",
			1106 => x"0f004104",
			1107 => x"fff211a9",
			1108 => x"000511a9",
			1109 => x"01001408",
			1110 => x"05000f04",
			1111 => x"000011a9",
			1112 => x"ffcc11a9",
			1113 => x"000011a9",
			1114 => x"08001c08",
			1115 => x"0000aa04",
			1116 => x"007111a9",
			1117 => x"fff811a9",
			1118 => x"0c002008",
			1119 => x"03002704",
			1120 => x"000611a9",
			1121 => x"ffd311a9",
			1122 => x"0a003b04",
			1123 => x"002811a9",
			1124 => x"fff311a9",
			1125 => x"0b001a04",
			1126 => x"ffba11a9",
			1127 => x"03003904",
			1128 => x"002711a9",
			1129 => x"fff911a9",
			1130 => x"0200ae38",
			1131 => x"02002004",
			1132 => x"fe78121d",
			1133 => x"04001c18",
			1134 => x"0c001104",
			1135 => x"fe57121d",
			1136 => x"06007010",
			1137 => x"02005008",
			1138 => x"09002a04",
			1139 => x"0197121d",
			1140 => x"fee7121d",
			1141 => x"0a001604",
			1142 => x"fe78121d",
			1143 => x"010d121d",
			1144 => x"fe9a121d",
			1145 => x"08001d14",
			1146 => x"0c001a0c",
			1147 => x"05004108",
			1148 => x"0c001604",
			1149 => x"ff33121d",
			1150 => x"00ec121d",
			1151 => x"fe6d121d",
			1152 => x"05004704",
			1153 => x"0198121d",
			1154 => x"feea121d",
			1155 => x"09002404",
			1156 => x"fe6d121d",
			1157 => x"fda7121d",
			1158 => x"fe69121d",
			1159 => x"0e006148",
			1160 => x"0c001b28",
			1161 => x"05004024",
			1162 => x"08001b14",
			1163 => x"0c001104",
			1164 => x"ff7412b1",
			1165 => x"0f005408",
			1166 => x"00007504",
			1167 => x"007f12b1",
			1168 => x"ff2d12b1",
			1169 => x"0000b804",
			1170 => x"00df12b1",
			1171 => x"fff312b1",
			1172 => x"0e00410c",
			1173 => x"0c001604",
			1174 => x"ff5e12b1",
			1175 => x"00002804",
			1176 => x"ffe212b1",
			1177 => x"00c112b1",
			1178 => x"ff0512b1",
			1179 => x"ff0c12b1",
			1180 => x"01000a10",
			1181 => x"0a00270c",
			1182 => x"0c001c08",
			1183 => x"03001004",
			1184 => x"fffc12b1",
			1185 => x"000812b1",
			1186 => x"ffde12b1",
			1187 => x"00fe12b1",
			1188 => x"0000940c",
			1189 => x"06002808",
			1190 => x"07002304",
			1191 => x"002512b1",
			1192 => x"ff9012b1",
			1193 => x"00a912b1",
			1194 => x"ff7112b1",
			1195 => x"ff1912b1",
			1196 => x"0f007844",
			1197 => x"0500413c",
			1198 => x"03001c20",
			1199 => x"05001514",
			1200 => x"01000404",
			1201 => x"0056133d",
			1202 => x"0a001108",
			1203 => x"05000b04",
			1204 => x"000b133d",
			1205 => x"ffce133d",
			1206 => x"02006e04",
			1207 => x"0022133d",
			1208 => x"fff3133d",
			1209 => x"05001b04",
			1210 => x"ff90133d",
			1211 => x"05001c04",
			1212 => x"001f133d",
			1213 => x"ffd8133d",
			1214 => x"04001c0c",
			1215 => x"00003904",
			1216 => x"fffb133d",
			1217 => x"05002504",
			1218 => x"0095133d",
			1219 => x"000a133d",
			1220 => x"08001c0c",
			1221 => x"09001d08",
			1222 => x"00009404",
			1223 => x"ffb6133d",
			1224 => x"000b133d",
			1225 => x"007d133d",
			1226 => x"ffa9133d",
			1227 => x"0b001a04",
			1228 => x"ff8a133d",
			1229 => x"003e133d",
			1230 => x"ffa3133d",
			1231 => x"0000aa3c",
			1232 => x"02002004",
			1233 => x"fe5313c1",
			1234 => x"00005c18",
			1235 => x"0b001204",
			1236 => x"fe7613c1",
			1237 => x"0100100c",
			1238 => x"01000504",
			1239 => x"027413c1",
			1240 => x"01000e04",
			1241 => x"01c813c1",
			1242 => x"015213c1",
			1243 => x"04001804",
			1244 => x"017b13c1",
			1245 => x"fe2113c1",
			1246 => x"08001604",
			1247 => x"01ac13c1",
			1248 => x"0c001a10",
			1249 => x"01000608",
			1250 => x"07002404",
			1251 => x"00ad13c1",
			1252 => x"ff8013c1",
			1253 => x"0e003804",
			1254 => x"007313c1",
			1255 => x"fe7313c1",
			1256 => x"03003a08",
			1257 => x"0a002304",
			1258 => x"ff8a13c1",
			1259 => x"020613c1",
			1260 => x"fe2a13c1",
			1261 => x"05001c04",
			1262 => x"007113c1",
			1263 => x"fe5f13c1",
			1264 => x"0e00614c",
			1265 => x"08001b20",
			1266 => x"0500411c",
			1267 => x"0c001104",
			1268 => x"fee7145d",
			1269 => x"0f004b10",
			1270 => x"02004608",
			1271 => x"00002104",
			1272 => x"ffcd145d",
			1273 => x"015d145d",
			1274 => x"03001f04",
			1275 => x"fed0145d",
			1276 => x"0088145d",
			1277 => x"0b001304",
			1278 => x"0085145d",
			1279 => x"0171145d",
			1280 => x"fec3145d",
			1281 => x"0b001910",
			1282 => x"0e00380c",
			1283 => x"0b001504",
			1284 => x"fef0145d",
			1285 => x"00002804",
			1286 => x"ffb0145d",
			1287 => x"0136145d",
			1288 => x"fe8c145d",
			1289 => x"01000808",
			1290 => x"03001a04",
			1291 => x"fff3145d",
			1292 => x"013e145d",
			1293 => x"04001e0c",
			1294 => x"00003304",
			1295 => x"ff2f145d",
			1296 => x"00009404",
			1297 => x"0146145d",
			1298 => x"ff35145d",
			1299 => x"0a003204",
			1300 => x"ffc6145d",
			1301 => x"fea4145d",
			1302 => x"fe87145d",
			1303 => x"0f006e48",
			1304 => x"0c001308",
			1305 => x"0f002504",
			1306 => x"000c14f1",
			1307 => x"ffbe14f1",
			1308 => x"0500261c",
			1309 => x"0a00160c",
			1310 => x"00005208",
			1311 => x"00002504",
			1312 => x"ffeb14f1",
			1313 => x"004014f1",
			1314 => x"ffc114f1",
			1315 => x"04001c0c",
			1316 => x"00003504",
			1317 => x"fff314f1",
			1318 => x"0000a104",
			1319 => x"008114f1",
			1320 => x"fffd14f1",
			1321 => x"fff914f1",
			1322 => x"0c001910",
			1323 => x"0600610c",
			1324 => x"01000708",
			1325 => x"0e004c04",
			1326 => x"001514f1",
			1327 => x"ffe614f1",
			1328 => x"ff9414f1",
			1329 => x"001114f1",
			1330 => x"08001d0c",
			1331 => x"04003808",
			1332 => x"0a003104",
			1333 => x"000314f1",
			1334 => x"007414f1",
			1335 => x"ffea14f1",
			1336 => x"09002e04",
			1337 => x"ffc714f1",
			1338 => x"000b14f1",
			1339 => x"ff9b14f1",
			1340 => x"0200ae48",
			1341 => x"05004140",
			1342 => x"03001c20",
			1343 => x"05001510",
			1344 => x"0b001004",
			1345 => x"ffcf1585",
			1346 => x"0c001704",
			1347 => x"009a1585",
			1348 => x"0d001304",
			1349 => x"ffd11585",
			1350 => x"001b1585",
			1351 => x"08002304",
			1352 => x"ff4a1585",
			1353 => x"0d001c04",
			1354 => x"00061585",
			1355 => x"08002604",
			1356 => x"00031585",
			1357 => x"fff71585",
			1358 => x"01000a0c",
			1359 => x"08001c08",
			1360 => x"06007704",
			1361 => x"00a71585",
			1362 => x"ffec1585",
			1363 => x"ffeb1585",
			1364 => x"0c001804",
			1365 => x"ff631585",
			1366 => x"00004508",
			1367 => x"0b002004",
			1368 => x"000f1585",
			1369 => x"ffb81585",
			1370 => x"00007f04",
			1371 => x"007b1585",
			1372 => x"fff71585",
			1373 => x"0c001b04",
			1374 => x"ff3d1585",
			1375 => x"00441585",
			1376 => x"ff571585",
			1377 => x"0e006150",
			1378 => x"04001c38",
			1379 => x"03001c24",
			1380 => x"04000e10",
			1381 => x"00002104",
			1382 => x"ff0a1629",
			1383 => x"00005204",
			1384 => x"016f1629",
			1385 => x"07002204",
			1386 => x"fef31629",
			1387 => x"009f1629",
			1388 => x"0a001c10",
			1389 => x"05001208",
			1390 => x"03001004",
			1391 => x"ffc91629",
			1392 => x"003a1629",
			1393 => x"03001a04",
			1394 => x"fea11629",
			1395 => x"fff91629",
			1396 => x"ffe81629",
			1397 => x"01000a04",
			1398 => x"01981629",
			1399 => x"0000940c",
			1400 => x"09002004",
			1401 => x"ffcb1629",
			1402 => x"00003d04",
			1403 => x"ff921629",
			1404 => x"01651629",
			1405 => x"ff121629",
			1406 => x"08001d14",
			1407 => x"06004104",
			1408 => x"00e91629",
			1409 => x"0c001b0c",
			1410 => x"08001604",
			1411 => x"00971629",
			1412 => x"05003704",
			1413 => x"ff801629",
			1414 => x"fe741629",
			1415 => x"00c21629",
			1416 => x"fe561629",
			1417 => x"fe751629",
			1418 => x"0e006164",
			1419 => x"04001430",
			1420 => x"03001a24",
			1421 => x"04000c10",
			1422 => x"08001804",
			1423 => x"013616f7",
			1424 => x"0d001304",
			1425 => x"ff8016f7",
			1426 => x"02006e04",
			1427 => x"00d016f7",
			1428 => x"ff7616f7",
			1429 => x"05001b0c",
			1430 => x"00004f08",
			1431 => x"00003504",
			1432 => x"ff6016f7",
			1433 => x"008516f7",
			1434 => x"fea916f7",
			1435 => x"07002d04",
			1436 => x"00fa16f7",
			1437 => x"ffc316f7",
			1438 => x"01000a04",
			1439 => x"018616f7",
			1440 => x"0d001804",
			1441 => x"000416f7",
			1442 => x"00cc16f7",
			1443 => x"01000a1c",
			1444 => x"0c001b14",
			1445 => x"00006e04",
			1446 => x"00c116f7",
			1447 => x"0f006708",
			1448 => x"0a003104",
			1449 => x"feac16f7",
			1450 => x"ffc916f7",
			1451 => x"08001b04",
			1452 => x"00fb16f7",
			1453 => x"ff1816f7",
			1454 => x"02009904",
			1455 => x"017316f7",
			1456 => x"000516f7",
			1457 => x"0b002714",
			1458 => x"08001b04",
			1459 => x"ffe116f7",
			1460 => x"04001908",
			1461 => x"0a001e04",
			1462 => x"ff6416f7",
			1463 => x"006a16f7",
			1464 => x"0a002704",
			1465 => x"ff8816f7",
			1466 => x"fe8616f7",
			1467 => x"008016f7",
			1468 => x"fe7f16f7",
			1469 => x"00007c18",
			1470 => x"0b00150c",
			1471 => x"01000404",
			1472 => x"002e1769",
			1473 => x"0e002404",
			1474 => x"00021769",
			1475 => x"ffb61769",
			1476 => x"06002808",
			1477 => x"07002304",
			1478 => x"00221769",
			1479 => x"ffc51769",
			1480 => x"00821769",
			1481 => x"0d001314",
			1482 => x"06004d04",
			1483 => x"ffc01769",
			1484 => x"09001704",
			1485 => x"ffda1769",
			1486 => x"0f007808",
			1487 => x"04003104",
			1488 => x"00911769",
			1489 => x"fff51769",
			1490 => x"ffe01769",
			1491 => x"0c001b08",
			1492 => x"01000404",
			1493 => x"00021769",
			1494 => x"ff821769",
			1495 => x"02009904",
			1496 => x"002d1769",
			1497 => x"ffd01769",
			1498 => x"05002b20",
			1499 => x"0000750c",
			1500 => x"0b001204",
			1501 => x"ffe517e5",
			1502 => x"02002004",
			1503 => x"ffef17e5",
			1504 => x"006517e5",
			1505 => x"0f005604",
			1506 => x"ffb117e5",
			1507 => x"09001704",
			1508 => x"ffe617e5",
			1509 => x"0f007a08",
			1510 => x"08001b04",
			1511 => x"005e17e5",
			1512 => x"000217e5",
			1513 => x"ffe817e5",
			1514 => x"0c001b10",
			1515 => x"0e003c04",
			1516 => x"000d17e5",
			1517 => x"08001604",
			1518 => x"000b17e5",
			1519 => x"01000404",
			1520 => x"000017e5",
			1521 => x"ff9c17e5",
			1522 => x"08001d08",
			1523 => x"04003704",
			1524 => x"004317e5",
			1525 => x"fff517e5",
			1526 => x"04002004",
			1527 => x"001017e5",
			1528 => x"ffcb17e5",
			1529 => x"0c001b34",
			1530 => x"0e003a14",
			1531 => x"0b00150c",
			1532 => x"0f002004",
			1533 => x"00411871",
			1534 => x"03001c04",
			1535 => x"ffa01871",
			1536 => x"00051871",
			1537 => x"00002804",
			1538 => x"fff21871",
			1539 => x"00801871",
			1540 => x"0800160c",
			1541 => x"0d001004",
			1542 => x"ffe41871",
			1543 => x"0000af04",
			1544 => x"00401871",
			1545 => x"fff61871",
			1546 => x"0100040c",
			1547 => x"09001d08",
			1548 => x"0d001104",
			1549 => x"ffd71871",
			1550 => x"00471871",
			1551 => x"ffd41871",
			1552 => x"0d001004",
			1553 => x"00011871",
			1554 => x"ff601871",
			1555 => x"0200990c",
			1556 => x"06002808",
			1557 => x"07002304",
			1558 => x"00111871",
			1559 => x"ffc51871",
			1560 => x"00911871",
			1561 => x"01000704",
			1562 => x"00161871",
			1563 => x"ffbe1871",
			1564 => x"0700252c",
			1565 => x"02006b18",
			1566 => x"0c001408",
			1567 => x"0d000f04",
			1568 => x"00711905",
			1569 => x"fe471905",
			1570 => x"05002d0c",
			1571 => x"06003008",
			1572 => x"0f002e04",
			1573 => x"06791905",
			1574 => x"055f1905",
			1575 => x"08101905",
			1576 => x"031e1905",
			1577 => x"01000608",
			1578 => x"0a002704",
			1579 => x"04871905",
			1580 => x"fe461905",
			1581 => x"0f005f08",
			1582 => x"09001f04",
			1583 => x"fe411905",
			1584 => x"ff771905",
			1585 => x"004e1905",
			1586 => x"0200a218",
			1587 => x"00002f04",
			1588 => x"fe421905",
			1589 => x"02008b08",
			1590 => x"0c001b04",
			1591 => x"02261905",
			1592 => x"06b41905",
			1593 => x"08001b04",
			1594 => x"02521905",
			1595 => x"0c001b04",
			1596 => x"fe481905",
			1597 => x"00311905",
			1598 => x"05001c04",
			1599 => x"ff8b1905",
			1600 => x"fe431905",
			1601 => x"07002528",
			1602 => x"02006b14",
			1603 => x"0b001204",
			1604 => x"fe511991",
			1605 => x"05002d0c",
			1606 => x"0c001504",
			1607 => x"01c31991",
			1608 => x"0e002d04",
			1609 => x"03921991",
			1610 => x"04541991",
			1611 => x"00b01991",
			1612 => x"01000608",
			1613 => x"07002104",
			1614 => x"fe3a1991",
			1615 => x"02581991",
			1616 => x"02007404",
			1617 => x"013f1991",
			1618 => x"06005904",
			1619 => x"fe4a1991",
			1620 => x"ff631991",
			1621 => x"0200a218",
			1622 => x"00002f04",
			1623 => x"fe4d1991",
			1624 => x"0a003b10",
			1625 => x"0900240c",
			1626 => x"0c001604",
			1627 => x"fe391991",
			1628 => x"08001c04",
			1629 => x"031a1991",
			1630 => x"ff471991",
			1631 => x"04251991",
			1632 => x"fe281991",
			1633 => x"05001c04",
			1634 => x"ff7d1991",
			1635 => x"fe4c1991",
			1636 => x"08001b28",
			1637 => x"0b001208",
			1638 => x"00009b04",
			1639 => x"ff891a25",
			1640 => x"00221a25",
			1641 => x"05004118",
			1642 => x"0f007914",
			1643 => x"0f005410",
			1644 => x"0f003208",
			1645 => x"00002104",
			1646 => x"fff71a25",
			1647 => x"00aa1a25",
			1648 => x"01000804",
			1649 => x"ff7a1a25",
			1650 => x"00331a25",
			1651 => x"00dc1a25",
			1652 => x"ffb81a25",
			1653 => x"0e004d04",
			1654 => x"00281a25",
			1655 => x"ff951a25",
			1656 => x"0b001910",
			1657 => x"0e003708",
			1658 => x"0a002004",
			1659 => x"ffc11a25",
			1660 => x"00271a25",
			1661 => x"04001204",
			1662 => x"ffff1a25",
			1663 => x"ff191a25",
			1664 => x"02009910",
			1665 => x"06002808",
			1666 => x"07002304",
			1667 => x"00251a25",
			1668 => x"ffab1a25",
			1669 => x"03001704",
			1670 => x"fffc1a25",
			1671 => x"00961a25",
			1672 => x"ff911a25",
			1673 => x"0c001b40",
			1674 => x"0e003a18",
			1675 => x"0b001510",
			1676 => x"00004608",
			1677 => x"0b001204",
			1678 => x"ffdd1ac9",
			1679 => x"005d1ac9",
			1680 => x"03001c04",
			1681 => x"ffa81ac9",
			1682 => x"fff61ac9",
			1683 => x"00002804",
			1684 => x"fff21ac9",
			1685 => x"00861ac9",
			1686 => x"0800160c",
			1687 => x"0d001004",
			1688 => x"ffe31ac9",
			1689 => x"07002904",
			1690 => x"003f1ac9",
			1691 => x"fff81ac9",
			1692 => x"0100040c",
			1693 => x"0b001404",
			1694 => x"ffd11ac9",
			1695 => x"0b001604",
			1696 => x"00461ac9",
			1697 => x"ffdb1ac9",
			1698 => x"0b001908",
			1699 => x"0d001004",
			1700 => x"00011ac9",
			1701 => x"ff511ac9",
			1702 => x"0d001504",
			1703 => x"00131ac9",
			1704 => x"ffe51ac9",
			1705 => x"0200990c",
			1706 => x"06002808",
			1707 => x"07002304",
			1708 => x"00111ac9",
			1709 => x"ffc31ac9",
			1710 => x"00961ac9",
			1711 => x"01000704",
			1712 => x"00161ac9",
			1713 => x"ffbb1ac9",
			1714 => x"0700252c",
			1715 => x"02005810",
			1716 => x"0b001204",
			1717 => x"fe4c1b5d",
			1718 => x"01001008",
			1719 => x"01000404",
			1720 => x"05861b5d",
			1721 => x"04841b5d",
			1722 => x"02bc1b5d",
			1723 => x"01000b14",
			1724 => x"0200a510",
			1725 => x"0a001604",
			1726 => x"fe441b5d",
			1727 => x"05003c08",
			1728 => x"07002104",
			1729 => x"02591b5d",
			1730 => x"055e1b5d",
			1731 => x"fe521b5d",
			1732 => x"fe3a1b5d",
			1733 => x"0b001804",
			1734 => x"fe411b5d",
			1735 => x"ffa41b5d",
			1736 => x"0200a218",
			1737 => x"00002f04",
			1738 => x"fe481b5d",
			1739 => x"0a003b10",
			1740 => x"02008004",
			1741 => x"04bf1b5d",
			1742 => x"08001b04",
			1743 => x"03091b5d",
			1744 => x"0e005604",
			1745 => x"fe3e1b5d",
			1746 => x"01861b5d",
			1747 => x"fe221b5d",
			1748 => x"05001c04",
			1749 => x"ff611b5d",
			1750 => x"fe481b5d",
			1751 => x"0500150c",
			1752 => x"0b001004",
			1753 => x"fff11be9",
			1754 => x"00002104",
			1755 => x"fff21be9",
			1756 => x"00461be9",
			1757 => x"0c001614",
			1758 => x"0800160c",
			1759 => x"0c001304",
			1760 => x"fff11be9",
			1761 => x"06007004",
			1762 => x"000c1be9",
			1763 => x"fffb1be9",
			1764 => x"0e002d04",
			1765 => x"00051be9",
			1766 => x"ffab1be9",
			1767 => x"07002208",
			1768 => x"0a001e04",
			1769 => x"fffd1be9",
			1770 => x"00471be9",
			1771 => x"06004708",
			1772 => x"04001204",
			1773 => x"00031be9",
			1774 => x"ffc51be9",
			1775 => x"0d00130c",
			1776 => x"04002d08",
			1777 => x"0000be04",
			1778 => x"004f1be9",
			1779 => x"fffc1be9",
			1780 => x"ffec1be9",
			1781 => x"02008b04",
			1782 => x"00261be9",
			1783 => x"09002404",
			1784 => x"ffbd1be9",
			1785 => x"00091be9",
			1786 => x"0700273c",
			1787 => x"00007c24",
			1788 => x"0b001510",
			1789 => x"00004608",
			1790 => x"0b001204",
			1791 => x"fe891c9d",
			1792 => x"02491c9d",
			1793 => x"08001904",
			1794 => x"00791c9d",
			1795 => x"fe3d1c9d",
			1796 => x"00002804",
			1797 => x"fe1c1c9d",
			1798 => x"08001d08",
			1799 => x"05002304",
			1800 => x"01d11c9d",
			1801 => x"02961c9d",
			1802 => x"05001f04",
			1803 => x"01de1c9d",
			1804 => x"006d1c9d",
			1805 => x"0100060c",
			1806 => x"03002d08",
			1807 => x"0200af04",
			1808 => x"01751c9d",
			1809 => x"fe691c9d",
			1810 => x"fe5f1c9d",
			1811 => x"0a003808",
			1812 => x"0f006104",
			1813 => x"fe501c9d",
			1814 => x"ff411c9d",
			1815 => x"00801c9d",
			1816 => x"0000aa1c",
			1817 => x"0e00340c",
			1818 => x"07002808",
			1819 => x"01000a04",
			1820 => x"fe861c9d",
			1821 => x"ffb51c9d",
			1822 => x"fe5e1c9d",
			1823 => x"03003a0c",
			1824 => x"07002a08",
			1825 => x"01000b04",
			1826 => x"00c01c9d",
			1827 => x"fec91c9d",
			1828 => x"023c1c9d",
			1829 => x"fe351c9d",
			1830 => x"fe5e1c9d",
			1831 => x"0c001510",
			1832 => x"06002204",
			1833 => x"00281d31",
			1834 => x"08001608",
			1835 => x"08001504",
			1836 => x"fff81d31",
			1837 => x"00001d31",
			1838 => x"ff901d31",
			1839 => x"0e003914",
			1840 => x"00002804",
			1841 => x"ffe71d31",
			1842 => x"0000750c",
			1843 => x"03001308",
			1844 => x"0b001604",
			1845 => x"fff41d31",
			1846 => x"000e1d31",
			1847 => x"007e1d31",
			1848 => x"fff31d31",
			1849 => x"0f005208",
			1850 => x"05003004",
			1851 => x"ff981d31",
			1852 => x"00091d31",
			1853 => x"0d00130c",
			1854 => x"0f007808",
			1855 => x"04003104",
			1856 => x"00881d31",
			1857 => x"fff51d31",
			1858 => x"ffed1d31",
			1859 => x"0c001b08",
			1860 => x"01000404",
			1861 => x"00021d31",
			1862 => x"ff991d31",
			1863 => x"0a003708",
			1864 => x"0000be04",
			1865 => x"004f1d31",
			1866 => x"fff51d31",
			1867 => x"ffdf1d31",
			1868 => x"01000a30",
			1869 => x"0e005020",
			1870 => x"0b001204",
			1871 => x"ff981ded",
			1872 => x"08001d14",
			1873 => x"0500210c",
			1874 => x"02005808",
			1875 => x"00002104",
			1876 => x"ffe11ded",
			1877 => x"00b31ded",
			1878 => x"ffc61ded",
			1879 => x"02009704",
			1880 => x"00c01ded",
			1881 => x"fff91ded",
			1882 => x"00004904",
			1883 => x"000a1ded",
			1884 => x"ffce1ded",
			1885 => x"02009704",
			1886 => x"ff3b1ded",
			1887 => x"05003c08",
			1888 => x"06007204",
			1889 => x"00e21ded",
			1890 => x"ff9d1ded",
			1891 => x"ff611ded",
			1892 => x"0e003d20",
			1893 => x"01001014",
			1894 => x"0b001608",
			1895 => x"00004804",
			1896 => x"fffe1ded",
			1897 => x"ffc41ded",
			1898 => x"07002708",
			1899 => x"00007c04",
			1900 => x"00a21ded",
			1901 => x"ffeb1ded",
			1902 => x"ffe41ded",
			1903 => x"04001708",
			1904 => x"00003904",
			1905 => x"ffea1ded",
			1906 => x"002b1ded",
			1907 => x"ff9d1ded",
			1908 => x"09003008",
			1909 => x"08001804",
			1910 => x"00281ded",
			1911 => x"fefd1ded",
			1912 => x"0a003b04",
			1913 => x"00591ded",
			1914 => x"ffe71ded",
			1915 => x"0200ae24",
			1916 => x"05000904",
			1917 => x"01ee1e39",
			1918 => x"0c001304",
			1919 => x"fe711e39",
			1920 => x"00002504",
			1921 => x"fe891e39",
			1922 => x"02005008",
			1923 => x"01001004",
			1924 => x"01901e39",
			1925 => x"00c01e39",
			1926 => x"01000a08",
			1927 => x"0c001b04",
			1928 => x"003c1e39",
			1929 => x"01711e39",
			1930 => x"0c001804",
			1931 => x"fe781e39",
			1932 => x"ffec1e39",
			1933 => x"fe6c1e39",
			1934 => x"0700252c",
			1935 => x"02006b18",
			1936 => x"0b001204",
			1937 => x"fe571ed5",
			1938 => x"0e003810",
			1939 => x"0100100c",
			1940 => x"0a000a04",
			1941 => x"04241ed5",
			1942 => x"0b001504",
			1943 => x"018d1ed5",
			1944 => x"031d1ed5",
			1945 => x"01c51ed5",
			1946 => x"ffe01ed5",
			1947 => x"08001b10",
			1948 => x"0200a50c",
			1949 => x"06004e04",
			1950 => x"ff821ed5",
			1951 => x"05002504",
			1952 => x"047a1ed5",
			1953 => x"00911ed5",
			1954 => x"fe4d1ed5",
			1955 => x"fe4d1ed5",
			1956 => x"0200a21c",
			1957 => x"00002f04",
			1958 => x"fe511ed5",
			1959 => x"02008b08",
			1960 => x"04001904",
			1961 => x"037a1ed5",
			1962 => x"01301ed5",
			1963 => x"0400320c",
			1964 => x"04001a04",
			1965 => x"fe3a1ed5",
			1966 => x"01000c04",
			1967 => x"03771ed5",
			1968 => x"ff8d1ed5",
			1969 => x"fe481ed5",
			1970 => x"05001c04",
			1971 => x"ffe41ed5",
			1972 => x"fe501ed5",
			1973 => x"0c001510",
			1974 => x"06002204",
			1975 => x"00291f71",
			1976 => x"08001608",
			1977 => x"08001504",
			1978 => x"fff71f71",
			1979 => x"00001f71",
			1980 => x"ff8d1f71",
			1981 => x"0e003914",
			1982 => x"00002804",
			1983 => x"ffe71f71",
			1984 => x"0000750c",
			1985 => x"03001308",
			1986 => x"0b001604",
			1987 => x"fff31f71",
			1988 => x"000e1f71",
			1989 => x"00831f71",
			1990 => x"fff31f71",
			1991 => x"0f00520c",
			1992 => x"0c001904",
			1993 => x"ff941f71",
			1994 => x"0c001c04",
			1995 => x"002a1f71",
			1996 => x"ffdc1f71",
			1997 => x"0d00130c",
			1998 => x"0f007808",
			1999 => x"04003104",
			2000 => x"008a1f71",
			2001 => x"fff51f71",
			2002 => x"ffed1f71",
			2003 => x"0c001b08",
			2004 => x"01000404",
			2005 => x"00021f71",
			2006 => x"ff961f71",
			2007 => x"0a003708",
			2008 => x"0000be04",
			2009 => x"00501f71",
			2010 => x"fff51f71",
			2011 => x"ffde1f71",
			2012 => x"0e00391c",
			2013 => x"0b00150c",
			2014 => x"06002204",
			2015 => x"00712035",
			2016 => x"00004604",
			2017 => x"fff62035",
			2018 => x"ff3d2035",
			2019 => x"07002308",
			2020 => x"00007504",
			2021 => x"00fe2035",
			2022 => x"ffdd2035",
			2023 => x"06002904",
			2024 => x"ff7e2035",
			2025 => x"00392035",
			2026 => x"0c001b34",
			2027 => x"08001814",
			2028 => x"03001f08",
			2029 => x"06008004",
			2030 => x"00692035",
			2031 => x"fff92035",
			2032 => x"01000a08",
			2033 => x"01000304",
			2034 => x"00072035",
			2035 => x"ff8b2035",
			2036 => x"002b2035",
			2037 => x"05002510",
			2038 => x"05002308",
			2039 => x"0d001104",
			2040 => x"00032035",
			2041 => x"ff482035",
			2042 => x"0000d604",
			2043 => x"00712035",
			2044 => x"fff32035",
			2045 => x"0c001a04",
			2046 => x"fed22035",
			2047 => x"0d001708",
			2048 => x"08001b04",
			2049 => x"002a2035",
			2050 => x"ff802035",
			2051 => x"00282035",
			2052 => x"0d001608",
			2053 => x"04003704",
			2054 => x"00ca2035",
			2055 => x"ffc82035",
			2056 => x"09003004",
			2057 => x"ff702035",
			2058 => x"0a003b04",
			2059 => x"004b2035",
			2060 => x"ffe22035",
			2061 => x"02008020",
			2062 => x"05002b18",
			2063 => x"0b001204",
			2064 => x"ffd320d1",
			2065 => x"02002004",
			2066 => x"ffe620d1",
			2067 => x"0000750c",
			2068 => x"07002e08",
			2069 => x"04000704",
			2070 => x"000220d1",
			2071 => x"009c20d1",
			2072 => x"fffb20d1",
			2073 => x"000320d1",
			2074 => x"09001e04",
			2075 => x"ffc220d1",
			2076 => x"002020d1",
			2077 => x"0c001b20",
			2078 => x"0d00131c",
			2079 => x"09001704",
			2080 => x"ffb320d1",
			2081 => x"0800160c",
			2082 => x"04001e04",
			2083 => x"ffd820d1",
			2084 => x"03002d04",
			2085 => x"001420d1",
			2086 => x"fffa20d1",
			2087 => x"0a002808",
			2088 => x"0200ae04",
			2089 => x"006920d1",
			2090 => x"fff920d1",
			2091 => x"ffe820d1",
			2092 => x"ff6c20d1",
			2093 => x"01000a08",
			2094 => x"05004704",
			2095 => x"006420d1",
			2096 => x"fff120d1",
			2097 => x"09003a04",
			2098 => x"ffb820d1",
			2099 => x"001920d1",
			2100 => x"0200ae34",
			2101 => x"08001d1c",
			2102 => x"05004618",
			2103 => x"0c001104",
			2104 => x"fe8c213d",
			2105 => x"0a000a04",
			2106 => x"01bb213d",
			2107 => x"0c001508",
			2108 => x"08001804",
			2109 => x"002d213d",
			2110 => x"fe90213d",
			2111 => x"00002804",
			2112 => x"fed2213d",
			2113 => x"00c5213d",
			2114 => x"fe9d213d",
			2115 => x"04001c14",
			2116 => x"02003808",
			2117 => x"05001004",
			2118 => x"0015213d",
			2119 => x"feb3213d",
			2120 => x"00009408",
			2121 => x"0c001a04",
			2122 => x"ff56213d",
			2123 => x"017c213d",
			2124 => x"fee0213d",
			2125 => x"fe17213d",
			2126 => x"fe6f213d",
			2127 => x"0c001304",
			2128 => x"ffba21c1",
			2129 => x"08001b20",
			2130 => x"05004118",
			2131 => x"0f007914",
			2132 => x"0a00140c",
			2133 => x"00005208",
			2134 => x"00002504",
			2135 => x"fffb21c1",
			2136 => x"002121c1",
			2137 => x"ffd521c1",
			2138 => x"05001704",
			2139 => x"ffff21c1",
			2140 => x"006f21c1",
			2141 => x"ffe721c1",
			2142 => x"0b001904",
			2143 => x"ffcb21c1",
			2144 => x"001021c1",
			2145 => x"0b001910",
			2146 => x"0e00380c",
			2147 => x"07001d04",
			2148 => x"fff121c1",
			2149 => x"00003d04",
			2150 => x"fff721c1",
			2151 => x"001a21c1",
			2152 => x"ff9d21c1",
			2153 => x"0200990c",
			2154 => x"06002808",
			2155 => x"07002304",
			2156 => x"000d21c1",
			2157 => x"ffd621c1",
			2158 => x"004f21c1",
			2159 => x"ffd821c1",
			2160 => x"0200ae34",
			2161 => x"00002504",
			2162 => x"fe83222d",
			2163 => x"04001414",
			2164 => x"0b001308",
			2165 => x"0d000f04",
			2166 => x"00fd222d",
			2167 => x"fe57222d",
			2168 => x"00006504",
			2169 => x"0198222d",
			2170 => x"06004e04",
			2171 => x"fe8b222d",
			2172 => x"01dd222d",
			2173 => x"08001d10",
			2174 => x"0c001b0c",
			2175 => x"05004108",
			2176 => x"0c001604",
			2177 => x"ff28222d",
			2178 => x"00be222d",
			2179 => x"fe6e222d",
			2180 => x"016b222d",
			2181 => x"04001c08",
			2182 => x"0a002704",
			2183 => x"ff07222d",
			2184 => x"0161222d",
			2185 => x"fe1e222d",
			2186 => x"fe6a222d",
			2187 => x"0f006e40",
			2188 => x"0b001928",
			2189 => x"08001b18",
			2190 => x"05004114",
			2191 => x"0c001104",
			2192 => x"ffcc22b1",
			2193 => x"0f005408",
			2194 => x"0f003204",
			2195 => x"006422b1",
			2196 => x"ffc522b1",
			2197 => x"0000b004",
			2198 => x"008e22b1",
			2199 => x"fffb22b1",
			2200 => x"ffbf22b1",
			2201 => x"0f003c0c",
			2202 => x"0a002008",
			2203 => x"0a000b04",
			2204 => x"000222b1",
			2205 => x"ffe722b1",
			2206 => x"001322b1",
			2207 => x"ff9722b1",
			2208 => x"06002808",
			2209 => x"07002304",
			2210 => x"001322b1",
			2211 => x"ffcb22b1",
			2212 => x"0300390c",
			2213 => x"0000aa08",
			2214 => x"0a002104",
			2215 => x"000722b1",
			2216 => x"008b22b1",
			2217 => x"fff522b1",
			2218 => x"ffe022b1",
			2219 => x"ff9722b1",
			2220 => x"0200a548",
			2221 => x"0c001b30",
			2222 => x"0800180c",
			2223 => x"06004508",
			2224 => x"02004604",
			2225 => x"00992345",
			2226 => x"ff982345",
			2227 => x"00c42345",
			2228 => x"0e003810",
			2229 => x"0b001508",
			2230 => x"06002304",
			2231 => x"00302345",
			2232 => x"ff532345",
			2233 => x"00002804",
			2234 => x"ffcf2345",
			2235 => x"00f62345",
			2236 => x"0200940c",
			2237 => x"04001404",
			2238 => x"fff62345",
			2239 => x"0a003104",
			2240 => x"fec62345",
			2241 => x"ffc72345",
			2242 => x"08001b04",
			2243 => x"00a42345",
			2244 => x"ff782345",
			2245 => x"06002808",
			2246 => x"07002304",
			2247 => x"00342345",
			2248 => x"ff712345",
			2249 => x"0a002a08",
			2250 => x"00008b04",
			2251 => x"00ab2345",
			2252 => x"ff7c2345",
			2253 => x"00007804",
			2254 => x"001c2345",
			2255 => x"010f2345",
			2256 => x"fee02345",
			2257 => x"05002b34",
			2258 => x"0b001208",
			2259 => x"09001704",
			2260 => x"ff802401",
			2261 => x"002f2401",
			2262 => x"06007028",
			2263 => x"0a001b14",
			2264 => x"0000520c",
			2265 => x"07002404",
			2266 => x"00852401",
			2267 => x"06002204",
			2268 => x"ffd42401",
			2269 => x"00082401",
			2270 => x"01000e04",
			2271 => x"ff902401",
			2272 => x"00082401",
			2273 => x"00003504",
			2274 => x"fff72401",
			2275 => x"00007508",
			2276 => x"07001c04",
			2277 => x"000a2401",
			2278 => x"00cc2401",
			2279 => x"09001d04",
			2280 => x"00692401",
			2281 => x"ffe52401",
			2282 => x"ffaf2401",
			2283 => x"0c001b1c",
			2284 => x"08001608",
			2285 => x"03002d04",
			2286 => x"003b2401",
			2287 => x"fff72401",
			2288 => x"0f004304",
			2289 => x"fff82401",
			2290 => x"0b001908",
			2291 => x"0d001104",
			2292 => x"fffa2401",
			2293 => x"ff132401",
			2294 => x"0d001504",
			2295 => x"00182401",
			2296 => x"ffd62401",
			2297 => x"08001d08",
			2298 => x"04003704",
			2299 => x"00af2401",
			2300 => x"ffe22401",
			2301 => x"04001f04",
			2302 => x"00192401",
			2303 => x"ff892401",
			2304 => x"0200ae40",
			2305 => x"0c001614",
			2306 => x"00004608",
			2307 => x"0b001204",
			2308 => x"ffcb2485",
			2309 => x"00a12485",
			2310 => x"08001604",
			2311 => x"002b2485",
			2312 => x"00009f04",
			2313 => x"ff072485",
			2314 => x"00002485",
			2315 => x"05004628",
			2316 => x"0a001b10",
			2317 => x"00006b08",
			2318 => x"00002804",
			2319 => x"ffb62485",
			2320 => x"006c2485",
			2321 => x"01000e04",
			2322 => x"ff872485",
			2323 => x"fffd2485",
			2324 => x"01000b0c",
			2325 => x"08001d08",
			2326 => x"05002104",
			2327 => x"00292485",
			2328 => x"00de2485",
			2329 => x"ffd72485",
			2330 => x"05003108",
			2331 => x"00008804",
			2332 => x"00882485",
			2333 => x"fffb2485",
			2334 => x"ff7f2485",
			2335 => x"ff652485",
			2336 => x"ff262485",
			2337 => x"0200a530",
			2338 => x"02002004",
			2339 => x"fe6824e9",
			2340 => x"0f003314",
			2341 => x"05002110",
			2342 => x"0b001204",
			2343 => x"feaa24e9",
			2344 => x"07002e08",
			2345 => x"02004e04",
			2346 => x"01b224e9",
			2347 => x"00f024e9",
			2348 => x"fed024e9",
			2349 => x"ff9424e9",
			2350 => x"05004614",
			2351 => x"07001d04",
			2352 => x"fe6024e9",
			2353 => x"0c001a08",
			2354 => x"08001604",
			2355 => x"014424e9",
			2356 => x"ffbe24e9",
			2357 => x"0c001c04",
			2358 => x"018824e9",
			2359 => x"005524e9",
			2360 => x"fe7124e9",
			2361 => x"fe6424e9",
			2362 => x"0e005040",
			2363 => x"08001d28",
			2364 => x"0b001204",
			2365 => x"ff5825b5",
			2366 => x"0200921c",
			2367 => x"03001510",
			2368 => x"07001b08",
			2369 => x"02003104",
			2370 => x"00ca25b5",
			2371 => x"000025b5",
			2372 => x"0a000a04",
			2373 => x"001925b5",
			2374 => x"ff5c25b5",
			2375 => x"01000b08",
			2376 => x"04003104",
			2377 => x"010125b5",
			2378 => x"002225b5",
			2379 => x"fff425b5",
			2380 => x"0e004b04",
			2381 => x"ff5a25b5",
			2382 => x"009125b5",
			2383 => x"04001c14",
			2384 => x"0a002110",
			2385 => x"0500160c",
			2386 => x"00006e08",
			2387 => x"00003504",
			2388 => x"ffec25b5",
			2389 => x"004c25b5",
			2390 => x"ffd325b5",
			2391 => x"ff8925b5",
			2392 => x"007e25b5",
			2393 => x"ff1725b5",
			2394 => x"0a002810",
			2395 => x"0c001608",
			2396 => x"0d000f04",
			2397 => x"006125b5",
			2398 => x"ff3025b5",
			2399 => x"0f007d04",
			2400 => x"00e125b5",
			2401 => x"ffd425b5",
			2402 => x"09003a14",
			2403 => x"08001608",
			2404 => x"0d001104",
			2405 => x"001d25b5",
			2406 => x"ffe025b5",
			2407 => x"0c001b04",
			2408 => x"fec625b5",
			2409 => x"0c001c04",
			2410 => x"000225b5",
			2411 => x"ff7725b5",
			2412 => x"004225b5",
			2413 => x"0e005b50",
			2414 => x"0b001930",
			2415 => x"09001f28",
			2416 => x"0c001818",
			2417 => x"05002b10",
			2418 => x"0c001308",
			2419 => x"06002304",
			2420 => x"00352661",
			2421 => x"ff362661",
			2422 => x"0f004b04",
			2423 => x"00002661",
			2424 => x"00c22661",
			2425 => x"01000704",
			2426 => x"fff32661",
			2427 => x"ff0d2661",
			2428 => x"0000a60c",
			2429 => x"03001a08",
			2430 => x"05001004",
			2431 => x"00052661",
			2432 => x"ffe82661",
			2433 => x"00ee2661",
			2434 => x"ffd82661",
			2435 => x"0c001b04",
			2436 => x"ff082661",
			2437 => x"ffe32661",
			2438 => x"01000a0c",
			2439 => x"0a001908",
			2440 => x"05001004",
			2441 => x"00062661",
			2442 => x"fff22661",
			2443 => x"00f92661",
			2444 => x"0000810c",
			2445 => x"06002808",
			2446 => x"07002304",
			2447 => x"00342661",
			2448 => x"ff802661",
			2449 => x"00ad2661",
			2450 => x"07002d04",
			2451 => x"ff682661",
			2452 => x"00092661",
			2453 => x"08003504",
			2454 => x"fed72661",
			2455 => x"00212661",
			2456 => x"0e005d44",
			2457 => x"0c001308",
			2458 => x"06002404",
			2459 => x"001226f5",
			2460 => x"ffad26f5",
			2461 => x"05002b20",
			2462 => x"00002808",
			2463 => x"03000c04",
			2464 => x"000126f5",
			2465 => x"ffe126f5",
			2466 => x"0000a10c",
			2467 => x"0a001608",
			2468 => x"0a000a04",
			2469 => x"003426f5",
			2470 => x"ffdc26f5",
			2471 => x"009e26f5",
			2472 => x"07002908",
			2473 => x"07002504",
			2474 => x"000426f5",
			2475 => x"ffe826f5",
			2476 => x"001026f5",
			2477 => x"0c001b10",
			2478 => x"0f004304",
			2479 => x"001926f5",
			2480 => x"06006104",
			2481 => x"ff8326f5",
			2482 => x"0d001304",
			2483 => x"001e26f5",
			2484 => x"ffeb26f5",
			2485 => x"0d001704",
			2486 => x"007826f5",
			2487 => x"07003004",
			2488 => x"ffc826f5",
			2489 => x"000326f5",
			2490 => x"07002704",
			2491 => x"fffb26f5",
			2492 => x"ff9b26f5",
			2493 => x"0200ae34",
			2494 => x"02002004",
			2495 => x"fe5d2761",
			2496 => x"00005c14",
			2497 => x"0b002010",
			2498 => x"0b001204",
			2499 => x"fe962761",
			2500 => x"01000e08",
			2501 => x"02002d04",
			2502 => x"023e2761",
			2503 => x"01a92761",
			2504 => x"01022761",
			2505 => x"ff932761",
			2506 => x"05004618",
			2507 => x"05001b08",
			2508 => x"06004c04",
			2509 => x"fe5b2761",
			2510 => x"ffe12761",
			2511 => x"08001d08",
			2512 => x"0c001604",
			2513 => x"fff02761",
			2514 => x"015e2761",
			2515 => x"04001e04",
			2516 => x"00e22761",
			2517 => x"fe472761",
			2518 => x"fe632761",
			2519 => x"fe622761",
			2520 => x"0e005d40",
			2521 => x"0c001308",
			2522 => x"0f002504",
			2523 => x"001327ed",
			2524 => x"ffb227ed",
			2525 => x"05004130",
			2526 => x"0f00551c",
			2527 => x"02008010",
			2528 => x"0b001508",
			2529 => x"02004c04",
			2530 => x"003d27ed",
			2531 => x"ffca27ed",
			2532 => x"00002804",
			2533 => x"ffdc27ed",
			2534 => x"007127ed",
			2535 => x"0d001504",
			2536 => x"ff9b27ed",
			2537 => x"0d001704",
			2538 => x"001627ed",
			2539 => x"ffe727ed",
			2540 => x"08001b08",
			2541 => x"0000b004",
			2542 => x"00a627ed",
			2543 => x"fffb27ed",
			2544 => x"08002308",
			2545 => x"00009f04",
			2546 => x"ffd527ed",
			2547 => x"000b27ed",
			2548 => x"001d27ed",
			2549 => x"0c001b04",
			2550 => x"ffa027ed",
			2551 => x"002a27ed",
			2552 => x"0a002004",
			2553 => x"000127ed",
			2554 => x"ffa227ed",
			2555 => x"0200ae40",
			2556 => x"0c001308",
			2557 => x"0a001204",
			2558 => x"00282871",
			2559 => x"fe612871",
			2560 => x"0400141c",
			2561 => x"00002504",
			2562 => x"fe972871",
			2563 => x"03001a0c",
			2564 => x"00005204",
			2565 => x"018d2871",
			2566 => x"06004904",
			2567 => x"fe862871",
			2568 => x"00672871",
			2569 => x"0a002004",
			2570 => x"01df2871",
			2571 => x"0a002304",
			2572 => x"00b82871",
			2573 => x"01752871",
			2574 => x"08001d10",
			2575 => x"0c001b0c",
			2576 => x"05004108",
			2577 => x"0c001804",
			2578 => x"ffc32871",
			2579 => x"00f62871",
			2580 => x"fe732871",
			2581 => x"01542871",
			2582 => x"04001c08",
			2583 => x"0a002704",
			2584 => x"fee72871",
			2585 => x"01552871",
			2586 => x"fe2a2871",
			2587 => x"fe6b2871",
			2588 => x"05002b40",
			2589 => x"0b001208",
			2590 => x"09001704",
			2591 => x"ff7a2945",
			2592 => x"00302945",
			2593 => x"06007034",
			2594 => x"0a001b1c",
			2595 => x"05000f0c",
			2596 => x"00002104",
			2597 => x"fff32945",
			2598 => x"00005e04",
			2599 => x"00842945",
			2600 => x"fffa2945",
			2601 => x"03001a08",
			2602 => x"08002404",
			2603 => x"ff952945",
			2604 => x"00052945",
			2605 => x"08002604",
			2606 => x"000b2945",
			2607 => x"fffc2945",
			2608 => x"09001e08",
			2609 => x"07001c04",
			2610 => x"00072945",
			2611 => x"00b82945",
			2612 => x"00007508",
			2613 => x"00003d04",
			2614 => x"fff72945",
			2615 => x"00672945",
			2616 => x"07002a04",
			2617 => x"ffb12945",
			2618 => x"00432945",
			2619 => x"ffac2945",
			2620 => x"0c001b1c",
			2621 => x"08001608",
			2622 => x"0000f204",
			2623 => x"003a2945",
			2624 => x"fffb2945",
			2625 => x"0b00190c",
			2626 => x"06004004",
			2627 => x"ffde2945",
			2628 => x"0d001104",
			2629 => x"fff92945",
			2630 => x"ff092945",
			2631 => x"0f006c04",
			2632 => x"00182945",
			2633 => x"fff02945",
			2634 => x"08001d08",
			2635 => x"04003704",
			2636 => x"00b72945",
			2637 => x"ffe12945",
			2638 => x"04001f04",
			2639 => x"00192945",
			2640 => x"ff842945",
			2641 => x"0e006150",
			2642 => x"04001424",
			2643 => x"03001a20",
			2644 => x"04000c10",
			2645 => x"00002104",
			2646 => x"fef229e9",
			2647 => x"00005204",
			2648 => x"019d29e9",
			2649 => x"0a001104",
			2650 => x"fee229e9",
			2651 => x"00da29e9",
			2652 => x"07002008",
			2653 => x"0a001404",
			2654 => x"ff1929e9",
			2655 => x"00e529e9",
			2656 => x"08002404",
			2657 => x"fe8629e9",
			2658 => x"005429e9",
			2659 => x"019f29e9",
			2660 => x"08001d1c",
			2661 => x"0c001a10",
			2662 => x"0500410c",
			2663 => x"0c001404",
			2664 => x"fece29e9",
			2665 => x"0e003904",
			2666 => x"016129e9",
			2667 => x"000529e9",
			2668 => x"fe7e29e9",
			2669 => x"04003808",
			2670 => x"05002c04",
			2671 => x"004429e9",
			2672 => x"01a229e9",
			2673 => x"fedc29e9",
			2674 => x"04001c0c",
			2675 => x"0a002708",
			2676 => x"01000c04",
			2677 => x"ffbf29e9",
			2678 => x"feda29e9",
			2679 => x"014529e9",
			2680 => x"fe2b29e9",
			2681 => x"fe7029e9",
			2682 => x"0000aa3c",
			2683 => x"02002004",
			2684 => x"fe572a6d",
			2685 => x"00005c18",
			2686 => x"0b001204",
			2687 => x"fe7a2a6d",
			2688 => x"0100100c",
			2689 => x"01000504",
			2690 => x"02602a6d",
			2691 => x"01000e04",
			2692 => x"01b92a6d",
			2693 => x"013d2a6d",
			2694 => x"04001804",
			2695 => x"01632a6d",
			2696 => x"fe342a6d",
			2697 => x"0500461c",
			2698 => x"08001d10",
			2699 => x"05001808",
			2700 => x"04000c04",
			2701 => x"ff672a6d",
			2702 => x"fe442a6d",
			2703 => x"0c001804",
			2704 => x"00682a6d",
			2705 => x"01b92a6d",
			2706 => x"04001d08",
			2707 => x"08002204",
			2708 => x"fe792a6d",
			2709 => x"019a2a6d",
			2710 => x"fe382a6d",
			2711 => x"fe5e2a6d",
			2712 => x"05001c04",
			2713 => x"007b2a6d",
			2714 => x"fe602a6d",
			2715 => x"0200a53c",
			2716 => x"02002004",
			2717 => x"fe6c2ae9",
			2718 => x"02006b18",
			2719 => x"05002d14",
			2720 => x"0b001204",
			2721 => x"fea72ae9",
			2722 => x"0b001508",
			2723 => x"08001b04",
			2724 => x"019b2ae9",
			2725 => x"fe9d2ae9",
			2726 => x"00002804",
			2727 => x"feb22ae9",
			2728 => x"01ac2ae9",
			2729 => x"ff7f2ae9",
			2730 => x"0b001910",
			2731 => x"08001b0c",
			2732 => x"06004e04",
			2733 => x"fec32ae9",
			2734 => x"04002904",
			2735 => x"01162ae9",
			2736 => x"fe6e2ae9",
			2737 => x"fe622ae9",
			2738 => x"0a002708",
			2739 => x"03001604",
			2740 => x"ffe02ae9",
			2741 => x"fea02ae9",
			2742 => x"03003a04",
			2743 => x"01a62ae9",
			2744 => x"fea52ae9",
			2745 => x"fe652ae9",
			2746 => x"0e00614c",
			2747 => x"01000a28",
			2748 => x"04003320",
			2749 => x"0b001204",
			2750 => x"ff532b85",
			2751 => x"08001d10",
			2752 => x"0b001908",
			2753 => x"03002c04",
			2754 => x"00dc2b85",
			2755 => x"fefc2b85",
			2756 => x"00002f04",
			2757 => x"ffb82b85",
			2758 => x"01872b85",
			2759 => x"00004f08",
			2760 => x"00001b04",
			2761 => x"ffd72b85",
			2762 => x"00a22b85",
			2763 => x"fefc2b85",
			2764 => x"07002404",
			2765 => x"00662b85",
			2766 => x"fea52b85",
			2767 => x"0c001808",
			2768 => x"04001204",
			2769 => x"ffcd2b85",
			2770 => x"fe882b85",
			2771 => x"07002308",
			2772 => x"02006b04",
			2773 => x"01742b85",
			2774 => x"002b2b85",
			2775 => x"06002a04",
			2776 => x"fe642b85",
			2777 => x"00009408",
			2778 => x"0a002f04",
			2779 => x"012a2b85",
			2780 => x"00552b85",
			2781 => x"0f006b04",
			2782 => x"fe962b85",
			2783 => x"00962b85",
			2784 => x"fe782b85",
			2785 => x"0200ae44",
			2786 => x"02002004",
			2787 => x"fe642c11",
			2788 => x"05002b24",
			2789 => x"00007514",
			2790 => x"0b001204",
			2791 => x"fe812c11",
			2792 => x"04001108",
			2793 => x"06001f04",
			2794 => x"021b2c11",
			2795 => x"01982c11",
			2796 => x"0b001504",
			2797 => x"ffdc2c11",
			2798 => x"018b2c11",
			2799 => x"0f005404",
			2800 => x"fe4a2c11",
			2801 => x"06007008",
			2802 => x"08001b04",
			2803 => x"01a02c11",
			2804 => x"00282c11",
			2805 => x"fe7e2c11",
			2806 => x"08001d10",
			2807 => x"0c001a08",
			2808 => x"04002b04",
			2809 => x"00252c11",
			2810 => x"fe602c11",
			2811 => x"04003804",
			2812 => x"02182c11",
			2813 => x"feb12c11",
			2814 => x"07002c08",
			2815 => x"07002504",
			2816 => x"fd9a2c11",
			2817 => x"fe622c11",
			2818 => x"ff162c11",
			2819 => x"fe642c11",
			2820 => x"0e006158",
			2821 => x"04001424",
			2822 => x"0c001104",
			2823 => x"fee32cc7",
			2824 => x"02002004",
			2825 => x"ff222cc7",
			2826 => x"03001a10",
			2827 => x"00005208",
			2828 => x"05001304",
			2829 => x"015d2cc7",
			2830 => x"00432cc7",
			2831 => x"0f004f04",
			2832 => x"fed52cc7",
			2833 => x"008d2cc7",
			2834 => x"01000a04",
			2835 => x"017b2cc7",
			2836 => x"01000c04",
			2837 => x"00092cc7",
			2838 => x"00ca2cc7",
			2839 => x"0c001a18",
			2840 => x"0d001310",
			2841 => x"05002304",
			2842 => x"ff152cc7",
			2843 => x"03002d08",
			2844 => x"0c001604",
			2845 => x"ffa82cc7",
			2846 => x"01522cc7",
			2847 => x"fee92cc7",
			2848 => x"01000604",
			2849 => x"ffea2cc7",
			2850 => x"fe9a2cc7",
			2851 => x"00004508",
			2852 => x"0d001a04",
			2853 => x"002b2cc7",
			2854 => x"feb12cc7",
			2855 => x"02009204",
			2856 => x"014b2cc7",
			2857 => x"06006108",
			2858 => x"09002404",
			2859 => x"feeb2cc7",
			2860 => x"00822cc7",
			2861 => x"04003904",
			2862 => x"010e2cc7",
			2863 => x"ff7b2cc7",
			2864 => x"fe832cc7",
			2865 => x"00007c1c",
			2866 => x"0c001710",
			2867 => x"0e002c08",
			2868 => x"0b001204",
			2869 => x"ffc92d49",
			2870 => x"00812d49",
			2871 => x"0f004204",
			2872 => x"ff732d49",
			2873 => x"00172d49",
			2874 => x"06002808",
			2875 => x"07002304",
			2876 => x"002a2d49",
			2877 => x"ffaf2d49",
			2878 => x"00ab2d49",
			2879 => x"01000614",
			2880 => x"0e005208",
			2881 => x"07002304",
			2882 => x"fff52d49",
			2883 => x"00792d49",
			2884 => x"0200a104",
			2885 => x"ffa42d49",
			2886 => x"0200ae04",
			2887 => x"004a2d49",
			2888 => x"ffe42d49",
			2889 => x"0b002f10",
			2890 => x"0e004308",
			2891 => x"06004004",
			2892 => x"fff02d49",
			2893 => x"00242d49",
			2894 => x"08001604",
			2895 => x"001a2d49",
			2896 => x"ff522d49",
			2897 => x"00272d49",
			2898 => x"05002b24",
			2899 => x"00007510",
			2900 => x"0b001204",
			2901 => x"ffe52dcd",
			2902 => x"02002004",
			2903 => x"ffef2dcd",
			2904 => x"04000704",
			2905 => x"00032dcd",
			2906 => x"00622dcd",
			2907 => x"0f005604",
			2908 => x"ffb42dcd",
			2909 => x"09001704",
			2910 => x"ffe62dcd",
			2911 => x"0f007a08",
			2912 => x"08001b04",
			2913 => x"005b2dcd",
			2914 => x"00012dcd",
			2915 => x"ffe82dcd",
			2916 => x"0c001b10",
			2917 => x"0e003c04",
			2918 => x"000c2dcd",
			2919 => x"08001604",
			2920 => x"000b2dcd",
			2921 => x"01000404",
			2922 => x"00002dcd",
			2923 => x"ff9f2dcd",
			2924 => x"08001d08",
			2925 => x"04003704",
			2926 => x"00422dcd",
			2927 => x"fff52dcd",
			2928 => x"04002004",
			2929 => x"00102dcd",
			2930 => x"ffcc2dcd",
			2931 => x"00007c20",
			2932 => x"0c001710",
			2933 => x"00004608",
			2934 => x"0b001204",
			2935 => x"ffda2e59",
			2936 => x"00732e59",
			2937 => x"0f004604",
			2938 => x"ff772e59",
			2939 => x"00022e59",
			2940 => x"06002808",
			2941 => x"07002304",
			2942 => x"00292e59",
			2943 => x"ffb32e59",
			2944 => x"05001504",
			2945 => x"00062e59",
			2946 => x"00ab2e59",
			2947 => x"08001b20",
			2948 => x"06004e04",
			2949 => x"ffa62e59",
			2950 => x"0e005b10",
			2951 => x"05003d08",
			2952 => x"07002204",
			2953 => x"ffff2e59",
			2954 => x"00982e59",
			2955 => x"0000a804",
			2956 => x"ffc52e59",
			2957 => x"00142e59",
			2958 => x"0c001604",
			2959 => x"ffaf2e59",
			2960 => x"09001b04",
			2961 => x"002c2e59",
			2962 => x"ffec2e59",
			2963 => x"0b002f04",
			2964 => x"ff512e59",
			2965 => x"00262e59",
			2966 => x"05002b28",
			2967 => x"00007510",
			2968 => x"0b001204",
			2969 => x"ffe42eed",
			2970 => x"02002004",
			2971 => x"ffef2eed",
			2972 => x"09002a04",
			2973 => x"00662eed",
			2974 => x"00012eed",
			2975 => x"06004e04",
			2976 => x"ffac2eed",
			2977 => x"09001704",
			2978 => x"ffe52eed",
			2979 => x"0f007a0c",
			2980 => x"08001b04",
			2981 => x"00692eed",
			2982 => x"0b001a04",
			2983 => x"ffe22eed",
			2984 => x"000f2eed",
			2985 => x"ffe72eed",
			2986 => x"0c001b14",
			2987 => x"08001608",
			2988 => x"03002d04",
			2989 => x"00112eed",
			2990 => x"fffb2eed",
			2991 => x"0f004304",
			2992 => x"00032eed",
			2993 => x"0b001904",
			2994 => x"ffa22eed",
			2995 => x"ffff2eed",
			2996 => x"0d001608",
			2997 => x"04003904",
			2998 => x"00482eed",
			2999 => x"fff52eed",
			3000 => x"04001f04",
			3001 => x"00102eed",
			3002 => x"ffcb2eed",
			3003 => x"02009a30",
			3004 => x"0c00181c",
			3005 => x"0d000f04",
			3006 => x"003d2f59",
			3007 => x"0e002c08",
			3008 => x"0b001304",
			3009 => x"ffe92f59",
			3010 => x"003e2f59",
			3011 => x"05002304",
			3012 => x"ff7f2f59",
			3013 => x"05002b04",
			3014 => x"00442f59",
			3015 => x"0f005a04",
			3016 => x"ffaf2f59",
			3017 => x"00042f59",
			3018 => x"04003110",
			3019 => x"00002f04",
			3020 => x"ffdd2f59",
			3021 => x"0a001608",
			3022 => x"0a001004",
			3023 => x"00072f59",
			3024 => x"fffb2f59",
			3025 => x"007d2f59",
			3026 => x"ffdf2f59",
			3027 => x"08001604",
			3028 => x"fff92f59",
			3029 => x"ff892f59",
			3030 => x"0700252c",
			3031 => x"0f003210",
			3032 => x"0c001408",
			3033 => x"0d001004",
			3034 => x"d9f72fed",
			3035 => x"d8d72fed",
			3036 => x"0c001604",
			3037 => x"e7b02fed",
			3038 => x"eabb2fed",
			3039 => x"01000a14",
			3040 => x"0c001810",
			3041 => x"0a002a0c",
			3042 => x"0f005a08",
			3043 => x"0a001b04",
			3044 => x"d8d72fed",
			3045 => x"ddac2fed",
			3046 => x"e4b82fed",
			3047 => x"d8d22fed",
			3048 => x"e5662fed",
			3049 => x"02006b04",
			3050 => x"db862fed",
			3051 => x"d8cf2fed",
			3052 => x"0200a218",
			3053 => x"00002f04",
			3054 => x"d8cc2fed",
			3055 => x"00007c04",
			3056 => x"e8ae2fed",
			3057 => x"0c001b08",
			3058 => x"08001904",
			3059 => x"dec92fed",
			3060 => x"d8cf2fed",
			3061 => x"0a003704",
			3062 => x"e14b2fed",
			3063 => x"db132fed",
			3064 => x"05001c04",
			3065 => x"d9e62fed",
			3066 => x"d8cb2fed",
			3067 => x"01000a34",
			3068 => x"0c001510",
			3069 => x"0d000f08",
			3070 => x"0b001004",
			3071 => x"ffe23089",
			3072 => x"00493089",
			3073 => x"08001604",
			3074 => x"00083089",
			3075 => x"ffa13089",
			3076 => x"04003318",
			3077 => x"0f007914",
			3078 => x"0a00180c",
			3079 => x"00006b08",
			3080 => x"00002504",
			3081 => x"fff73089",
			3082 => x"00183089",
			3083 => x"ffe43089",
			3084 => x"08001d04",
			3085 => x"00743089",
			3086 => x"fff83089",
			3087 => x"ffea3089",
			3088 => x"0c001b04",
			3089 => x"ffce3089",
			3090 => x"0c001c04",
			3091 => x"00143089",
			3092 => x"fffa3089",
			3093 => x"09003014",
			3094 => x"08001804",
			3095 => x"000f3089",
			3096 => x"05000d04",
			3097 => x"00053089",
			3098 => x"05003f04",
			3099 => x"ff953089",
			3100 => x"05004004",
			3101 => x"00193089",
			3102 => x"ffe23089",
			3103 => x"04001b04",
			3104 => x"00293089",
			3105 => x"fff33089",
			3106 => x"05001508",
			3107 => x"0f001b04",
			3108 => x"fff130f5",
			3109 => x"003b30f5",
			3110 => x"0c001608",
			3111 => x"00004804",
			3112 => x"000030f5",
			3113 => x"ffb230f5",
			3114 => x"07002208",
			3115 => x"0a001e04",
			3116 => x"fffd30f5",
			3117 => x"004730f5",
			3118 => x"06004708",
			3119 => x"04001204",
			3120 => x"000330f5",
			3121 => x"ffc230f5",
			3122 => x"0d00130c",
			3123 => x"04002d08",
			3124 => x"0000be04",
			3125 => x"005130f5",
			3126 => x"fffc30f5",
			3127 => x"ffec30f5",
			3128 => x"02008b04",
			3129 => x"002730f5",
			3130 => x"09002404",
			3131 => x"ffb930f5",
			3132 => x"000930f5",
			3133 => x"04001c28",
			3134 => x"03001c20",
			3135 => x"04000c0c",
			3136 => x"00002104",
			3137 => x"fff63189",
			3138 => x"04000504",
			3139 => x"ffff3189",
			3140 => x"00313189",
			3141 => x"05001b0c",
			3142 => x"08002308",
			3143 => x"08001f04",
			3144 => x"ffbc3189",
			3145 => x"00003189",
			3146 => x"00043189",
			3147 => x"05001c04",
			3148 => x"00113189",
			3149 => x"ffee3189",
			3150 => x"06007104",
			3151 => x"005a3189",
			3152 => x"fff13189",
			3153 => x"01000b20",
			3154 => x"06004104",
			3155 => x"00323189",
			3156 => x"0a003610",
			3157 => x"06006108",
			3158 => x"09001c04",
			3159 => x"00033189",
			3160 => x"ffb03189",
			3161 => x"08001904",
			3162 => x"00163189",
			3163 => x"fff93189",
			3164 => x"05004608",
			3165 => x"0b001704",
			3166 => x"fff83189",
			3167 => x"00403189",
			3168 => x"ffe63189",
			3169 => x"ffc03189",
			3170 => x"02009a34",
			3171 => x"0c001104",
			3172 => x"ffc8320d",
			3173 => x"07002218",
			3174 => x"05002b10",
			3175 => x"01000c08",
			3176 => x"04000704",
			3177 => x"0002320d",
			3178 => x"0092320d",
			3179 => x"0c001904",
			3180 => x"ffe7320d",
			3181 => x"000c320d",
			3182 => x"04002604",
			3183 => x"ffcc320d",
			3184 => x"0022320d",
			3185 => x"0c001b10",
			3186 => x"0200940c",
			3187 => x"0b001908",
			3188 => x"00007204",
			3189 => x"0002320d",
			3190 => x"ff88320d",
			3191 => x"0009320d",
			3192 => x"0033320d",
			3193 => x"06002804",
			3194 => x"ffcd320d",
			3195 => x"006e320d",
			3196 => x"05001c04",
			3197 => x"0021320d",
			3198 => x"09002404",
			3199 => x"ff8f320d",
			3200 => x"09002504",
			3201 => x"0012320d",
			3202 => x"ffec320d",
			3203 => x"0700252c",
			3204 => x"02006b18",
			3205 => x"0b001204",
			3206 => x"fe5c32a9",
			3207 => x"0e003810",
			3208 => x"0100100c",
			3209 => x"0a000a04",
			3210 => x"039a32a9",
			3211 => x"0b001504",
			3212 => x"015432a9",
			3213 => x"02b932a9",
			3214 => x"018032a9",
			3215 => x"ffe932a9",
			3216 => x"08001b10",
			3217 => x"0200a50c",
			3218 => x"06004e04",
			3219 => x"ff9132a9",
			3220 => x"03002404",
			3221 => x"03a332a9",
			3222 => x"005a32a9",
			3223 => x"fe5432a9",
			3224 => x"fe5232a9",
			3225 => x"0200a21c",
			3226 => x"00002f04",
			3227 => x"fe5532a9",
			3228 => x"0c001b0c",
			3229 => x"03002f08",
			3230 => x"0c001604",
			3231 => x"fe4a32a9",
			3232 => x"01d432a9",
			3233 => x"fe4232a9",
			3234 => x"0a003b08",
			3235 => x"0a002704",
			3236 => x"015a32a9",
			3237 => x"03b032a9",
			3238 => x"ff0e32a9",
			3239 => x"05001c04",
			3240 => x"fffb32a9",
			3241 => x"fe5332a9",
			3242 => x"05002b38",
			3243 => x"03001c20",
			3244 => x"05001510",
			3245 => x"0f001b04",
			3246 => x"ffe23365",
			3247 => x"00005204",
			3248 => x"006d3365",
			3249 => x"06003f04",
			3250 => x"ffd03365",
			3251 => x"00353365",
			3252 => x"0a001e0c",
			3253 => x"08002404",
			3254 => x"ff6e3365",
			3255 => x"08002604",
			3256 => x"00043365",
			3257 => x"fffa3365",
			3258 => x"00013365",
			3259 => x"0f007a14",
			3260 => x"01000a04",
			3261 => x"00b63365",
			3262 => x"0d001908",
			3263 => x"02005c04",
			3264 => x"000d3365",
			3265 => x"ffc03365",
			3266 => x"00003d04",
			3267 => x"fff93365",
			3268 => x"003c3365",
			3269 => x"ffb83365",
			3270 => x"0c001b18",
			3271 => x"0f004304",
			3272 => x"00123365",
			3273 => x"08001608",
			3274 => x"01000504",
			3275 => x"fffc3365",
			3276 => x"00223365",
			3277 => x"0d001104",
			3278 => x"00043365",
			3279 => x"0b001904",
			3280 => x"ff233365",
			3281 => x"fff33365",
			3282 => x"08001d08",
			3283 => x"05004a04",
			3284 => x"00a23365",
			3285 => x"fff13365",
			3286 => x"04001f04",
			3287 => x"001a3365",
			3288 => x"ff923365",
			3289 => x"0f007830",
			3290 => x"05004128",
			3291 => x"08001c14",
			3292 => x"0c001104",
			3293 => x"ffd533c9",
			3294 => x"08001504",
			3295 => x"fff033c9",
			3296 => x"00002104",
			3297 => x"fff333c9",
			3298 => x"01000b04",
			3299 => x"008633c9",
			3300 => x"fff833c9",
			3301 => x"04001c10",
			3302 => x"0c001704",
			3303 => x"ffe633c9",
			3304 => x"00003304",
			3305 => x"fff133c9",
			3306 => x"00009404",
			3307 => x"004b33c9",
			3308 => x"fff333c9",
			3309 => x"ffbc33c9",
			3310 => x"0b001a04",
			3311 => x"ffac33c9",
			3312 => x"002a33c9",
			3313 => x"ffc433c9",
			3314 => x"0700252c",
			3315 => x"02006b18",
			3316 => x"0b001204",
			3317 => x"fe5f3465",
			3318 => x"01000404",
			3319 => x"03843465",
			3320 => x"0c001504",
			3321 => x"ff6d3465",
			3322 => x"0b001504",
			3323 => x"014d3465",
			3324 => x"0f003104",
			3325 => x"024e3465",
			3326 => x"03313465",
			3327 => x"04001304",
			3328 => x"fe4f3465",
			3329 => x"05002608",
			3330 => x"0f005904",
			3331 => x"00933465",
			3332 => x"02823465",
			3333 => x"00008804",
			3334 => x"015a3465",
			3335 => x"fe513465",
			3336 => x"0200a21c",
			3337 => x"00002f04",
			3338 => x"fe583465",
			3339 => x"03003914",
			3340 => x"0c001b0c",
			3341 => x"0d001304",
			3342 => x"01553465",
			3343 => x"06005504",
			3344 => x"ffd13465",
			3345 => x"fe463465",
			3346 => x"0a002c04",
			3347 => x"010b3465",
			3348 => x"03ae3465",
			3349 => x"fe173465",
			3350 => x"05001c04",
			3351 => x"ffe43465",
			3352 => x"fe553465",
			3353 => x"01000a30",
			3354 => x"0b001208",
			3355 => x"00009b04",
			3356 => x"ffd83501",
			3357 => x"000f3501",
			3358 => x"06006f24",
			3359 => x"0500411c",
			3360 => x"0a00180c",
			3361 => x"00005208",
			3362 => x"00002104",
			3363 => x"fff53501",
			3364 => x"00323501",
			3365 => x"ffcf3501",
			3366 => x"08001c08",
			3367 => x"09001e04",
			3368 => x"00673501",
			3369 => x"000a3501",
			3370 => x"09001e04",
			3371 => x"fff63501",
			3372 => x"00023501",
			3373 => x"0c001b04",
			3374 => x"ffd73501",
			3375 => x"001a3501",
			3376 => x"ffea3501",
			3377 => x"04001c14",
			3378 => x"0b001b0c",
			3379 => x"0e002308",
			3380 => x"08001c04",
			3381 => x"00083501",
			3382 => x"ffff3501",
			3383 => x"ffeb3501",
			3384 => x"00003704",
			3385 => x"fff93501",
			3386 => x"002c3501",
			3387 => x"08001b08",
			3388 => x"08001904",
			3389 => x"000b3501",
			3390 => x"00003501",
			3391 => x"ffb53501",
			3392 => x"0e005244",
			3393 => x"0c00181c",
			3394 => x"05002b14",
			3395 => x"0c001304",
			3396 => x"ff2635cd",
			3397 => x"0f004b0c",
			3398 => x"02006b08",
			3399 => x"0a001404",
			3400 => x"fff335cd",
			3401 => x"00c735cd",
			3402 => x"ff1a35cd",
			3403 => x"00db35cd",
			3404 => x"0f005a04",
			3405 => x"fef835cd",
			3406 => x"fffb35cd",
			3407 => x"08001d18",
			3408 => x"04001810",
			3409 => x"07002204",
			3410 => x"008435cd",
			3411 => x"07002804",
			3412 => x"ff6035cd",
			3413 => x"0a000f04",
			3414 => x"001035cd",
			3415 => x"fff735cd",
			3416 => x"02009704",
			3417 => x"011635cd",
			3418 => x"fffd35cd",
			3419 => x"04001c0c",
			3420 => x"00007c08",
			3421 => x"00003504",
			3422 => x"ffb535cd",
			3423 => x"00db35cd",
			3424 => x"ff9e35cd",
			3425 => x"ff4535cd",
			3426 => x"0a002810",
			3427 => x"0c001608",
			3428 => x"0d001004",
			3429 => x"007235cd",
			3430 => x"fefa35cd",
			3431 => x"0f007d04",
			3432 => x"00d935cd",
			3433 => x"ffcd35cd",
			3434 => x"08001608",
			3435 => x"05003204",
			3436 => x"ffe135cd",
			3437 => x"004d35cd",
			3438 => x"0c001b04",
			3439 => x"feb435cd",
			3440 => x"0000ad04",
			3441 => x"005e35cd",
			3442 => x"ff4035cd",
			3443 => x"0e005b40",
			3444 => x"0c001b24",
			3445 => x"03002e20",
			3446 => x"0800180c",
			3447 => x"06004e08",
			3448 => x"02004604",
			3449 => x"00bc3661",
			3450 => x"ff933661",
			3451 => x"012a3661",
			3452 => x"0c001504",
			3453 => x"fef63661",
			3454 => x"06003808",
			3455 => x"0a001104",
			3456 => x"ffde3661",
			3457 => x"00f03661",
			3458 => x"09001d04",
			3459 => x"00773661",
			3460 => x"ff5b3661",
			3461 => x"fede3661",
			3462 => x"06002808",
			3463 => x"07002304",
			3464 => x"005a3661",
			3465 => x"ff2d3661",
			3466 => x"0a002a08",
			3467 => x"00008304",
			3468 => x"00d73661",
			3469 => x"ff363661",
			3470 => x"03003908",
			3471 => x"0000ad04",
			3472 => x"01603661",
			3473 => x"ffe23661",
			3474 => x"ff8f3661",
			3475 => x"0a002004",
			3476 => x"00063661",
			3477 => x"0c002d04",
			3478 => x"feaa3661",
			3479 => x"00323661",
			3480 => x"07002528",
			3481 => x"0c001304",
			3482 => x"ff8c3725",
			3483 => x"05002d1c",
			3484 => x"0a00140c",
			3485 => x"00005208",
			3486 => x"07001b04",
			3487 => x"004c3725",
			3488 => x"00003725",
			3489 => x"ffad3725",
			3490 => x"09001e08",
			3491 => x"01000b04",
			3492 => x"00c93725",
			3493 => x"ffe73725",
			3494 => x"00006b04",
			3495 => x"00473725",
			3496 => x"ffcf3725",
			3497 => x"0b001504",
			3498 => x"ffa93725",
			3499 => x"00293725",
			3500 => x"0c001b1c",
			3501 => x"08001608",
			3502 => x"05003004",
			3503 => x"fff23725",
			3504 => x"002c3725",
			3505 => x"0a002410",
			3506 => x"03001c08",
			3507 => x"03000e04",
			3508 => x"00023725",
			3509 => x"ffb63725",
			3510 => x"08001904",
			3511 => x"00463725",
			3512 => x"fffa3725",
			3513 => x"ff443725",
			3514 => x"01000a10",
			3515 => x"03002708",
			3516 => x"05001004",
			3517 => x"00003725",
			3518 => x"ffe13725",
			3519 => x"03003e04",
			3520 => x"00943725",
			3521 => x"fff13725",
			3522 => x"09003308",
			3523 => x"07002704",
			3524 => x"00083725",
			3525 => x"ff963725",
			3526 => x"03003404",
			3527 => x"001d3725",
			3528 => x"fff83725",
			3529 => x"0c001304",
			3530 => x"ffbc37a9",
			3531 => x"08001b20",
			3532 => x"05004118",
			3533 => x"0f007914",
			3534 => x"0a00140c",
			3535 => x"00005208",
			3536 => x"00002504",
			3537 => x"fffb37a9",
			3538 => x"002137a9",
			3539 => x"ffd637a9",
			3540 => x"05001704",
			3541 => x"000037a9",
			3542 => x"006a37a9",
			3543 => x"ffe737a9",
			3544 => x"0b001904",
			3545 => x"ffcd37a9",
			3546 => x"001037a9",
			3547 => x"0b001910",
			3548 => x"0e00380c",
			3549 => x"07001d04",
			3550 => x"fff137a9",
			3551 => x"00003d04",
			3552 => x"fff737a9",
			3553 => x"001a37a9",
			3554 => x"ffa037a9",
			3555 => x"0200990c",
			3556 => x"06002808",
			3557 => x"07002304",
			3558 => x"000d37a9",
			3559 => x"ffd737a9",
			3560 => x"004d37a9",
			3561 => x"ffd837a9",
			3562 => x"07002534",
			3563 => x"02005818",
			3564 => x"0b001204",
			3565 => x"fe6a3845",
			3566 => x"05002410",
			3567 => x"08001804",
			3568 => x"02e13845",
			3569 => x"06001f04",
			3570 => x"015d3845",
			3571 => x"07001a04",
			3572 => x"01bb3845",
			3573 => x"021d3845",
			3574 => x"00de3845",
			3575 => x"01000b14",
			3576 => x"0200a510",
			3577 => x"0a001604",
			3578 => x"fe5b3845",
			3579 => x"04002b08",
			3580 => x"0c001704",
			3581 => x"015b3845",
			3582 => x"02b23845",
			3583 => x"fe6d3845",
			3584 => x"fe613845",
			3585 => x"0b001804",
			3586 => x"fe4f3845",
			3587 => x"00713845",
			3588 => x"0200ae18",
			3589 => x"00002f04",
			3590 => x"fe5e3845",
			3591 => x"04003310",
			3592 => x"0c001604",
			3593 => x"fe4c3845",
			3594 => x"0d001404",
			3595 => x"02c23845",
			3596 => x"00009404",
			3597 => x"01613845",
			3598 => x"ff0a3845",
			3599 => x"fe533845",
			3600 => x"fe5a3845",
			3601 => x"07002530",
			3602 => x"0c001304",
			3603 => x"ff863919",
			3604 => x"01000a18",
			3605 => x"0a001408",
			3606 => x"00005204",
			3607 => x"00313919",
			3608 => x"ffb33919",
			3609 => x"05003c0c",
			3610 => x"08001c08",
			3611 => x"0200a504",
			3612 => x"00ca3919",
			3613 => x"fff83919",
			3614 => x"fff93919",
			3615 => x"ffea3919",
			3616 => x"0b001708",
			3617 => x"05002704",
			3618 => x"00073919",
			3619 => x"ff9b3919",
			3620 => x"08002208",
			3621 => x"00007c04",
			3622 => x"005f3919",
			3623 => x"fff33919",
			3624 => x"ffdd3919",
			3625 => x"0c001b1c",
			3626 => x"08001608",
			3627 => x"05003004",
			3628 => x"fff13919",
			3629 => x"002e3919",
			3630 => x"0a002410",
			3631 => x"03001c08",
			3632 => x"03000e04",
			3633 => x"00023919",
			3634 => x"ffb33919",
			3635 => x"08001904",
			3636 => x"00483919",
			3637 => x"fffa3919",
			3638 => x"ff3a3919",
			3639 => x"01000a10",
			3640 => x"03002708",
			3641 => x"07002a04",
			3642 => x"ffdf3919",
			3643 => x"00013919",
			3644 => x"03003e04",
			3645 => x"00993919",
			3646 => x"fff03919",
			3647 => x"09003308",
			3648 => x"07002704",
			3649 => x"00083919",
			3650 => x"ff923919",
			3651 => x"03003404",
			3652 => x"001e3919",
			3653 => x"fff83919",
			3654 => x"0e00503c",
			3655 => x"08001d24",
			3656 => x"0b001204",
			3657 => x"ff4d39dd",
			3658 => x"02009718",
			3659 => x"0a00190c",
			3660 => x"00004d08",
			3661 => x"00002104",
			3662 => x"ffba39dd",
			3663 => x"00e439dd",
			3664 => x"ff4a39dd",
			3665 => x"01000b08",
			3666 => x"04003104",
			3667 => x"010639dd",
			3668 => x"002439dd",
			3669 => x"fffe39dd",
			3670 => x"0e004b04",
			3671 => x"ff7339dd",
			3672 => x"005a39dd",
			3673 => x"04001c14",
			3674 => x"0a002110",
			3675 => x"0500160c",
			3676 => x"00006e08",
			3677 => x"00003504",
			3678 => x"ffeb39dd",
			3679 => x"005039dd",
			3680 => x"ffd039dd",
			3681 => x"ff8139dd",
			3682 => x"008339dd",
			3683 => x"ff0c39dd",
			3684 => x"0a002810",
			3685 => x"0c001608",
			3686 => x"0d000f04",
			3687 => x"006739dd",
			3688 => x"ff2639dd",
			3689 => x"0f007d04",
			3690 => x"00ec39dd",
			3691 => x"ffd339dd",
			3692 => x"09003a14",
			3693 => x"08001608",
			3694 => x"0d001104",
			3695 => x"002039dd",
			3696 => x"ffde39dd",
			3697 => x"0c001b04",
			3698 => x"febc39dd",
			3699 => x"0c001c04",
			3700 => x"fffe39dd",
			3701 => x"ff7039dd",
			3702 => x"004539dd",
			3703 => x"01000620",
			3704 => x"03001c0c",
			3705 => x"05001508",
			3706 => x"0c001704",
			3707 => x"00883ab1",
			3708 => x"ffda3ab1",
			3709 => x"ff633ab1",
			3710 => x"0f004b04",
			3711 => x"fff83ab1",
			3712 => x"0e00610c",
			3713 => x"04003308",
			3714 => x"0200af04",
			3715 => x"00d53ab1",
			3716 => x"fff63ab1",
			3717 => x"ffd43ab1",
			3718 => x"ffc73ab1",
			3719 => x"0e003d24",
			3720 => x"0b001508",
			3721 => x"04001104",
			3722 => x"000b3ab1",
			3723 => x"ff883ab1",
			3724 => x"0b00200c",
			3725 => x"02007408",
			3726 => x"00002804",
			3727 => x"ffea3ab1",
			3728 => x"00d73ab1",
			3729 => x"ffe63ab1",
			3730 => x"08002304",
			3731 => x"00093ab1",
			3732 => x"03001a08",
			3733 => x"03001804",
			3734 => x"ffff3ab1",
			3735 => x"00033ab1",
			3736 => x"ffb23ab1",
			3737 => x"0c001b10",
			3738 => x"08001604",
			3739 => x"001d3ab1",
			3740 => x"05002508",
			3741 => x"05002404",
			3742 => x"ffc73ab1",
			3743 => x"00333ab1",
			3744 => x"feef3ab1",
			3745 => x"0a003b14",
			3746 => x"0a002f08",
			3747 => x"07003a04",
			3748 => x"ffbe3ab1",
			3749 => x"001e3ab1",
			3750 => x"07003404",
			3751 => x"007f3ab1",
			3752 => x"07004004",
			3753 => x"ffe53ab1",
			3754 => x"001b3ab1",
			3755 => x"ffa53ab1",
			3756 => x"0200ae40",
			3757 => x"0c001614",
			3758 => x"00004608",
			3759 => x"0b001204",
			3760 => x"ffcd3b35",
			3761 => x"009b3b35",
			3762 => x"08001604",
			3763 => x"00293b35",
			3764 => x"00009f04",
			3765 => x"ff123b35",
			3766 => x"fffe3b35",
			3767 => x"05004628",
			3768 => x"0a001b10",
			3769 => x"00006b08",
			3770 => x"00002804",
			3771 => x"ffba3b35",
			3772 => x"00673b35",
			3773 => x"01000e04",
			3774 => x"ff8b3b35",
			3775 => x"fffd3b35",
			3776 => x"01000b0c",
			3777 => x"08001d08",
			3778 => x"05002104",
			3779 => x"00273b35",
			3780 => x"00cf3b35",
			3781 => x"ffd83b35",
			3782 => x"05003108",
			3783 => x"00008804",
			3784 => x"00823b35",
			3785 => x"fffd3b35",
			3786 => x"ff853b35",
			3787 => x"ff6e3b35",
			3788 => x"ff2f3b35",
			3789 => x"0e006144",
			3790 => x"04001418",
			3791 => x"0c001104",
			3792 => x"fec73bc1",
			3793 => x"02002004",
			3794 => x"ff0a3bc1",
			3795 => x"02005004",
			3796 => x"016d3bc1",
			3797 => x"03001a08",
			3798 => x"06004a04",
			3799 => x"fec13bc1",
			3800 => x"00533bc1",
			3801 => x"01503bc1",
			3802 => x"08001d1c",
			3803 => x"0c001b14",
			3804 => x"0e003908",
			3805 => x"0b001504",
			3806 => x"ff693bc1",
			3807 => x"017c3bc1",
			3808 => x"01000304",
			3809 => x"00fa3bc1",
			3810 => x"0f006704",
			3811 => x"fec53bc1",
			3812 => x"00293bc1",
			3813 => x"0c001c04",
			3814 => x"016f3bc1",
			3815 => x"fede3bc1",
			3816 => x"04001c0c",
			3817 => x"0a002708",
			3818 => x"01000c04",
			3819 => x"ffe33bc1",
			3820 => x"ff053bc1",
			3821 => x"00f43bc1",
			3822 => x"fe6d3bc1",
			3823 => x"fe7a3bc1",
			3824 => x"0200ae34",
			3825 => x"0500412c",
			3826 => x"05003a28",
			3827 => x"01000a14",
			3828 => x"0b001204",
			3829 => x"fede3c2d",
			3830 => x"02006b08",
			3831 => x"00002104",
			3832 => x"ff713c2d",
			3833 => x"010f3c2d",
			3834 => x"0f005804",
			3835 => x"ff373c2d",
			3836 => x"009b3c2d",
			3837 => x"04001c0c",
			3838 => x"0a002708",
			3839 => x"05001504",
			3840 => x"00593c2d",
			3841 => x"ff443c2d",
			3842 => x"01093c2d",
			3843 => x"04001e04",
			3844 => x"ffd73c2d",
			3845 => x"feb93c2d",
			3846 => x"010c3c2d",
			3847 => x"09002204",
			3848 => x"feb03c2d",
			3849 => x"00673c2d",
			3850 => x"fe8f3c2d",
			3851 => x"0e005b50",
			3852 => x"0b001930",
			3853 => x"09001f28",
			3854 => x"0c001818",
			3855 => x"05002b10",
			3856 => x"0c001308",
			3857 => x"06002304",
			3858 => x"00303cd9",
			3859 => x"ff3e3cd9",
			3860 => x"08001c04",
			3861 => x"007b3cd9",
			3862 => x"ff973cd9",
			3863 => x"01000704",
			3864 => x"fff43cd9",
			3865 => x"ff193cd9",
			3866 => x"0000a60c",
			3867 => x"03001a08",
			3868 => x"00007804",
			3869 => x"00283cd9",
			3870 => x"ffc73cd9",
			3871 => x"00e23cd9",
			3872 => x"ffda3cd9",
			3873 => x"0c001b04",
			3874 => x"ff133cd9",
			3875 => x"ffe53cd9",
			3876 => x"01000a0c",
			3877 => x"0a001908",
			3878 => x"05001004",
			3879 => x"00063cd9",
			3880 => x"fff33cd9",
			3881 => x"00ef3cd9",
			3882 => x"0000810c",
			3883 => x"06002808",
			3884 => x"07002304",
			3885 => x"00323cd9",
			3886 => x"ff863cd9",
			3887 => x"00a53cd9",
			3888 => x"07002d04",
			3889 => x"ff713cd9",
			3890 => x"000a3cd9",
			3891 => x"08003504",
			3892 => x"fee13cd9",
			3893 => x"00213cd9",
			3894 => x"0f007838",
			3895 => x"0a003734",
			3896 => x"08001c18",
			3897 => x"0a003614",
			3898 => x"05003c10",
			3899 => x"00009b08",
			3900 => x"07002504",
			3901 => x"00613d4d",
			3902 => x"fee93d4d",
			3903 => x"06005604",
			3904 => x"ff4d3d4d",
			3905 => x"01543d4d",
			3906 => x"ff043d4d",
			3907 => x"01293d4d",
			3908 => x"0b00190c",
			3909 => x"06002408",
			3910 => x"0e001504",
			3911 => x"fff83d4d",
			3912 => x"00123d4d",
			3913 => x"feee3d4d",
			3914 => x"06002808",
			3915 => x"07002304",
			3916 => x"007c3d4d",
			3917 => x"ff183d4d",
			3918 => x"00009404",
			3919 => x"010f3d4d",
			3920 => x"ff553d4d",
			3921 => x"fedc3d4d",
			3922 => x"feae3d4d",
			3923 => x"0200a550",
			3924 => x"0c001b38",
			3925 => x"08001c28",
			3926 => x"02006b10",
			3927 => x"0b001204",
			3928 => x"ff8e3df1",
			3929 => x"01000a08",
			3930 => x"03001304",
			3931 => x"002c3df1",
			3932 => x"01113df1",
			3933 => x"fff83df1",
			3934 => x"00009b10",
			3935 => x"04001408",
			3936 => x"01000704",
			3937 => x"00343df1",
			3938 => x"ffdc3df1",
			3939 => x"0a003104",
			3940 => x"ff0b3df1",
			3941 => x"fffb3df1",
			3942 => x"0d001304",
			3943 => x"00cb3df1",
			3944 => x"ffae3df1",
			3945 => x"06002408",
			3946 => x"00002f04",
			3947 => x"fffb3df1",
			3948 => x"001d3df1",
			3949 => x"04001204",
			3950 => x"fff13df1",
			3951 => x"ff1e3df1",
			3952 => x"06002808",
			3953 => x"07002304",
			3954 => x"00323df1",
			3955 => x"ff783df1",
			3956 => x"0a002a08",
			3957 => x"00008b04",
			3958 => x"00a53df1",
			3959 => x"ff853df1",
			3960 => x"00007804",
			3961 => x"001b3df1",
			3962 => x"01043df1",
			3963 => x"feea3df1",
			3964 => x"0200ae38",
			3965 => x"02002004",
			3966 => x"fe733e65",
			3967 => x"04001c18",
			3968 => x"0c001104",
			3969 => x"fe4a3e65",
			3970 => x"06007010",
			3971 => x"02005008",
			3972 => x"09002a04",
			3973 => x"019d3e65",
			3974 => x"fedf3e65",
			3975 => x"0a001604",
			3976 => x"fe713e65",
			3977 => x"01213e65",
			3978 => x"fe903e65",
			3979 => x"08001d14",
			3980 => x"0c001a0c",
			3981 => x"05004108",
			3982 => x"0c001604",
			3983 => x"ff223e65",
			3984 => x"01053e65",
			3985 => x"fe653e65",
			3986 => x"05004704",
			3987 => x"01b03e65",
			3988 => x"fee13e65",
			3989 => x"09002404",
			3990 => x"fe683e65",
			3991 => x"fd833e65",
			3992 => x"fe683e65",
			3993 => x"0e006140",
			3994 => x"08001b20",
			3995 => x"0500411c",
			3996 => x"0c001104",
			3997 => x"feef3ee9",
			3998 => x"0f004b10",
			3999 => x"02004608",
			4000 => x"00002104",
			4001 => x"ffd13ee9",
			4002 => x"01533ee9",
			4003 => x"0c001704",
			4004 => x"ff463ee9",
			4005 => x"00f13ee9",
			4006 => x"0b001304",
			4007 => x"00783ee9",
			4008 => x"01683ee9",
			4009 => x"fecd3ee9",
			4010 => x"0b001504",
			4011 => x"feb53ee9",
			4012 => x"07002308",
			4013 => x"0e003704",
			4014 => x"013e3ee9",
			4015 => x"fff73ee9",
			4016 => x"0c001b08",
			4017 => x"0a000d04",
			4018 => x"ffe23ee9",
			4019 => x"fe9e3ee9",
			4020 => x"06002904",
			4021 => x"fec33ee9",
			4022 => x"02009904",
			4023 => x"00df3ee9",
			4024 => x"ff103ee9",
			4025 => x"fe8c3ee9",
			4026 => x"0e00613c",
			4027 => x"05004638",
			4028 => x"01000a18",
			4029 => x"02005008",
			4030 => x"00002104",
			4031 => x"fec83f65",
			4032 => x"019c3f65",
			4033 => x"05001804",
			4034 => x"feef3f65",
			4035 => x"04001404",
			4036 => x"01a23f65",
			4037 => x"0b001904",
			4038 => x"00123f65",
			4039 => x"01a83f65",
			4040 => x"0c001808",
			4041 => x"04001204",
			4042 => x"ffdc3f65",
			4043 => x"fe783f65",
			4044 => x"07002608",
			4045 => x"00007c04",
			4046 => x"01843f65",
			4047 => x"fee43f65",
			4048 => x"0e005008",
			4049 => x"0a002804",
			4050 => x"fe8c3f65",
			4051 => x"ffa63f65",
			4052 => x"05003404",
			4053 => x"015b3f65",
			4054 => x"fef03f65",
			4055 => x"fe8a3f65",
			4056 => x"fe6d3f65",
			4057 => x"0200a548",
			4058 => x"0700252c",
			4059 => x"0c001820",
			4060 => x"01000a18",
			4061 => x"02006b0c",
			4062 => x"0b001204",
			4063 => x"fea33ff9",
			4064 => x"00004804",
			4065 => x"01da3ff9",
			4066 => x"01193ff9",
			4067 => x"06004e04",
			4068 => x"fe453ff9",
			4069 => x"05004104",
			4070 => x"00f83ff9",
			4071 => x"ff023ff9",
			4072 => x"06002704",
			4073 => x"ffc13ff9",
			4074 => x"fe643ff9",
			4075 => x"02007408",
			4076 => x"0a001204",
			4077 => x"00a63ff9",
			4078 => x"01b83ff9",
			4079 => x"fffb3ff9",
			4080 => x"00002f04",
			4081 => x"fe793ff9",
			4082 => x"04003214",
			4083 => x"09001b04",
			4084 => x"fe6e3ff9",
			4085 => x"0f005208",
			4086 => x"00008b04",
			4087 => x"00ad3ff9",
			4088 => x"fe6a3ff9",
			4089 => x"0b001904",
			4090 => x"00543ff9",
			4091 => x"01a63ff9",
			4092 => x"fe6e3ff9",
			4093 => x"fe673ff9",
			4094 => x"0200ae40",
			4095 => x"02002004",
			4096 => x"fe61407d",
			4097 => x"05002b20",
			4098 => x"00007510",
			4099 => x"0b001204",
			4100 => x"fe7c407d",
			4101 => x"01000404",
			4102 => x"0233407d",
			4103 => x"0b001504",
			4104 => x"0010407d",
			4105 => x"01a8407d",
			4106 => x"0f005404",
			4107 => x"fe41407d",
			4108 => x"06007008",
			4109 => x"08001b04",
			4110 => x"01c3407d",
			4111 => x"002d407d",
			4112 => x"fe76407d",
			4113 => x"08001d10",
			4114 => x"0c001a08",
			4115 => x"05004104",
			4116 => x"0020407d",
			4117 => x"fe57407d",
			4118 => x"04003804",
			4119 => x"0246407d",
			4120 => x"fea7407d",
			4121 => x"07002504",
			4122 => x"fd85407d",
			4123 => x"07002c04",
			4124 => x"fe5a407d",
			4125 => x"fefa407d",
			4126 => x"fe63407d",
			4127 => x"0200ae48",
			4128 => x"0c001b30",
			4129 => x"03002e2c",
			4130 => x"0800180c",
			4131 => x"06004e08",
			4132 => x"02004604",
			4133 => x"00cc4111",
			4134 => x"ff844111",
			4135 => x"00ec4111",
			4136 => x"06003810",
			4137 => x"0b001508",
			4138 => x"0e002404",
			4139 => x"00304111",
			4140 => x"ff3c4111",
			4141 => x"00002804",
			4142 => x"ffb54111",
			4143 => x"01044111",
			4144 => x"00009b08",
			4145 => x"07002304",
			4146 => x"fec04111",
			4147 => x"ffba4111",
			4148 => x"0e005404",
			4149 => x"00714111",
			4150 => x"ffa24111",
			4151 => x"fec94111",
			4152 => x"06002808",
			4153 => x"07002304",
			4154 => x"005e4111",
			4155 => x"ff224111",
			4156 => x"03003a0c",
			4157 => x"0a002a08",
			4158 => x"00008304",
			4159 => x"00e04111",
			4160 => x"ff2d4111",
			4161 => x"01624111",
			4162 => x"ff824111",
			4163 => x"feb24111",
			4164 => x"0e006148",
			4165 => x"08001d28",
			4166 => x"05004624",
			4167 => x"0a00361c",
			4168 => x"08001810",
			4169 => x"06003d08",
			4170 => x"06002604",
			4171 => x"00ae41a5",
			4172 => x"ff5f41a5",
			4173 => x"0200af04",
			4174 => x"010a41a5",
			4175 => x"ffe441a5",
			4176 => x"0c001504",
			4177 => x"ff1941a5",
			4178 => x"0e003804",
			4179 => x"00d941a5",
			4180 => x"ffde41a5",
			4181 => x"0b001704",
			4182 => x"ffbb41a5",
			4183 => x"014f41a5",
			4184 => x"ff3441a5",
			4185 => x"04001c1c",
			4186 => x"0b001b10",
			4187 => x"0600310c",
			4188 => x"02003608",
			4189 => x"0a000f04",
			4190 => x"000541a5",
			4191 => x"ffdd41a5",
			4192 => x"003541a5",
			4193 => x"ff7d41a5",
			4194 => x"00003704",
			4195 => x"ffb541a5",
			4196 => x"00009f04",
			4197 => x"00fb41a5",
			4198 => x"ffd741a5",
			4199 => x"fede41a5",
			4200 => x"fecb41a5",
			4201 => x"0e006150",
			4202 => x"0c001b30",
			4203 => x"0500402c",
			4204 => x"08001b1c",
			4205 => x"03001c0c",
			4206 => x"05001508",
			4207 => x"0c001704",
			4208 => x"009a4249",
			4209 => x"ffd64249",
			4210 => x"ff544249",
			4211 => x"0f005408",
			4212 => x"0e003904",
			4213 => x"00794249",
			4214 => x"ffb44249",
			4215 => x"0000b804",
			4216 => x"010a4249",
			4217 => x"fff14249",
			4218 => x"0e00410c",
			4219 => x"0c001604",
			4220 => x"ff664249",
			4221 => x"08001d04",
			4222 => x"00bf4249",
			4223 => x"ffef4249",
			4224 => x"ff0e4249",
			4225 => x"ff174249",
			4226 => x"01000a10",
			4227 => x"0a00270c",
			4228 => x"0c001c08",
			4229 => x"04000b04",
			4230 => x"ffff4249",
			4231 => x"00054249",
			4232 => x"ffe04249",
			4233 => x"00f34249",
			4234 => x"0000940c",
			4235 => x"06002808",
			4236 => x"07002304",
			4237 => x"00244249",
			4238 => x"ff954249",
			4239 => x"00a14249",
			4240 => x"ff784249",
			4241 => x"ff234249",
			4242 => x"0e006144",
			4243 => x"0a003740",
			4244 => x"08001810",
			4245 => x"0b001204",
			4246 => x"ffb242d7",
			4247 => x"09001a04",
			4248 => x"013342d7",
			4249 => x"03002304",
			4250 => x"ff8f42d7",
			4251 => x"00b642d7",
			4252 => x"0c001714",
			4253 => x"00009710",
			4254 => x"0e002c08",
			4255 => x"07001704",
			4256 => x"ff9542d7",
			4257 => x"008742d7",
			4258 => x"07002304",
			4259 => x"febd42d7",
			4260 => x"ffb342d7",
			4261 => x"008d42d7",
			4262 => x"00007c10",
			4263 => x"06002808",
			4264 => x"07002304",
			4265 => x"00c942d7",
			4266 => x"fef642d7",
			4267 => x"0a001b04",
			4268 => x"004d42d7",
			4269 => x"016442d7",
			4270 => x"0f005804",
			4271 => x"fecb42d7",
			4272 => x"0c001b04",
			4273 => x"ffc142d7",
			4274 => x"012542d7",
			4275 => x"fed942d7",
			4276 => x"fea742d7",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1469, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2865, initial_addr_3'length));
	end generate gen_rom_11;

	gen_rom_12: if SELECT_ROM = 12 generate
		bank <= (
			0 => x"00002804",
			1 => x"0106000d",
			2 => x"fea4000d",
			3 => x"00002804",
			4 => x"00400019",
			5 => x"ffbe0019",
			6 => x"00002808",
			7 => x"08001904",
			8 => x"0212002d",
			9 => x"0350002d",
			10 => x"fe34002d",
			11 => x"00002808",
			12 => x"08001904",
			13 => x"ffdb0041",
			14 => x"01b70041",
			15 => x"fe5e0041",
			16 => x"00002808",
			17 => x"05000d04",
			18 => x"ff800055",
			19 => x"01a30055",
			20 => x"fe620055",
			21 => x"00002808",
			22 => x"0b001804",
			23 => x"ff530069",
			24 => x"016a0069",
			25 => x"fe780069",
			26 => x"00002808",
			27 => x"08001904",
			28 => x"ff85007d",
			29 => x"0145007d",
			30 => x"fe87007d",
			31 => x"00002808",
			32 => x"08001904",
			33 => x"ffce0091",
			34 => x"00c40091",
			35 => x"fef10091",
			36 => x"02002508",
			37 => x"03000c04",
			38 => x"ffd900a5",
			39 => x"009100a5",
			40 => x"ff3700a5",
			41 => x"00002808",
			42 => x"08001904",
			43 => x"ffdb00b9",
			44 => x"008a00b9",
			45 => x"ff4d00b9",
			46 => x"02002508",
			47 => x"0a000b04",
			48 => x"000200cd",
			49 => x"007a00cd",
			50 => x"ff6100cd",
			51 => x"00002808",
			52 => x"0a000b04",
			53 => x"ffe000e1",
			54 => x"006700e1",
			55 => x"ff8000e1",
			56 => x"00002808",
			57 => x"0b001804",
			58 => x"ffe000f5",
			59 => x"005e00f5",
			60 => x"ff8e00f5",
			61 => x"00002808",
			62 => x"08001904",
			63 => x"ffe80109",
			64 => x"00570109",
			65 => x"ff9f0109",
			66 => x"00002808",
			67 => x"08001904",
			68 => x"ffeb011d",
			69 => x"0052011d",
			70 => x"ffaa011d",
			71 => x"00002808",
			72 => x"08001904",
			73 => x"ffed0131",
			74 => x"00460131",
			75 => x"ffb80131",
			76 => x"00002808",
			77 => x"0a000b04",
			78 => x"fff50145",
			79 => x"003f0145",
			80 => x"ffc20145",
			81 => x"00002808",
			82 => x"08001904",
			83 => x"fff20159",
			84 => x"00390159",
			85 => x"ffcb0159",
			86 => x"00002808",
			87 => x"02002104",
			88 => x"ed5b016d",
			89 => x"eb2a016d",
			90 => x"e26a016d",
			91 => x"00002508",
			92 => x"08001904",
			93 => x"01dc0189",
			94 => x"022d0189",
			95 => x"00002c04",
			96 => x"ff860189",
			97 => x"fe4b0189",
			98 => x"00002504",
			99 => x"019a01a5",
			100 => x"09003404",
			101 => x"fe6401a5",
			102 => x"0b002804",
			103 => x"009301a5",
			104 => x"fecd01a5",
			105 => x"02002004",
			106 => x"019401c1",
			107 => x"0b002404",
			108 => x"fe6001c1",
			109 => x"00005c04",
			110 => x"017501c1",
			111 => x"fea701c1",
			112 => x"02002004",
			113 => x"018d01dd",
			114 => x"0b002404",
			115 => x"fe6701dd",
			116 => x"00005c04",
			117 => x"014901dd",
			118 => x"febe01dd",
			119 => x"02002004",
			120 => x"010801f9",
			121 => x"0b002104",
			122 => x"fe9d01f9",
			123 => x"00005c04",
			124 => x"008801f9",
			125 => x"ff8001f9",
			126 => x"02002004",
			127 => x"00d30215",
			128 => x"0b002404",
			129 => x"fec20215",
			130 => x"00005c04",
			131 => x"00540215",
			132 => x"ffc70215",
			133 => x"02002004",
			134 => x"00ba0231",
			135 => x"0b002404",
			136 => x"fedb0231",
			137 => x"00005c04",
			138 => x"004b0231",
			139 => x"ffcf0231",
			140 => x"02002004",
			141 => x"0095024d",
			142 => x"0b002404",
			143 => x"ff05024d",
			144 => x"00005c04",
			145 => x"0033024d",
			146 => x"ffde024d",
			147 => x"00002504",
			148 => x"00780269",
			149 => x"09003404",
			150 => x"ff660269",
			151 => x"0c002b04",
			152 => x"00090269",
			153 => x"fffb0269",
			154 => x"02002004",
			155 => x"004b0285",
			156 => x"0b002104",
			157 => x"ff8b0285",
			158 => x"00005c04",
			159 => x"00230285",
			160 => x"fff10285",
			161 => x"02002004",
			162 => x"003f02a1",
			163 => x"0b002104",
			164 => x"ffa002a1",
			165 => x"00005c04",
			166 => x"001e02a1",
			167 => x"fff302a1",
			168 => x"02002004",
			169 => x"002f02bd",
			170 => x"0b002104",
			171 => x"ffb902bd",
			172 => x"00005c04",
			173 => x"001702bd",
			174 => x"fff802bd",
			175 => x"02002004",
			176 => x"002d02d9",
			177 => x"09003004",
			178 => x"ffbe02d9",
			179 => x"08002b04",
			180 => x"000b02d9",
			181 => x"ffff02d9",
			182 => x"00002508",
			183 => x"0b001804",
			184 => x"016602fd",
			185 => x"01e402fd",
			186 => x"09003404",
			187 => x"fe5302fd",
			188 => x"0a003904",
			189 => x"00d002fd",
			190 => x"fe6802fd",
			191 => x"00002508",
			192 => x"08001904",
			193 => x"00f50321",
			194 => x"01c20321",
			195 => x"09003604",
			196 => x"fe5a0321",
			197 => x"09003a04",
			198 => x"ffff0321",
			199 => x"fe8a0321",
			200 => x"00002508",
			201 => x"02002004",
			202 => x"019f0345",
			203 => x"00120345",
			204 => x"09003404",
			205 => x"fe630345",
			206 => x"0c002b04",
			207 => x"00dd0345",
			208 => x"febe0345",
			209 => x"02002004",
			210 => x"01210369",
			211 => x"0b002408",
			212 => x"0d002104",
			213 => x"fe920369",
			214 => x"ffd90369",
			215 => x"00005c04",
			216 => x"00860369",
			217 => x"ff990369",
			218 => x"02002004",
			219 => x"017a0395",
			220 => x"0b00240c",
			221 => x"0b002104",
			222 => x"fe6e0395",
			223 => x"0b002204",
			224 => x"ffec0395",
			225 => x"ff7c0395",
			226 => x"00005c04",
			227 => x"011e0395",
			228 => x"ff030395",
			229 => x"02002004",
			230 => x"014203c1",
			231 => x"0b00240c",
			232 => x"0b002104",
			233 => x"fe8203c1",
			234 => x"0b002204",
			235 => x"fffa03c1",
			236 => x"ffbf03c1",
			237 => x"00005c04",
			238 => x"00b703c1",
			239 => x"ff6603c1",
			240 => x"02002004",
			241 => x"016903f7",
			242 => x"0b002410",
			243 => x"0b002104",
			244 => x"fe7403f7",
			245 => x"0b002208",
			246 => x"0d002104",
			247 => x"ffd303f7",
			248 => x"002703f7",
			249 => x"ff9003f7",
			250 => x"00005c04",
			251 => x"00f803f7",
			252 => x"ff2f03f7",
			253 => x"00002804",
			254 => x"00fb0401",
			255 => x"feab0401",
			256 => x"00002808",
			257 => x"07002704",
			258 => x"04840415",
			259 => x"05660415",
			260 => x"fe200415",
			261 => x"00002504",
			262 => x"02530429",
			263 => x"00002c04",
			264 => x"ff7d0429",
			265 => x"fe460429",
			266 => x"00002808",
			267 => x"08001904",
			268 => x"000d043d",
			269 => x"01b2043d",
			270 => x"fe5f043d",
			271 => x"00002808",
			272 => x"05000d04",
			273 => x"ff8e0451",
			274 => x"01a10451",
			275 => x"fe630451",
			276 => x"00002808",
			277 => x"08001904",
			278 => x"ff820465",
			279 => x"01650465",
			280 => x"fe7a0465",
			281 => x"00002808",
			282 => x"08001904",
			283 => x"ff8f0479",
			284 => x"013c0479",
			285 => x"fe8c0479",
			286 => x"00002808",
			287 => x"08001904",
			288 => x"ffd1048d",
			289 => x"00bc048d",
			290 => x"fefa048d",
			291 => x"02002508",
			292 => x"03000c04",
			293 => x"ffdb04a1",
			294 => x"008c04a1",
			295 => x"ff3f04a1",
			296 => x"00002808",
			297 => x"08001904",
			298 => x"ffe104b5",
			299 => x"008604b5",
			300 => x"ff5604b5",
			301 => x"00002808",
			302 => x"0b001804",
			303 => x"ffe004c9",
			304 => x"007804c9",
			305 => x"ff6f04c9",
			306 => x"00002808",
			307 => x"0a000b04",
			308 => x"ffe104dd",
			309 => x"006404dd",
			310 => x"ff8404dd",
			311 => x"00002808",
			312 => x"0a000b04",
			313 => x"ffe504f1",
			314 => x"005f04f1",
			315 => x"ff9304f1",
			316 => x"00002808",
			317 => x"08001904",
			318 => x"ffe90505",
			319 => x"00540505",
			320 => x"ffa20505",
			321 => x"00002808",
			322 => x"0b001804",
			323 => x"ffea0519",
			324 => x"00470519",
			325 => x"ffb50519",
			326 => x"00002808",
			327 => x"08001904",
			328 => x"ffed052d",
			329 => x"0044052d",
			330 => x"ffba052d",
			331 => x"00002808",
			332 => x"0a000b04",
			333 => x"fff00541",
			334 => x"003e0541",
			335 => x"ffc30541",
			336 => x"00002808",
			337 => x"08001904",
			338 => x"fff20555",
			339 => x"00380555",
			340 => x"ffcc0555",
			341 => x"02002508",
			342 => x"05000d04",
			343 => x"02100571",
			344 => x"02dc0571",
			345 => x"00002f04",
			346 => x"fec30571",
			347 => x"fe3b0571",
			348 => x"00002508",
			349 => x"02002004",
			350 => x"020e058d",
			351 => x"01ba058d",
			352 => x"02002b04",
			353 => x"ff96058d",
			354 => x"fe4f058d",
			355 => x"00002504",
			356 => x"019805a9",
			357 => x"09003404",
			358 => x"fe6505a9",
			359 => x"0b002804",
			360 => x"008b05a9",
			361 => x"fedb05a9",
			362 => x"02002004",
			363 => x"019205c5",
			364 => x"0b002404",
			365 => x"fe6205c5",
			366 => x"00005c04",
			367 => x"016805c5",
			368 => x"feab05c5",
			369 => x"02002004",
			370 => x"018b05e1",
			371 => x"0b002404",
			372 => x"fe6905e1",
			373 => x"00005c04",
			374 => x"013e05e1",
			375 => x"fec905e1",
			376 => x"02002004",
			377 => x"00e705fd",
			378 => x"0b002104",
			379 => x"feb405fd",
			380 => x"00005c04",
			381 => x"006b05fd",
			382 => x"ffa205fd",
			383 => x"02002004",
			384 => x"00ca0619",
			385 => x"0b002104",
			386 => x"fecc0619",
			387 => x"00005c04",
			388 => x"005f0619",
			389 => x"ffb30619",
			390 => x"02002004",
			391 => x"00b30635",
			392 => x"0b002404",
			393 => x"fee40635",
			394 => x"00005c04",
			395 => x"00480635",
			396 => x"ffd20635",
			397 => x"02002004",
			398 => x"00870651",
			399 => x"0b002404",
			400 => x"ff1b0651",
			401 => x"00005c04",
			402 => x"00340651",
			403 => x"ffdf0651",
			404 => x"02002004",
			405 => x"005a066d",
			406 => x"0b002104",
			407 => x"ff6a066d",
			408 => x"00005c04",
			409 => x"0029066d",
			410 => x"ffe9066d",
			411 => x"02002004",
			412 => x"00490689",
			413 => x"0b002104",
			414 => x"ff8f0689",
			415 => x"00005c04",
			416 => x"00230689",
			417 => x"fff10689",
			418 => x"02002004",
			419 => x"003b06a5",
			420 => x"0b002104",
			421 => x"ffa306a5",
			422 => x"00005c04",
			423 => x"001b06a5",
			424 => x"fff306a5",
			425 => x"02002004",
			426 => x"002e06c1",
			427 => x"0b002104",
			428 => x"ffbb06c1",
			429 => x"00005c04",
			430 => x"001706c1",
			431 => x"fff806c1",
			432 => x"02002004",
			433 => x"002b06dd",
			434 => x"0b002404",
			435 => x"ffc506dd",
			436 => x"08002a04",
			437 => x"000606dd",
			438 => x"ffff06dd",
			439 => x"00002508",
			440 => x"03000c04",
			441 => x"01440701",
			442 => x"01d50701",
			443 => x"09003404",
			444 => x"fe550701",
			445 => x"03003304",
			446 => x"00c00701",
			447 => x"fe6c0701",
			448 => x"00002508",
			449 => x"02002004",
			450 => x"01a80725",
			451 => x"008f0725",
			452 => x"09003404",
			453 => x"fe600725",
			454 => x"01001604",
			455 => x"00cd0725",
			456 => x"fe900725",
			457 => x"00002508",
			458 => x"02002004",
			459 => x"019c0749",
			460 => x"000a0749",
			461 => x"09003404",
			462 => x"fe640749",
			463 => x"07004104",
			464 => x"00cf0749",
			465 => x"fec90749",
			466 => x"02002004",
			467 => x"01840775",
			468 => x"0b00240c",
			469 => x"0b002104",
			470 => x"fe6a0775",
			471 => x"0b002204",
			472 => x"ffe00775",
			473 => x"ff5a0775",
			474 => x"00005c04",
			475 => x"01340775",
			476 => x"fee70775",
			477 => x"02002004",
			478 => x"017507a1",
			479 => x"0b00240c",
			480 => x"0b002104",
			481 => x"fe6f07a1",
			482 => x"0b002204",
			483 => x"fff107a1",
			484 => x"ff8307a1",
			485 => x"00005c04",
			486 => x"011107a1",
			487 => x"ff1707a1",
			488 => x"02002004",
			489 => x"012a07cf",
			490 => x"0b00240c",
			491 => x"0b002104",
			492 => x"fe8d07cf",
			493 => x"0b002204",
			494 => x"ffff07cf",
			495 => x"ffcf07cf",
			496 => x"00005c04",
			497 => x"008d07cf",
			498 => x"ff9107cf",
			499 => x"00002804",
			500 => x"004107d9",
			501 => x"ffbc07d9",
			502 => x"00002504",
			503 => x"040707ed",
			504 => x"00002c04",
			505 => x"ffce07ed",
			506 => x"fe2b07ed",
			507 => x"00002808",
			508 => x"08001904",
			509 => x"ffe30801",
			510 => x"01bd0801",
			511 => x"fe5c0801",
			512 => x"00002808",
			513 => x"08001904",
			514 => x"00020815",
			515 => x"01ad0815",
			516 => x"fe600815",
			517 => x"00002808",
			518 => x"08001904",
			519 => x"ff470829",
			520 => x"01750829",
			521 => x"fe730829",
			522 => x"00002808",
			523 => x"08001904",
			524 => x"ff8c083d",
			525 => x"015d083d",
			526 => x"fe7d083d",
			527 => x"00002808",
			528 => x"0d001304",
			529 => x"ff910851",
			530 => x"011e0851",
			531 => x"fe990851",
			532 => x"00002808",
			533 => x"08001904",
			534 => x"ffd10865",
			535 => x"00a70865",
			536 => x"ff170865",
			537 => x"00002808",
			538 => x"08001904",
			539 => x"ffd90879",
			540 => x"008f0879",
			541 => x"ff450879",
			542 => x"00002808",
			543 => x"0b001804",
			544 => x"ffe1088d",
			545 => x"0082088d",
			546 => x"ff5e088d",
			547 => x"00002808",
			548 => x"0a000b04",
			549 => x"ffdf08a1",
			550 => x"007308a1",
			551 => x"ff7508a1",
			552 => x"00002808",
			553 => x"0b001804",
			554 => x"ffe008b5",
			555 => x"006108b5",
			556 => x"ff8a08b5",
			557 => x"00002808",
			558 => x"0a000b04",
			559 => x"ffe508c9",
			560 => x"005c08c9",
			561 => x"ff9708c9",
			562 => x"00002808",
			563 => x"08001904",
			564 => x"ffea08dd",
			565 => x"005308dd",
			566 => x"ffa708dd",
			567 => x"00002808",
			568 => x"0b001804",
			569 => x"ffea08f1",
			570 => x"004508f1",
			571 => x"ffb708f1",
			572 => x"00002808",
			573 => x"0a000b04",
			574 => x"fff40905",
			575 => x"00400905",
			576 => x"ffc00905",
			577 => x"00002808",
			578 => x"0a000b04",
			579 => x"fff00919",
			580 => x"003d0919",
			581 => x"ffc40919",
			582 => x"00002808",
			583 => x"08001904",
			584 => x"fff4092d",
			585 => x"0036092d",
			586 => x"ffd1092d",
			587 => x"02002508",
			588 => x"08001904",
			589 => x"01cc0949",
			590 => x"028d0949",
			591 => x"00002f04",
			592 => x"fed90949",
			593 => x"fe410949",
			594 => x"00002508",
			595 => x"02002004",
			596 => x"01f70965",
			597 => x"01970965",
			598 => x"02002b04",
			599 => x"ff9a0965",
			600 => x"fe520965",
			601 => x"02002004",
			602 => x"01960981",
			603 => x"0b002404",
			604 => x"fe5e0981",
			605 => x"00005c04",
			606 => x"017c0981",
			607 => x"fe9f0981",
			608 => x"02002004",
			609 => x"0190099d",
			610 => x"0b002404",
			611 => x"fe65099d",
			612 => x"00005c04",
			613 => x"015d099d",
			614 => x"feb6099d",
			615 => x"02002004",
			616 => x"018809b9",
			617 => x"0b002404",
			618 => x"fe6c09b9",
			619 => x"00005c04",
			620 => x"014009b9",
			621 => x"feda09b9",
			622 => x"02002004",
			623 => x"00dc09d5",
			624 => x"09003004",
			625 => x"febb09d5",
			626 => x"00006504",
			627 => x"005409d5",
			628 => x"ffcc09d5",
			629 => x"02002004",
			630 => x"00c209f1",
			631 => x"0b002104",
			632 => x"fed509f1",
			633 => x"00005c04",
			634 => x"005c09f1",
			635 => x"ffb609f1",
			636 => x"02002004",
			637 => x"009c0a0d",
			638 => x"0b002404",
			639 => x"fefb0a0d",
			640 => x"00005c04",
			641 => x"00340a0d",
			642 => x"ffdd0a0d",
			643 => x"02002004",
			644 => x"00830a29",
			645 => x"0b002404",
			646 => x"ff240a29",
			647 => x"00005c04",
			648 => x"00320a29",
			649 => x"ffe10a29",
			650 => x"02002004",
			651 => x"00570a45",
			652 => x"0b002104",
			653 => x"ff700a45",
			654 => x"00005c04",
			655 => x"00280a45",
			656 => x"ffea0a45",
			657 => x"02002004",
			658 => x"00410a61",
			659 => x"0b002104",
			660 => x"ff9d0a61",
			661 => x"00005c04",
			662 => x"001f0a61",
			663 => x"fff30a61",
			664 => x"02002004",
			665 => x"003a0a7d",
			666 => x"0b002104",
			667 => x"ffa60a7d",
			668 => x"00005c04",
			669 => x"001b0a7d",
			670 => x"fff40a7d",
			671 => x"02002004",
			672 => x"002d0a99",
			673 => x"09003004",
			674 => x"ffbc0a99",
			675 => x"08002b04",
			676 => x"000b0a99",
			677 => x"ffff0a99",
			678 => x"02002004",
			679 => x"002a0ab5",
			680 => x"0b002404",
			681 => x"ffc70ab5",
			682 => x"08002a04",
			683 => x"00060ab5",
			684 => x"ffff0ab5",
			685 => x"00002508",
			686 => x"08001904",
			687 => x"01140ad9",
			688 => x"01cb0ad9",
			689 => x"09003604",
			690 => x"fe580ad9",
			691 => x"09003a04",
			692 => x"fff80ad9",
			693 => x"fe800ad9",
			694 => x"00002508",
			695 => x"0a000b04",
			696 => x"00660afd",
			697 => x"01a40afd",
			698 => x"09003404",
			699 => x"fe610afd",
			700 => x"01001604",
			701 => x"00bf0afd",
			702 => x"fe980afd",
			703 => x"00002508",
			704 => x"0a000b04",
			705 => x"ffe30b21",
			706 => x"009c0b21",
			707 => x"09003404",
			708 => x"ff1c0b21",
			709 => x"0c002b04",
			710 => x"00140b21",
			711 => x"fff50b21",
			712 => x"02002004",
			713 => x"017f0b4d",
			714 => x"0b00240c",
			715 => x"0b002104",
			716 => x"fe6c0b4d",
			717 => x"0b002204",
			718 => x"ffe60b4d",
			719 => x"ff700b4d",
			720 => x"00005c04",
			721 => x"012a0b4d",
			722 => x"fef50b4d",
			723 => x"02002004",
			724 => x"014b0b79",
			725 => x"0b00240c",
			726 => x"0b002104",
			727 => x"fe7f0b79",
			728 => x"0b002204",
			729 => x"fff90b79",
			730 => x"ffba0b79",
			731 => x"00005c04",
			732 => x"00c20b79",
			733 => x"ff5d0b79",
			734 => x"02002004",
			735 => x"00f00ba7",
			736 => x"0b00240c",
			737 => x"0d002104",
			738 => x"fead0ba7",
			739 => x"0d002204",
			740 => x"00030ba7",
			741 => x"ffe50ba7",
			742 => x"00005c04",
			743 => x"00630ba7",
			744 => x"ffbc0ba7",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(253, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(499, initial_addr_3'length));
	end generate gen_rom_12;

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
