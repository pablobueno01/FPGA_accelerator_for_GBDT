-------------------------------------------------------------------------------
-- Synchronous ROM with generic memory and data sizes
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
    generic(ADDRESS_BITS: positive;
            DATA_LENGTH:  positive;
            SELECT_ROM:  integer := 0); -- Select which ROM to use
    port(-- Control signals
         Clk: in std_logic;
         Re:  in std_logic;
         
         -- Input signals
         Addr: in std_logic_vector (ADDRESS_BITS - 1 downto 0);
         
         -- Output
         Dout: out std_logic_vector (DATA_LENGTH - 1 downto 0);
         initial_addr_2: out std_logic_vector (ADDRESS_BITS - 1 downto 0);
         initial_addr_3: out std_logic_vector (ADDRESS_BITS - 1 downto 0));
end rom;

architecture Behavioral of rom is

    type MemoryBank is array(0 to 2**ADDRESS_BITS - 1)
                    of std_logic_vector(DATA_LENGTH - 1 downto 0);
    signal bank: MemoryBank;


begin

	gen_rom_0: if SELECT_ROM = 0 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000000000000001110101",
			29 => "0000000000000001111001",
			30 => "0000000000000001111101",
			31 => "0000000000000010000001",
			32 => "0000000000000010000101",
			33 => "0000000000000010001001",
			34 => "0000000000000010001101",
			35 => "0000000000000010010001",
			36 => "0000000000000010010101",
			37 => "0011111010111000000100",
			38 => "0000000000000010100001",
			39 => "0000000000000010100001",
			40 => "0011110000001100000100",
			41 => "0000000000000010101101",
			42 => "0000000000000010101101",
			43 => "0000001100100100000100",
			44 => "0000000000000010111001",
			45 => "0000000000000010111001",
			46 => "0000001100100100000100",
			47 => "0000000000000011000101",
			48 => "0000000000000011000101",
			49 => "0011110000001100000100",
			50 => "0000000000000011010001",
			51 => "0000000000000011010001",
			52 => "0011110111001000001000",
			53 => "0011101001101000000100",
			54 => "0000000000000011100101",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0000000110100000001000",
			58 => "0011111100101100000100",
			59 => "0000000000000100000001",
			60 => "0000000000000100000001",
			61 => "0011101001101000000100",
			62 => "0000000000000100000001",
			63 => "0000000000000100000001",
			64 => "0000000101100100000100",
			65 => "0000000000000100011101",
			66 => "0001101100011000001000",
			67 => "0010011100100000000100",
			68 => "0000000000000100011101",
			69 => "0000000000000100011101",
			70 => "0000000000000100011101",
			71 => "0010011100100000001100",
			72 => "0001101100011000001000",
			73 => "0001010100011000000100",
			74 => "0000000000000100111001",
			75 => "0000000000000100111001",
			76 => "0000000000000100111001",
			77 => "0000000000000100111001",
			78 => "0000011110011100001100",
			79 => "0011101100011100000100",
			80 => "0000000000000101010101",
			81 => "0011111010111000000100",
			82 => "0000000000000101010101",
			83 => "0000000000000101010101",
			84 => "0000000000000101010101",
			85 => "0011111010111000001100",
			86 => "0011001110001100000100",
			87 => "0000000000000101110001",
			88 => "0011001101010100000100",
			89 => "0000000000000101110001",
			90 => "0000000000000101110001",
			91 => "0000000000000101110001",
			92 => "0011111010111000001100",
			93 => "0011001101010100001000",
			94 => "0011001100110000000100",
			95 => "0000000000000110001101",
			96 => "0000000000000110001101",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0010011100100000001100",
			100 => "0011111010111000001000",
			101 => "0000000101100100000100",
			102 => "0000000000000110101001",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0000000110100000001000",
			107 => "0010011100100000000100",
			108 => "0000000000000111001101",
			109 => "1111111000000111001101",
			110 => "0011000100001000001000",
			111 => "0000101110110100000100",
			112 => "0000000000000111001101",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0001000010100000000100",
			116 => "1111111000000111110001",
			117 => "0000101110010000001100",
			118 => "0000110001110100000100",
			119 => "0000000000000111110001",
			120 => "0010011100100000000100",
			121 => "0000001000000111110001",
			122 => "0000000000000111110001",
			123 => "0000000000000111110001",
			124 => "0000011110011100010000",
			125 => "0011001101010100001100",
			126 => "0001011110110000000100",
			127 => "0000000000001000010101",
			128 => "0011111010111000000100",
			129 => "0000000000001000010101",
			130 => "0000000000001000010101",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0011111010111000010000",
			134 => "0001110111001000001100",
			135 => "0011001100110000000100",
			136 => "0000000000001000111001",
			137 => "0010011100100000000100",
			138 => "0000000000001000111001",
			139 => "0000000000001000111001",
			140 => "0000000000001000111001",
			141 => "0000000000001000111001",
			142 => "0000011110011100010000",
			143 => "0011000001111100001100",
			144 => "0001110110000100000100",
			145 => "0000000000001001011101",
			146 => "0011111010111000000100",
			147 => "0000000000001001011101",
			148 => "0000000000001001011101",
			149 => "0000000000001001011101",
			150 => "0000000000001001011101",
			151 => "0011110111001000010000",
			152 => "0011101001101000000100",
			153 => "0000000000001010000001",
			154 => "0010011100100000001000",
			155 => "0011001101010100000100",
			156 => "0000000000001010000001",
			157 => "0000000000001010000001",
			158 => "0000000000001010000001",
			159 => "0000000000001010000001",
			160 => "0010011100100000010000",
			161 => "0011001110001100000100",
			162 => "0000000000001010100101",
			163 => "0011001101010100001000",
			164 => "0011110111001000000100",
			165 => "0000000000001010100101",
			166 => "0000000000001010100101",
			167 => "0000000000001010100101",
			168 => "0000000000001010100101",
			169 => "0000000010110100001000",
			170 => "0010011100100000000100",
			171 => "0000000000001011010001",
			172 => "0000000000001011010001",
			173 => "0011101001101000000100",
			174 => "0000000000001011010001",
			175 => "0011001101010100001000",
			176 => "0010011100100000000100",
			177 => "0000000000001011010001",
			178 => "0000000000001011010001",
			179 => "0000000000001011010001",
			180 => "0000000101100100000100",
			181 => "1111111000001011111101",
			182 => "0000011110011100001100",
			183 => "0011110111001000001000",
			184 => "0000101001100000000100",
			185 => "0000001000001011111101",
			186 => "0000000000001011111101",
			187 => "0000000000001011111101",
			188 => "0011110000001100000100",
			189 => "0000000000001011111101",
			190 => "0000000000001011111101",
			191 => "0000001101000100001100",
			192 => "0000011110011100001000",
			193 => "0011101011010100000100",
			194 => "1111111000001100110001",
			195 => "0000001000001100110001",
			196 => "1111111000001100110001",
			197 => "0000101100010100000100",
			198 => "0000001000001100110001",
			199 => "0001000001100000000100",
			200 => "1111111000001100110001",
			201 => "0000101110110100000100",
			202 => "0000001000001100110001",
			203 => "0000000000001100110001",
			204 => "0000001100100100001100",
			205 => "0010011100100000001000",
			206 => "0000110111000000000100",
			207 => "1111111000001101101101",
			208 => "0000010000001101101101",
			209 => "1111111000001101101101",
			210 => "0000100110010000001100",
			211 => "0011111010111100001000",
			212 => "0011110100001000000100",
			213 => "0000001000001101101101",
			214 => "0000001000001101101101",
			215 => "0000011000001101101101",
			216 => "0001111101010100000100",
			217 => "0000001000001101101101",
			218 => "1111111000001101101101",
			219 => "0000000010110100001000",
			220 => "0010011100100000000100",
			221 => "0000000000001110100001",
			222 => "1111111000001110100001",
			223 => "0011110000001100000100",
			224 => "0000001000001110100001",
			225 => "0001101100011000001000",
			226 => "0000100010000100000100",
			227 => "0000001000001110100001",
			228 => "0000000000001110100001",
			229 => "0010100010111100000100",
			230 => "1111111000001110100001",
			231 => "0000001000001110100001",
			232 => "0000000010110100001000",
			233 => "0010011100100000000100",
			234 => "0000000000001111011101",
			235 => "1111111000001111011101",
			236 => "0011000100001000001100",
			237 => "0000101110110100001000",
			238 => "0000000110100000000100",
			239 => "0000000000001111011101",
			240 => "0000001000001111011101",
			241 => "0000000000001111011101",
			242 => "0000100011001000000100",
			243 => "0000000000001111011101",
			244 => "0001101100011000000100",
			245 => "0000000000001111011101",
			246 => "0000000000001111011101",
			247 => "0010000101101100001000",
			248 => "0010011100100000000100",
			249 => "0000000000010000010001",
			250 => "1111111000010000010001",
			251 => "0000101100010100000100",
			252 => "0000001000010000010001",
			253 => "0001101100011000000100",
			254 => "0000001000010000010001",
			255 => "0010100010111100001000",
			256 => "0010111010111100000100",
			257 => "0000000000010000010001",
			258 => "1111111000010000010001",
			259 => "0000000000010000010001",
			260 => "0000000110100000001000",
			261 => "0011110000001100000100",
			262 => "0000000000010001000101",
			263 => "0000000000010001000101",
			264 => "0001110111001000010000",
			265 => "0011110111001000001100",
			266 => "0010011100100000000100",
			267 => "0000000000010001000101",
			268 => "0010011100100000000100",
			269 => "0000000000010001000101",
			270 => "0000000000010001000101",
			271 => "0000000000010001000101",
			272 => "0000000000010001000101",
			273 => "0000000010110100001000",
			274 => "0010011100100000000100",
			275 => "0000000000010001111001",
			276 => "0000000000010001111001",
			277 => "0011101001101000000100",
			278 => "0000000000010001111001",
			279 => "0011001101010100001100",
			280 => "0011110111001000001000",
			281 => "0010011100100000000100",
			282 => "0000000000010001111001",
			283 => "0000000000010001111001",
			284 => "0000000000010001111001",
			285 => "0000000000010001111001",
			286 => "0010011100100000010100",
			287 => "0001110111001000010000",
			288 => "0001011110110000000100",
			289 => "0000000000010010100101",
			290 => "0011111010111000001000",
			291 => "0010111110110000000100",
			292 => "0000000000010010100101",
			293 => "0000000000010010100101",
			294 => "0000000000010010100101",
			295 => "0000000000010010100101",
			296 => "0000000000010010100101",
			297 => "0011111010111000010100",
			298 => "0011101001101000000100",
			299 => "0000000000010011010001",
			300 => "0011001101010100001100",
			301 => "0000011110011100001000",
			302 => "0000011110011100000100",
			303 => "0000000000010011010001",
			304 => "0000000000010011010001",
			305 => "0000000000010011010001",
			306 => "0000000000010011010001",
			307 => "0000000000010011010001",
			308 => "0000001101000100001100",
			309 => "0010011100100000001000",
			310 => "0000111111001000000100",
			311 => "1111111000010100010101",
			312 => "0000001000010100010101",
			313 => "1111111000010100010101",
			314 => "0000100010000000001100",
			315 => "0001000000100100000100",
			316 => "0000001000010100010101",
			317 => "0000000111100000000100",
			318 => "0000001000010100010101",
			319 => "0000001000010100010101",
			320 => "0001101100011000000100",
			321 => "0000010000010100010101",
			322 => "0011011000011000000100",
			323 => "0000001000010100010101",
			324 => "1111111000010100010101",
			325 => "0000001100100100001100",
			326 => "0010011100100000001000",
			327 => "0000110111000000000100",
			328 => "1111111000010101011001",
			329 => "0000010000010101011001",
			330 => "1111111000010101011001",
			331 => "0000100110010000010000",
			332 => "0011101011010100001100",
			333 => "0000110010111100000100",
			334 => "0000001000010101011001",
			335 => "0011110001111100000100",
			336 => "0000001000010101011001",
			337 => "1111111000010101011001",
			338 => "0000010000010101011001",
			339 => "0001101010011000000100",
			340 => "0000001000010101011001",
			341 => "1111111000010101011001",
			342 => "0000000010110100001000",
			343 => "0010011100100000000100",
			344 => "0000000000010110011101",
			345 => "1111111000010110011101",
			346 => "0011000100001000001100",
			347 => "0000101110110100001000",
			348 => "0000000110100000000100",
			349 => "0000000000010110011101",
			350 => "0000001000010110011101",
			351 => "0000000000010110011101",
			352 => "0000100011001000000100",
			353 => "0000000000010110011101",
			354 => "0001101100011000000100",
			355 => "0000000000010110011101",
			356 => "0011011000011000000100",
			357 => "0000000000010110011101",
			358 => "0000000000010110011101",
			359 => "0000001101000100001100",
			360 => "0010011100100000001000",
			361 => "0000111111001000000100",
			362 => "1111111000010111101001",
			363 => "0000001000010111101001",
			364 => "1111111000010111101001",
			365 => "0000100010000000010000",
			366 => "0001000000100100000100",
			367 => "0000001000010111101001",
			368 => "0011110000001100000100",
			369 => "0000001000010111101001",
			370 => "0000000111100000000100",
			371 => "0000000000010111101001",
			372 => "0000001000010111101001",
			373 => "0001101100011000000100",
			374 => "0000001000010111101001",
			375 => "0011011000011000000100",
			376 => "0000000000010111101001",
			377 => "1111111000010111101001",
			378 => "0010011100100000011000",
			379 => "0001011110110000000100",
			380 => "0000000000011000100101",
			381 => "0000101100010100000100",
			382 => "0000001000011000100101",
			383 => "0011010100000100001000",
			384 => "0000011110011100000100",
			385 => "0000000000011000100101",
			386 => "0000000000011000100101",
			387 => "0011010000011100000100",
			388 => "0000000000011000100101",
			389 => "0000000000011000100101",
			390 => "0010100010111100000100",
			391 => "1111111000011000100101",
			392 => "0000000000011000100101",
			393 => "0010011100100000011000",
			394 => "0001110111001000010100",
			395 => "0001011110110000000100",
			396 => "0000000000011001100001",
			397 => "0011110111001000001100",
			398 => "0000011110011100001000",
			399 => "0000101001100000000100",
			400 => "0000001000011001100001",
			401 => "0000000000011001100001",
			402 => "0000000000011001100001",
			403 => "0000000000011001100001",
			404 => "0000000000011001100001",
			405 => "0010100010111100000100",
			406 => "1111111000011001100001",
			407 => "0000000000011001100001",
			408 => "0010011100100000011100",
			409 => "0001010100011000000100",
			410 => "1111111000011010100101",
			411 => "0011110000001100000100",
			412 => "0000001000011010100101",
			413 => "0001101100011000001000",
			414 => "0000000111100000000100",
			415 => "0000000000011010100101",
			416 => "0000001000011010100101",
			417 => "0001110001111100000100",
			418 => "0000001000011010100101",
			419 => "0010100010111100000100",
			420 => "1111111000011010100101",
			421 => "0000000000011010100101",
			422 => "0010100010111100000100",
			423 => "1111111000011010100101",
			424 => "0000000000011010100101",
			425 => "0000001110101000001100",
			426 => "0010011100100000001000",
			427 => "0000000101100100000100",
			428 => "1111111000011011111001",
			429 => "0000001000011011111001",
			430 => "1111111000011011111001",
			431 => "0010011100100000011000",
			432 => "0011010100000100010100",
			433 => "0000110010111100001000",
			434 => "0011110100001000000100",
			435 => "0000001000011011111001",
			436 => "0000001000011011111001",
			437 => "0001101010011000000100",
			438 => "0000001000011011111001",
			439 => "0000100110010000000100",
			440 => "0000000000011011111001",
			441 => "1111111000011011111001",
			442 => "0000010000011011111001",
			443 => "0000100010000000000100",
			444 => "0000001000011011111001",
			445 => "1111111000011011111001",
			446 => "0010011100100000100100",
			447 => "0000000110100000010000",
			448 => "0011101011010100001000",
			449 => "0010011100100000000100",
			450 => "0000000000011101001101",
			451 => "0000000000011101001101",
			452 => "0001100100110100000100",
			453 => "0000000000011101001101",
			454 => "0000000000011101001101",
			455 => "0001101101111100000100",
			456 => "0000010000011101001101",
			457 => "0011001010111100001100",
			458 => "0000001101000100000100",
			459 => "0000000000011101001101",
			460 => "0011111010111000000100",
			461 => "0000001000011101001101",
			462 => "0000000000011101001101",
			463 => "0000000000011101001101",
			464 => "0010100010111100000100",
			465 => "1111111000011101001101",
			466 => "0000000000011101001101",
			467 => "0000001110101000010100",
			468 => "0000011110011100010000",
			469 => "0011101011010100001000",
			470 => "0000001001010100000100",
			471 => "1111111000011110101001",
			472 => "0000000000011110101001",
			473 => "0010101000110000000100",
			474 => "0000001000011110101001",
			475 => "0000000000011110101001",
			476 => "1111111000011110101001",
			477 => "0000101110110100011000",
			478 => "0011100110001000010100",
			479 => "0000110010111100001000",
			480 => "0011110100001000000100",
			481 => "0000001000011110101001",
			482 => "0000000000011110101001",
			483 => "0000000101001000001000",
			484 => "0000011110011100000100",
			485 => "1111111000011110101001",
			486 => "0000000000011110101001",
			487 => "0000000000011110101001",
			488 => "0000010000011110101001",
			489 => "1111111000011110101001",
			490 => "0010011100100000101100",
			491 => "0000011110011100100000",
			492 => "0000001101000100010000",
			493 => "0011101011010100001000",
			494 => "0010011100100000000100",
			495 => "0000000000100000001101",
			496 => "0000000000100000001101",
			497 => "0001100100110100000100",
			498 => "0000000000100000001101",
			499 => "0000000000100000001101",
			500 => "0011001101010100001100",
			501 => "0000011110011100001000",
			502 => "0000101110110100000100",
			503 => "0000001000100000001101",
			504 => "0000000000100000001101",
			505 => "0000000000100000001101",
			506 => "0000000000100000001101",
			507 => "0001011010001100000100",
			508 => "0000000000100000001101",
			509 => "0010000110000100000100",
			510 => "0000010000100000001101",
			511 => "0000000000100000001101",
			512 => "0010001101111000000100",
			513 => "1111111000100000001101",
			514 => "0000000000100000001101",
			515 => "0000000101100100000100",
			516 => "1111111000100001001011",
			517 => "0001110111001000011000",
			518 => "0010011100100000010100",
			519 => "0011110111001000010000",
			520 => "0000011110011100001100",
			521 => "0000101001100000001000",
			522 => "0011001100110000000100",
			523 => "0000000000100001001011",
			524 => "0000001000100001001011",
			525 => "0000000000100001001011",
			526 => "0000000000100001001011",
			527 => "0000000000100001001011",
			528 => "0000000000100001001011",
			529 => "0000000000100001001011",
			530 => "0000000000100001001101",
			531 => "0000000000100001010001",
			532 => "0000000000100001010101",
			533 => "0000000000100001011001",
			534 => "0000000000100001011101",
			535 => "0000000000100001100001",
			536 => "0000000000100001100101",
			537 => "0000000000100001101001",
			538 => "0000000000100001101101",
			539 => "0000000000100001110001",
			540 => "0000000000100001110101",
			541 => "0000000000100001111001",
			542 => "0000000000100001111101",
			543 => "0000000000100010000001",
			544 => "0000000000100010000101",
			545 => "0000000000100010001001",
			546 => "0000000000100010001101",
			547 => "0000000000100010010001",
			548 => "0000000000100010010101",
			549 => "0000000000100010011001",
			550 => "0000000000100010011101",
			551 => "0000000000100010100001",
			552 => "0000000000100010100101",
			553 => "0000000000100010101001",
			554 => "0000000000100010101101",
			555 => "0000000000100010110001",
			556 => "0000000000100010110101",
			557 => "0000000000100010111001",
			558 => "0000000000100010111101",
			559 => "0000000000100011000001",
			560 => "0000000000100011000101",
			561 => "0000000000100011001001",
			562 => "0000000000100011001101",
			563 => "0000000000100011010001",
			564 => "0000000000100011010101",
			565 => "0000000000100011011001",
			566 => "0000000000100011011101",
			567 => "0011111010111000000100",
			568 => "0000000000100011101001",
			569 => "0000000000100011101001",
			570 => "0011110000001100000100",
			571 => "0000000000100011110101",
			572 => "0000000000100011110101",
			573 => "0000001100100100000100",
			574 => "0000000000100100000001",
			575 => "0000000000100100000001",
			576 => "0000001100100100000100",
			577 => "0000000000100100001101",
			578 => "0000000000100100001101",
			579 => "0011110000001100000100",
			580 => "0000000000100100011001",
			581 => "0000000000100100011001",
			582 => "0000000110100000001000",
			583 => "0011110000001100000100",
			584 => "0000000000100100101101",
			585 => "0000000000100100101101",
			586 => "0000000000100100101101",
			587 => "0000000110100000001000",
			588 => "0011111100101100000100",
			589 => "0000000000100101001001",
			590 => "0000000000100101001001",
			591 => "0011101001101000000100",
			592 => "0000000000100101001001",
			593 => "0000000000100101001001",
			594 => "0000011110011100001100",
			595 => "0000101001100000001000",
			596 => "0001011110110000000100",
			597 => "0000000000100101100101",
			598 => "0000000000100101100101",
			599 => "0000000000100101100101",
			600 => "0000000000100101100101",
			601 => "0000000111100000001100",
			602 => "0011111110001100000100",
			603 => "0000000000100110000001",
			604 => "0010100010111100000100",
			605 => "0000000000100110000001",
			606 => "0000000000100110000001",
			607 => "0000000000100110000001",
			608 => "0000011110011100001100",
			609 => "0011101100011100000100",
			610 => "0000000000100110011101",
			611 => "0011111010111000000100",
			612 => "0000000000100110011101",
			613 => "0000000000100110011101",
			614 => "0000000000100110011101",
			615 => "0011111010111000001100",
			616 => "0011001101010100001000",
			617 => "0011001100110000000100",
			618 => "0000000000100110111001",
			619 => "0000000000100110111001",
			620 => "0000000000100110111001",
			621 => "0000000000100110111001",
			622 => "0010011100100000001100",
			623 => "0011111010111000001000",
			624 => "0010001011000100000100",
			625 => "0000000000100111010101",
			626 => "0000000000100111010101",
			627 => "0000000000100111010101",
			628 => "0000000000100111010101",
			629 => "0011111010111000001100",
			630 => "0001110110000100000100",
			631 => "0000000000100111110001",
			632 => "0000011110011100000100",
			633 => "0000000000100111110001",
			634 => "0000000000100111110001",
			635 => "0000000000100111110001",
			636 => "0000000110100000001000",
			637 => "0010011100100000000100",
			638 => "0000000000101000010101",
			639 => "1111111000101000010101",
			640 => "0011000100001000001000",
			641 => "0000101110110100000100",
			642 => "0000000000101000010101",
			643 => "0000000000101000010101",
			644 => "0000000000101000010101",
			645 => "0011111010111000010000",
			646 => "0001101100011000001100",
			647 => "0001110110000100000100",
			648 => "0000000000101000111001",
			649 => "0010011100100000000100",
			650 => "0000000000101000111001",
			651 => "0000000000101000111001",
			652 => "0000000000101000111001",
			653 => "1111111000101000111001",
			654 => "0000000101100100000100",
			655 => "0000000000101001011101",
			656 => "0001101100011000001100",
			657 => "0010011100100000001000",
			658 => "0001111101111000000100",
			659 => "0000000000101001011101",
			660 => "0000000000101001011101",
			661 => "0000000000101001011101",
			662 => "0000000000101001011101",
			663 => "0000011110011100010000",
			664 => "0011000001111100001100",
			665 => "0001110110000100000100",
			666 => "0000000000101010000001",
			667 => "0011111010111000000100",
			668 => "0000000000101010000001",
			669 => "0000000000101010000001",
			670 => "0000000000101010000001",
			671 => "0000000000101010000001",
			672 => "0011111010111000010000",
			673 => "0011000100001000001100",
			674 => "0001110111001000001000",
			675 => "0011001100110000000100",
			676 => "0000000000101010100101",
			677 => "0000000000101010100101",
			678 => "0000000000101010100101",
			679 => "0000000000101010100101",
			680 => "0000000000101010100101",
			681 => "0011110111001000010000",
			682 => "0011101001101000000100",
			683 => "0000000000101011001001",
			684 => "0011001101010100001000",
			685 => "0001111110001100000100",
			686 => "0000000000101011001001",
			687 => "0000000000101011001001",
			688 => "0000000000101011001001",
			689 => "0000000000101011001001",
			690 => "0010011100100000010000",
			691 => "0011001110001100000100",
			692 => "0000000000101011101101",
			693 => "0011001101010100001000",
			694 => "0011110111001000000100",
			695 => "0000000000101011101101",
			696 => "0000000000101011101101",
			697 => "0000000000101011101101",
			698 => "0000000000101011101101",
			699 => "0000000110100000001000",
			700 => "0011111100101100000100",
			701 => "0000000000101100011001",
			702 => "0000000000101100011001",
			703 => "0011101001101000000100",
			704 => "0000000000101100011001",
			705 => "0011001101010100001000",
			706 => "0011000000001100000100",
			707 => "0000000000101100011001",
			708 => "0000000000101100011001",
			709 => "0000000000101100011001",
			710 => "0010011100100000010100",
			711 => "0000101010001000001000",
			712 => "0001011110110000000100",
			713 => "0000000000101101000101",
			714 => "0000000000101101000101",
			715 => "0001110001111100000100",
			716 => "0000000000101101000101",
			717 => "0011010100000100000100",
			718 => "0000000000101101000101",
			719 => "0000000000101101000101",
			720 => "1111111000101101000101",
			721 => "0000011110011100010000",
			722 => "0001011110110000000100",
			723 => "0000000000101101111001",
			724 => "0011111010111100001000",
			725 => "0011001101010100000100",
			726 => "0000001000101101111001",
			727 => "0000000000101101111001",
			728 => "0000000000101101111001",
			729 => "0010100010011000000100",
			730 => "1111111000101101111001",
			731 => "0011110100001000000100",
			732 => "0000000000101101111001",
			733 => "0000000000101101111001",
			734 => "0000000010110100001000",
			735 => "0010011100100000000100",
			736 => "0000000000101110101101",
			737 => "1111111000101110101101",
			738 => "0011110000001100000100",
			739 => "0000001000101110101101",
			740 => "0001101100011000001000",
			741 => "0000100010000100000100",
			742 => "0000001000101110101101",
			743 => "0000000000101110101101",
			744 => "0010100010111100000100",
			745 => "1111111000101110101101",
			746 => "0000001000101110101101",
			747 => "0000000110100000001000",
			748 => "0010011100100000000100",
			749 => "0000000000101111100001",
			750 => "1111111000101111100001",
			751 => "0000100011001000000100",
			752 => "0000001000101111100001",
			753 => "0001111101010100001000",
			754 => "0001111010111100000100",
			755 => "0000000000101111100001",
			756 => "0000000000101111100001",
			757 => "0001101100011000000100",
			758 => "0000000000101111100001",
			759 => "0000000000101111100001",
			760 => "0000011110011100011000",
			761 => "0001101100011000001100",
			762 => "0001010100011000000100",
			763 => "0000000000110000011101",
			764 => "0010011100100000000100",
			765 => "0000001000110000011101",
			766 => "0000000000110000011101",
			767 => "0010100010111100001000",
			768 => "0000101010001000000100",
			769 => "0000000000110000011101",
			770 => "0000000000110000011101",
			771 => "0000000000110000011101",
			772 => "0010100010111100000100",
			773 => "1111111000110000011101",
			774 => "0000000000110000011101",
			775 => "0010011100100000010100",
			776 => "0001110111001000010000",
			777 => "0001011110110000000100",
			778 => "0000000000110001010001",
			779 => "0011110111001000001000",
			780 => "0000011110011100000100",
			781 => "0000001000110001010001",
			782 => "0000000000110001010001",
			783 => "0000000000110001010001",
			784 => "0000000000110001010001",
			785 => "0010100010111100000100",
			786 => "1111111000110001010001",
			787 => "0000000000110001010001",
			788 => "0010000101101100001000",
			789 => "0010011100100000000100",
			790 => "0000000000110010000101",
			791 => "0000000000110010000101",
			792 => "0001110111001000010000",
			793 => "0010011100100000000100",
			794 => "0000000000110010000101",
			795 => "0011110111001000001000",
			796 => "0010011100100000000100",
			797 => "0000000000110010000101",
			798 => "0000000000110010000101",
			799 => "0000000000110010000101",
			800 => "0000000000110010000101",
			801 => "0011001110001100001000",
			802 => "0010001110001100000100",
			803 => "0000000000110010111001",
			804 => "0000000000110010111001",
			805 => "0001110111001000010000",
			806 => "0010011100100000001100",
			807 => "0011000100001000001000",
			808 => "0011110111001000000100",
			809 => "0000000000110010111001",
			810 => "0000000000110010111001",
			811 => "0000000000110010111001",
			812 => "0000000000110010111001",
			813 => "0000000000110010111001",
			814 => "0000000101100100000100",
			815 => "0000000000110011100101",
			816 => "0001110111001000010000",
			817 => "0010011100100000001100",
			818 => "0000011110011100001000",
			819 => "0011001100110000000100",
			820 => "0000000000110011100101",
			821 => "0000000000110011100101",
			822 => "0000000000110011100101",
			823 => "0000000000110011100101",
			824 => "0000000000110011100101",
			825 => "0011111010111000010100",
			826 => "0010011100100000010000",
			827 => "0011001101010100001100",
			828 => "0001010100011000000100",
			829 => "0000000000110100010001",
			830 => "0000011110011100000100",
			831 => "0000000000110100010001",
			832 => "0000000000110100010001",
			833 => "0000000000110100010001",
			834 => "0000000000110100010001",
			835 => "0000000000110100010001",
			836 => "0000000101100100000100",
			837 => "1111111000110101000101",
			838 => "0000011110011100010000",
			839 => "0011001101010100001100",
			840 => "0011110111001000001000",
			841 => "0000101001100000000100",
			842 => "0000001000110101000101",
			843 => "0000000000110101000101",
			844 => "0000000000110101000101",
			845 => "0000000000110101000101",
			846 => "0011110000001100000100",
			847 => "0000000000110101000101",
			848 => "0000000000110101000101",
			849 => "0000001100100100001100",
			850 => "0010011100100000001000",
			851 => "0000110111000000000100",
			852 => "1111111000110110001001",
			853 => "0000001000110110001001",
			854 => "1111111000110110001001",
			855 => "0000100110010000010000",
			856 => "0011101011010100001100",
			857 => "0000110010111100000100",
			858 => "0000001000110110001001",
			859 => "0011110001111100000100",
			860 => "0000001000110110001001",
			861 => "1111111000110110001001",
			862 => "0000010000110110001001",
			863 => "0001111101010100000100",
			864 => "0000001000110110001001",
			865 => "1111111000110110001001",
			866 => "0000000010110100001000",
			867 => "0000011110011100000100",
			868 => "0000000000110111001101",
			869 => "1111111000110111001101",
			870 => "0011000100001000001100",
			871 => "0000101110110100001000",
			872 => "0000000110100000000100",
			873 => "0000000000110111001101",
			874 => "0000001000110111001101",
			875 => "0000000000110111001101",
			876 => "0000100011001000000100",
			877 => "0000000000110111001101",
			878 => "0001101100011000000100",
			879 => "0000000000110111001101",
			880 => "0011011000011000000100",
			881 => "0000000000110111001101",
			882 => "0000000000110111001101",
			883 => "0010011100100000011000",
			884 => "0001010100011000000100",
			885 => "0000000000111000001001",
			886 => "0011110000001100000100",
			887 => "0000001000111000001001",
			888 => "0001101100011000001000",
			889 => "0000000111100000000100",
			890 => "0000000000111000001001",
			891 => "0000001000111000001001",
			892 => "0001110001111100000100",
			893 => "0000001000111000001001",
			894 => "1111111000111000001001",
			895 => "0010100010111100000100",
			896 => "1111111000111000001001",
			897 => "0000000000111000001001",
			898 => "0000001101000100011000",
			899 => "0010011100100000010100",
			900 => "0001100111101000001000",
			901 => "0011111001110000000100",
			902 => "0000000000111001010101",
			903 => "0000001000111001010101",
			904 => "0000011110011100001000",
			905 => "0010011100100000000100",
			906 => "0000000000111001010101",
			907 => "0000000000111001010101",
			908 => "1111111000111001010101",
			909 => "1111111000111001010101",
			910 => "0000101100010100000100",
			911 => "0000001000111001010101",
			912 => "0001101100011000000100",
			913 => "0000001000111001010101",
			914 => "0001000011100100000100",
			915 => "1111111000111001010101",
			916 => "0000000000111001010101",
			917 => "0000000101100100000100",
			918 => "1111111000111010011001",
			919 => "0001101100011000001100",
			920 => "0010011100100000001000",
			921 => "0001111101111000000100",
			922 => "0000000000111010011001",
			923 => "0000000000111010011001",
			924 => "0000000000111010011001",
			925 => "0001110001111100001000",
			926 => "0000110010011000000100",
			927 => "0000000000111010011001",
			928 => "0000000000111010011001",
			929 => "0001101101011000001000",
			930 => "0000111111000100000100",
			931 => "0000000000111010011001",
			932 => "0000000000111010011001",
			933 => "0000000000111010011001",
			934 => "0010011100100000011100",
			935 => "0001010100011000000100",
			936 => "0000000000111011011101",
			937 => "0011110000001100000100",
			938 => "0000001000111011011101",
			939 => "0001101100011000001000",
			940 => "0000000111100000000100",
			941 => "0000000000111011011101",
			942 => "0000001000111011011101",
			943 => "0001110001111100000100",
			944 => "0000001000111011011101",
			945 => "0010100010111100000100",
			946 => "1111111000111011011101",
			947 => "0000000000111011011101",
			948 => "0010100010111100000100",
			949 => "1111111000111011011101",
			950 => "0000000000111011011101",
			951 => "0000001110101000010100",
			952 => "0000011110011100010000",
			953 => "0011101011010100001000",
			954 => "0000001001010100000100",
			955 => "1111111000111100110001",
			956 => "0000000000111100110001",
			957 => "0010101000110000000100",
			958 => "0000010000111100110001",
			959 => "0000000000111100110001",
			960 => "1111111000111100110001",
			961 => "0000101110110100010100",
			962 => "0011100110001000010000",
			963 => "0000101100010100000100",
			964 => "0000001000111100110001",
			965 => "0001101010011000000100",
			966 => "0000001000111100110001",
			967 => "0010110111001000000100",
			968 => "0000001000111100110001",
			969 => "1111111000111100110001",
			970 => "0000010000111100110001",
			971 => "1111111000111100110001",
			972 => "0000001100100100010100",
			973 => "0010011100100000001000",
			974 => "0000001001010100000100",
			975 => "1111111000111110001101",
			976 => "0000110000111110001101",
			977 => "0010100010011000000100",
			978 => "1111111000111110001101",
			979 => "0010001100110000000100",
			980 => "1111111000111110001101",
			981 => "0000001000111110001101",
			982 => "0000101110110100011000",
			983 => "0011110111001000010100",
			984 => "0011001010111100001100",
			985 => "0011110001111100001000",
			986 => "0011110100001000000100",
			987 => "0000010000111110001101",
			988 => "0000001000111110001101",
			989 => "0000101000111110001101",
			990 => "0000101100010100000100",
			991 => "0000010000111110001101",
			992 => "1111111000111110001101",
			993 => "0000101000111110001101",
			994 => "1111111000111110001101",
			995 => "0000001101000100001100",
			996 => "0010011100100000001000",
			997 => "0000111111001000000100",
			998 => "1111111000111111100001",
			999 => "0000001000111111100001",
			1000 => "1111111000111111100001",
			1001 => "0000101001100000011100",
			1002 => "0011001010111100010100",
			1003 => "0010011100100000010000",
			1004 => "0011110001111100001000",
			1005 => "0000101100010100000100",
			1006 => "0000001000111111100001",
			1007 => "0000000000111111100001",
			1008 => "0010001110001100000100",
			1009 => "0000011000111111100001",
			1010 => "0000001000111111100001",
			1011 => "1111111000111111100001",
			1012 => "0000101100010100000100",
			1013 => "0000001000111111100001",
			1014 => "1111111000111111100001",
			1015 => "1111111000111111100001",
			1016 => "0000000101001000101100",
			1017 => "0000001100100100011100",
			1018 => "0010011100100000001000",
			1019 => "0010100111000100000100",
			1020 => "1100101001000001000101",
			1021 => "1101111001000001000101",
			1022 => "0010011100100000001000",
			1023 => "0010100111000100000100",
			1024 => "1100101001000001000101",
			1025 => "1101011001000001000101",
			1026 => "0010100010011000000100",
			1027 => "1100101001000001000101",
			1028 => "0010100010111100000100",
			1029 => "1100110001000001000101",
			1030 => "1100101001000001000101",
			1031 => "0000101100010100000100",
			1032 => "1111010001000001000101",
			1033 => "0011000100001000000100",
			1034 => "1101100001000001000101",
			1035 => "0000100010000000000100",
			1036 => "1100111001000001000101",
			1037 => "1100101001000001000101",
			1038 => "0011111010111100000100",
			1039 => "1111011001000001000101",
			1040 => "1101011001000001000101",
			1041 => "0000001101000100001100",
			1042 => "0010011100100000001000",
			1043 => "0000111011010100000100",
			1044 => "1111111001000010011011",
			1045 => "0000001001000010011011",
			1046 => "1111111001000010011011",
			1047 => "0011110111001000011100",
			1048 => "0010011100100000011000",
			1049 => "0000001101000100000100",
			1050 => "0000010001000010011011",
			1051 => "0000000111100000001000",
			1052 => "0000101100010100000100",
			1053 => "0000001001000010011011",
			1054 => "1111111001000010011011",
			1055 => "0011010100000100001000",
			1056 => "0011011010011100000100",
			1057 => "0000001001000010011011",
			1058 => "0000001001000010011011",
			1059 => "0000001001000010011011",
			1060 => "0000000001000010011011",
			1061 => "1111111001000010011011",
			1062 => "0000000001000010011101",
			1063 => "0000000001000010100001",
			1064 => "0000000001000010100101",
			1065 => "0000000001000010101001",
			1066 => "0000000001000010101101",
			1067 => "0000000001000010110001",
			1068 => "0000000001000010110101",
			1069 => "0000000001000010111001",
			1070 => "0000000001000010111101",
			1071 => "0000000001000011000001",
			1072 => "0000000001000011000101",
			1073 => "0000000001000011001001",
			1074 => "0000000001000011001101",
			1075 => "0000000001000011010001",
			1076 => "0000000001000011010101",
			1077 => "0000000001000011011001",
			1078 => "0000000001000011011101",
			1079 => "0000000001000011100001",
			1080 => "0000000001000011100101",
			1081 => "0000000001000011101001",
			1082 => "0000000001000011101101",
			1083 => "0000000001000011110001",
			1084 => "0000000001000011110101",
			1085 => "0000000001000011111001",
			1086 => "0000000001000011111101",
			1087 => "0000000001000100000001",
			1088 => "0000000001000100000101",
			1089 => "0000000001000100001001",
			1090 => "0000000001000100001101",
			1091 => "0000000001000100010001",
			1092 => "0000000001000100010101",
			1093 => "0000000001000100011001",
			1094 => "0000000001000100011101",
			1095 => "0000000001000100100001",
			1096 => "0000000001000100100101",
			1097 => "0000000001000100101001",
			1098 => "0000000001000100101101",
			1099 => "0011111010111000000100",
			1100 => "0000000001000100111001",
			1101 => "0000000001000100111001",
			1102 => "0011110000001100000100",
			1103 => "0000000001000101000101",
			1104 => "0000000001000101000101",
			1105 => "0000001100100100000100",
			1106 => "0000000001000101010001",
			1107 => "0000000001000101010001",
			1108 => "0011110000001100000100",
			1109 => "0000000001000101011101",
			1110 => "0000000001000101011101",
			1111 => "0000001001010100000100",
			1112 => "1111111001000101110001",
			1113 => "0000101010001000000100",
			1114 => "0000000001000101110001",
			1115 => "0000000001000101110001",
			1116 => "0011110000001100000100",
			1117 => "0000000001000110000101",
			1118 => "0010011100100000000100",
			1119 => "0000000001000110000101",
			1120 => "0000000001000110000101",
			1121 => "0000000101100100000100",
			1122 => "1111111001000110100001",
			1123 => "0000101110010000001000",
			1124 => "0010011100100000000100",
			1125 => "0000001001000110100001",
			1126 => "0000000001000110100001",
			1127 => "0000000001000110100001",
			1128 => "0000011110011100001100",
			1129 => "0001011110110000000100",
			1130 => "0000000001000110111101",
			1131 => "0001101100011000000100",
			1132 => "0000000001000110111101",
			1133 => "0000000001000110111101",
			1134 => "0000000001000110111101",
			1135 => "0000000111100000001100",
			1136 => "0011111110001100000100",
			1137 => "0000000001000111011001",
			1138 => "0010100010111100000100",
			1139 => "0000000001000111011001",
			1140 => "0000000001000111011001",
			1141 => "0000000001000111011001",
			1142 => "0000011110011100001100",
			1143 => "0001000010100000000100",
			1144 => "0000000001000111110101",
			1145 => "0011111010111000000100",
			1146 => "0000000001000111110101",
			1147 => "0000000001000111110101",
			1148 => "0000000001000111110101",
			1149 => "0011111010111000001100",
			1150 => "0011001101010100001000",
			1151 => "0011001100110000000100",
			1152 => "0000000001001000010001",
			1153 => "0000000001001000010001",
			1154 => "0000000001001000010001",
			1155 => "0000000001001000010001",
			1156 => "0010011100100000001100",
			1157 => "0011111010111000001000",
			1158 => "0000000101100100000100",
			1159 => "0000000001001000101101",
			1160 => "0000000001001000101101",
			1161 => "0000000001001000101101",
			1162 => "0000000001001000101101",
			1163 => "0010011100100000001100",
			1164 => "0000101110010000001000",
			1165 => "0001010100011000000100",
			1166 => "0000000001001001010001",
			1167 => "0000001001001001010001",
			1168 => "0000000001001001010001",
			1169 => "0010100010111100000100",
			1170 => "1111111001001001010001",
			1171 => "0000000001001001010001",
			1172 => "0000000110100000001000",
			1173 => "0011111100101100000100",
			1174 => "0000000001001001110101",
			1175 => "1111111001001001110101",
			1176 => "0011000100001000001000",
			1177 => "0000101110110100000100",
			1178 => "0000000001001001110101",
			1179 => "0000000001001001110101",
			1180 => "0000000001001001110101",
			1181 => "0011111010111000010000",
			1182 => "0001101100011000001100",
			1183 => "0011001100110000000100",
			1184 => "0000000001001010011001",
			1185 => "0010011100100000000100",
			1186 => "0000000001001010011001",
			1187 => "0000000001001010011001",
			1188 => "0000000001001010011001",
			1189 => "0000000001001010011001",
			1190 => "0011111010111000010000",
			1191 => "0001110111001000001100",
			1192 => "0011001100110000000100",
			1193 => "0000000001001010111101",
			1194 => "0010011100100000000100",
			1195 => "0000000001001010111101",
			1196 => "0000000001001010111101",
			1197 => "0000000001001010111101",
			1198 => "0000000001001010111101",
			1199 => "0000011110011100010000",
			1200 => "0011000001111100001100",
			1201 => "0001011110110000000100",
			1202 => "0000000001001011100001",
			1203 => "0011111010111000000100",
			1204 => "0000000001001011100001",
			1205 => "0000000001001011100001",
			1206 => "0000000001001011100001",
			1207 => "0000000001001011100001",
			1208 => "0011111010111000010000",
			1209 => "0011101001101000000100",
			1210 => "0000000001001100000101",
			1211 => "0010011100100000001000",
			1212 => "0011001101010100000100",
			1213 => "0000000001001100000101",
			1214 => "0000000001001100000101",
			1215 => "0000000001001100000101",
			1216 => "0000000001001100000101",
			1217 => "0011110111001000010000",
			1218 => "0011101001101000000100",
			1219 => "0000000001001100101001",
			1220 => "0011001101010100001000",
			1221 => "0001111110001100000100",
			1222 => "0000000001001100101001",
			1223 => "0000000001001100101001",
			1224 => "0000000001001100101001",
			1225 => "0000000001001100101001",
			1226 => "0000000110100000001000",
			1227 => "0010011100100000000100",
			1228 => "0000000001001101010101",
			1229 => "1111111001001101010101",
			1230 => "0000100011001000000100",
			1231 => "0000001001001101010101",
			1232 => "0001010001101000000100",
			1233 => "0000000001001101010101",
			1234 => "0000110011010000000100",
			1235 => "0000000001001101010101",
			1236 => "0000000001001101010101",
			1237 => "0011001110001100001000",
			1238 => "0010001110001100000100",
			1239 => "0000000001001110000001",
			1240 => "0000000001001110000001",
			1241 => "0001110111001000001100",
			1242 => "0010011100100000001000",
			1243 => "0011000100001000000100",
			1244 => "0000000001001110000001",
			1245 => "0000000001001110000001",
			1246 => "0000000001001110000001",
			1247 => "0000000001001110000001",
			1248 => "0001001101110000000100",
			1249 => "1111111001001110101101",
			1250 => "0001101100011000001000",
			1251 => "0010011100100000000100",
			1252 => "0000000001001110101101",
			1253 => "0000000001001110101101",
			1254 => "0000101010001000000100",
			1255 => "0000000001001110101101",
			1256 => "0011111101111000000100",
			1257 => "0000000001001110101101",
			1258 => "0000000001001110101101",
			1259 => "0010011100100000010100",
			1260 => "0001101100011000001000",
			1261 => "0000000001001000000100",
			1262 => "0000000001001111100001",
			1263 => "0000000001001111100001",
			1264 => "0011111101111000000100",
			1265 => "0000000001001111100001",
			1266 => "0000000010011100000100",
			1267 => "0000000001001111100001",
			1268 => "0000000001001111100001",
			1269 => "0011110000001100000100",
			1270 => "0000000001001111100001",
			1271 => "1111111001001111100001",
			1272 => "0000000010110100001000",
			1273 => "0010011100100000000100",
			1274 => "0000000001010000010101",
			1275 => "1111111001010000010101",
			1276 => "0011110000001100000100",
			1277 => "0000001001010000010101",
			1278 => "0001101100011000001000",
			1279 => "0000100010000100000100",
			1280 => "0000001001010000010101",
			1281 => "0000000001010000010101",
			1282 => "0001110001111100000100",
			1283 => "0000001001010000010101",
			1284 => "1111111001010000010101",
			1285 => "0010000101101100001000",
			1286 => "0000011110011100000100",
			1287 => "0000000001010001001001",
			1288 => "1111111001010001001001",
			1289 => "0000100011001000000100",
			1290 => "0000001001010001001001",
			1291 => "0001111101010100001000",
			1292 => "0011000100001000000100",
			1293 => "0000000001010001001001",
			1294 => "0000000001010001001001",
			1295 => "0001101100011000000100",
			1296 => "0000000001010001001001",
			1297 => "0000000001010001001001",
			1298 => "0000011110011100011000",
			1299 => "0001101100011000001100",
			1300 => "0001010100011000000100",
			1301 => "0000000001010010000101",
			1302 => "0010011100100000000100",
			1303 => "0000001001010010000101",
			1304 => "0000000001010010000101",
			1305 => "0010100010111100001000",
			1306 => "0000101010001000000100",
			1307 => "0000000001010010000101",
			1308 => "0000000001010010000101",
			1309 => "0000000001010010000101",
			1310 => "0010100010111100000100",
			1311 => "1111111001010010000101",
			1312 => "0000000001010010000101",
			1313 => "0011111010111000011000",
			1314 => "0001101100011000001100",
			1315 => "0001111110001100000100",
			1316 => "0000000001010010111001",
			1317 => "0010011100100000000100",
			1318 => "0000000001010010111001",
			1319 => "0000000001010010111001",
			1320 => "0001110001111100001000",
			1321 => "0001010001101000000100",
			1322 => "0000000001010010111001",
			1323 => "0000000001010010111001",
			1324 => "0000000001010010111001",
			1325 => "1111111001010010111001",
			1326 => "0000000110100000001000",
			1327 => "0011110000001100000100",
			1328 => "0000000001010011101101",
			1329 => "0000000001010011101101",
			1330 => "0000011110011100000100",
			1331 => "0000000001010011101101",
			1332 => "0011110111001000001100",
			1333 => "0010011100100000001000",
			1334 => "0000011110011100000100",
			1335 => "0000000001010011101101",
			1336 => "0000000001010011101101",
			1337 => "0000000001010011101101",
			1338 => "0000000001010011101101",
			1339 => "0000000101100100000100",
			1340 => "1111111001010100011001",
			1341 => "0011000100001000010000",
			1342 => "0000101110110100001100",
			1343 => "0010011100100000001000",
			1344 => "0001110111001000000100",
			1345 => "0000000001010100011001",
			1346 => "0000000001010100011001",
			1347 => "0000000001010100011001",
			1348 => "0000000001010100011001",
			1349 => "0000000001010100011001",
			1350 => "0010000011011100000100",
			1351 => "0000000001010101000101",
			1352 => "0011101001101000000100",
			1353 => "0000000001010101000101",
			1354 => "0010001100110000000100",
			1355 => "0000000001010101000101",
			1356 => "0011001101010100001000",
			1357 => "0011110111001000000100",
			1358 => "0000000001010101000101",
			1359 => "0000000001010101000101",
			1360 => "0000000001010101000101",
			1361 => "0011111010111000010100",
			1362 => "0010011100100000010000",
			1363 => "0011001101010100001100",
			1364 => "0001010100011000000100",
			1365 => "0000000001010101110001",
			1366 => "0000011110011100000100",
			1367 => "0000000001010101110001",
			1368 => "0000000001010101110001",
			1369 => "0000000001010101110001",
			1370 => "0000000001010101110001",
			1371 => "0000000001010101110001",
			1372 => "0010011100100000011000",
			1373 => "0000101010001000001000",
			1374 => "0001011110110000000100",
			1375 => "0000000001010110100101",
			1376 => "0000000001010110100101",
			1377 => "0011110001111100000100",
			1378 => "0000000001010110100101",
			1379 => "0011111010111000001000",
			1380 => "0001111110110000000100",
			1381 => "0000000001010110100101",
			1382 => "0000000001010110100101",
			1383 => "0000000001010110100101",
			1384 => "1111111001010110100101",
			1385 => "0000000110100000001100",
			1386 => "0010011100100000001000",
			1387 => "0010001011000100000100",
			1388 => "0000000001010111110001",
			1389 => "0000000001010111110001",
			1390 => "1111111001010111110001",
			1391 => "0011011010011100001100",
			1392 => "0010011100100000001000",
			1393 => "0010111010111000000100",
			1394 => "0000001001010111110001",
			1395 => "0000000001010111110001",
			1396 => "0000000001010111110001",
			1397 => "0001101100011000001000",
			1398 => "0000100010000100000100",
			1399 => "0000001001010111110001",
			1400 => "0000000001010111110001",
			1401 => "0000100011001000000100",
			1402 => "0000001001010111110001",
			1403 => "1111111001010111110001",
			1404 => "0010011100100000011100",
			1405 => "0011101001101000001100",
			1406 => "0000001111010000001000",
			1407 => "0010011100100000000100",
			1408 => "0000000001011000110101",
			1409 => "0000000001011000110101",
			1410 => "0000000001011000110101",
			1411 => "0000101001100000001100",
			1412 => "0011001101010100001000",
			1413 => "0000011110011100000100",
			1414 => "0000001001011000110101",
			1415 => "0000000001011000110101",
			1416 => "0000000001011000110101",
			1417 => "0000000001011000110101",
			1418 => "0010100010111100000100",
			1419 => "1111111001011000110101",
			1420 => "0000000001011000110101",
			1421 => "0010011100100000011000",
			1422 => "0001111110001100000100",
			1423 => "0000000001011001110001",
			1424 => "0000101100010100000100",
			1425 => "0000001001011001110001",
			1426 => "0011010100000100001000",
			1427 => "0000011110011100000100",
			1428 => "0000000001011001110001",
			1429 => "0000000001011001110001",
			1430 => "0011010000011100000100",
			1431 => "0000000001011001110001",
			1432 => "0000000001011001110001",
			1433 => "0010100010111100000100",
			1434 => "1111111001011001110001",
			1435 => "0000000001011001110001",
			1436 => "0000001101000100011000",
			1437 => "0010011100100000010100",
			1438 => "0001100111101000001000",
			1439 => "0011111001110000000100",
			1440 => "0000000001011010111101",
			1441 => "0000001001011010111101",
			1442 => "0000011110011100001000",
			1443 => "0010011100100000000100",
			1444 => "0000000001011010111101",
			1445 => "0000000001011010111101",
			1446 => "1111111001011010111101",
			1447 => "1111111001011010111101",
			1448 => "0000101100010100000100",
			1449 => "0000001001011010111101",
			1450 => "0001101100011000000100",
			1451 => "0000001001011010111101",
			1452 => "0001000011100100000100",
			1453 => "1111111001011010111101",
			1454 => "0000000001011010111101",
			1455 => "0000000101100100000100",
			1456 => "1111111001011011111001",
			1457 => "0000011110011100010100",
			1458 => "0011001101010100010000",
			1459 => "0011110111001000001100",
			1460 => "0000000110100000001000",
			1461 => "0000001110101100000100",
			1462 => "0000000001011011111001",
			1463 => "0000000001011011111001",
			1464 => "0000001001011011111001",
			1465 => "0000000001011011111001",
			1466 => "0000000001011011111001",
			1467 => "0011110000001100000100",
			1468 => "0000000001011011111001",
			1469 => "0000000001011011111001",
			1470 => "0001000010100000000100",
			1471 => "1111111001011100111101",
			1472 => "0000101010001000001100",
			1473 => "0000110001110100000100",
			1474 => "0000000001011100111101",
			1475 => "0010011100100000000100",
			1476 => "0000001001011100111101",
			1477 => "0000000001011100111101",
			1478 => "0010001100101100000100",
			1479 => "0000000001011100111101",
			1480 => "0000011110011100001100",
			1481 => "0011000001111100001000",
			1482 => "0000101110110100000100",
			1483 => "0000001001011100111101",
			1484 => "0000000001011100111101",
			1485 => "0000000001011100111101",
			1486 => "0000000001011100111101",
			1487 => "0000000110100000001100",
			1488 => "0010011100100000001000",
			1489 => "0011110101101100000100",
			1490 => "0000000001011110010001",
			1491 => "0000000001011110010001",
			1492 => "1111111001011110010001",
			1493 => "0011011010011100001000",
			1494 => "0010011100100000000100",
			1495 => "0000001001011110010001",
			1496 => "0000000001011110010001",
			1497 => "0000100011001000000100",
			1498 => "0000001001011110010001",
			1499 => "0001000101101000001100",
			1500 => "0011100111000100000100",
			1501 => "1111111001011110010001",
			1502 => "0011010001011000000100",
			1503 => "0000000001011110010001",
			1504 => "0000000001011110010001",
			1505 => "0000100010000100000100",
			1506 => "0000001001011110010001",
			1507 => "0000000001011110010001",
			1508 => "0000001101000100001100",
			1509 => "0010011100100000001000",
			1510 => "0000111011010100000100",
			1511 => "1111111001011111110101",
			1512 => "0000001001011111110101",
			1513 => "1111111001011111110101",
			1514 => "0000100110010000011100",
			1515 => "0011001010111100010000",
			1516 => "0011110001111100001100",
			1517 => "0011110000001100000100",
			1518 => "0000001001011111110101",
			1519 => "0011011010011100000100",
			1520 => "0000001001011111110101",
			1521 => "0000000001011111110101",
			1522 => "0000010001011111110101",
			1523 => "0000100011001000000100",
			1524 => "0000001001011111110101",
			1525 => "0010111110110000000100",
			1526 => "0000000001011111110101",
			1527 => "0000000001011111110101",
			1528 => "0001110111001000001000",
			1529 => "0010011100100000000100",
			1530 => "0000001001011111110101",
			1531 => "1111111001011111110101",
			1532 => "1111111001011111110101",
			1533 => "0010011100100000100100",
			1534 => "0000101010001000001000",
			1535 => "0001011110110000000100",
			1536 => "0000000001100001000001",
			1537 => "0000001001100001000001",
			1538 => "0011110001111100001100",
			1539 => "0001101100011000000100",
			1540 => "0000000001100001000001",
			1541 => "0010100010111100000100",
			1542 => "0000000001100001000001",
			1543 => "0000000001100001000001",
			1544 => "0010101111000100000100",
			1545 => "0000000001100001000001",
			1546 => "0011111010111000001000",
			1547 => "0001111110110000000100",
			1548 => "0000000001100001000001",
			1549 => "0000000001100001000001",
			1550 => "0000000001100001000001",
			1551 => "1111111001100001000001",
			1552 => "0000001110101000011000",
			1553 => "0000011110011100001100",
			1554 => "0000001001010100000100",
			1555 => "1111111001100010101101",
			1556 => "0010101101010000000100",
			1557 => "0000011001100010101101",
			1558 => "1111111001100010101101",
			1559 => "0010100010011000000100",
			1560 => "1111111001100010101101",
			1561 => "0010001100110000000100",
			1562 => "1111111001100010101101",
			1563 => "0000001001100010101101",
			1564 => "0000101110110100011100",
			1565 => "0011001101010100010100",
			1566 => "0011100110001000010000",
			1567 => "0000110011111100001100",
			1568 => "0011111010111100001000",
			1569 => "0011110100001000000100",
			1570 => "0000010001100010101101",
			1571 => "0000001001100010101101",
			1572 => "0000011001100010101101",
			1573 => "0000000001100010101101",
			1574 => "0000011001100010101101",
			1575 => "0000100010000000000100",
			1576 => "0000001001100010101101",
			1577 => "1111111001100010101101",
			1578 => "1111111001100010101101",
			1579 => "0000001101000100001100",
			1580 => "0010011100100000001000",
			1581 => "0000111011010100000100",
			1582 => "1111111001100100100011",
			1583 => "0000001001100100100011",
			1584 => "1111111001100100100011",
			1585 => "0011110111001000101100",
			1586 => "0011001010111100011100",
			1587 => "0000011110011100010000",
			1588 => "0011100110001000001100",
			1589 => "0000110010011000000100",
			1590 => "0000001001100100100011",
			1591 => "0000110010111100000100",
			1592 => "0000000001100100100011",
			1593 => "0000000001100100100011",
			1594 => "0000001001100100100011",
			1595 => "0000110010011000000100",
			1596 => "0000001001100100100011",
			1597 => "0001000101111100000100",
			1598 => "0000000001100100100011",
			1599 => "1111111001100100100011",
			1600 => "0001101010011000000100",
			1601 => "0000001001100100100011",
			1602 => "0001101101011000001000",
			1603 => "0010111010111000000100",
			1604 => "0000000001100100100011",
			1605 => "1111111001100100100011",
			1606 => "0000000001100100100011",
			1607 => "1111111001100100100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(530, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1062, initial_addr_3'length));
	end generate gen_rom_0;

	gen_rom_1: if SELECT_ROM = 1 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000000000000001110101",
			29 => "0000000000000001111001",
			30 => "0000000000000001111101",
			31 => "0000000000000010000001",
			32 => "0000000000000010000101",
			33 => "0000000000000010001001",
			34 => "0000000000000010001101",
			35 => "0000000000000010010001",
			36 => "0000000000000010010101",
			37 => "0000000000000010011001",
			38 => "0001110001111100000100",
			39 => "0000000000000010100101",
			40 => "0000000000000010100101",
			41 => "0001000010010000000100",
			42 => "0000000000000010110001",
			43 => "0000000000000010110001",
			44 => "0000010110000000000100",
			45 => "0000000000000010111101",
			46 => "0000000000000010111101",
			47 => "0010011110100000000100",
			48 => "0000000000000011001001",
			49 => "0000000000000011001001",
			50 => "0010010000011000000100",
			51 => "0000000000000011010101",
			52 => "0000000000000011010101",
			53 => "0001110001111100000100",
			54 => "0000000000000011100001",
			55 => "0000000000000011100001",
			56 => "0001010110100100001000",
			57 => "0001001111111000000100",
			58 => "0000000000000011110101",
			59 => "0000000000000011110101",
			60 => "0000000000000011110101",
			61 => "0000010000011000001000",
			62 => "0000101010001000000100",
			63 => "0000000000000100001001",
			64 => "0000000000000100001001",
			65 => "0000000000000100001001",
			66 => "0001110111001000001000",
			67 => "0000101100010000000100",
			68 => "0000000000000100011101",
			69 => "0000000000000100011101",
			70 => "0000000000000100011101",
			71 => "0010111110001100001000",
			72 => "0011101001101000000100",
			73 => "0000000000000100111001",
			74 => "0000000000000100111001",
			75 => "0001101101011000000100",
			76 => "0000000000000100111001",
			77 => "0000000000000100111001",
			78 => "0010011110100000001000",
			79 => "0000000111100000000100",
			80 => "0000000000000101010101",
			81 => "0000000000000101010101",
			82 => "0001000101001100000100",
			83 => "0000000000000101010101",
			84 => "0000000000000101010101",
			85 => "0010111110001100000100",
			86 => "0000000000000101110001",
			87 => "0001101101011000001000",
			88 => "0001101100011000000100",
			89 => "0000000000000101110001",
			90 => "0000000000000101110001",
			91 => "0000000000000101110001",
			92 => "0001110001111100000100",
			93 => "0000000000000110001101",
			94 => "0000101010001000000100",
			95 => "0000000000000110001101",
			96 => "0000101100111000000100",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0011011010011100001100",
			100 => "0011000100001000001000",
			101 => "0010111010111000000100",
			102 => "0000000000000110101001",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0001111110001100001000",
			107 => "0001001111111000000100",
			108 => "0000000000000111001101",
			109 => "0000000000000111001101",
			110 => "0001101101011000001000",
			111 => "0001101100011000000100",
			112 => "0000000000000111001101",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0001000010010000000100",
			116 => "1111111000000111110001",
			117 => "0011111010111000000100",
			118 => "0000000000000111110001",
			119 => "0011001001110000000100",
			120 => "0000000000000111110001",
			121 => "0000010010001100000100",
			122 => "0000000000000111110001",
			123 => "0000000000000111110001",
			124 => "0000100011001000000100",
			125 => "0000000000001000010101",
			126 => "0000010110000000001100",
			127 => "0010011100100000000100",
			128 => "0000000000001000010101",
			129 => "0011100001110000000100",
			130 => "0000000000001000010101",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0001110001111100000100",
			134 => "0000000000001000111001",
			135 => "0000011001111000001100",
			136 => "0010011100100000000100",
			137 => "0000000000001000111001",
			138 => "0011010001101000000100",
			139 => "0000000000001000111001",
			140 => "0000000000001000111001",
			141 => "0000000000001000111001",
			142 => "0001111110001100001000",
			143 => "0001000000100100000100",
			144 => "1111111000001001100101",
			145 => "0000000000001001100101",
			146 => "0000010010001100001100",
			147 => "0011110100001000000100",
			148 => "0000000000001001100101",
			149 => "0010001101111000000100",
			150 => "0000000000001001100101",
			151 => "0000000000001001100101",
			152 => "0000000000001001100101",
			153 => "0000010110000000010100",
			154 => "0011111101010100001000",
			155 => "0001101100011000000100",
			156 => "0000000000001010010001",
			157 => "0000000000001010010001",
			158 => "0011000011011100000100",
			159 => "0000000000001010010001",
			160 => "0000011110011100000100",
			161 => "0000000000001010010001",
			162 => "0000000000001010010001",
			163 => "1111111000001010010001",
			164 => "0001000101001100000100",
			165 => "1111111000001010111101",
			166 => "0001101100011000000100",
			167 => "0000000000001010111101",
			168 => "0000001111010000001100",
			169 => "0011110100010000001000",
			170 => "0011111101111000000100",
			171 => "0000000000001010111101",
			172 => "0000000000001010111101",
			173 => "0000000000001010111101",
			174 => "0000000000001010111101",
			175 => "0000010110000000011000",
			176 => "0011111101010100001000",
			177 => "0001101100011000000100",
			178 => "0000000000001011110001",
			179 => "0000000000001011110001",
			180 => "0000100101110000000100",
			181 => "0000000000001011110001",
			182 => "0000111111000100000100",
			183 => "0000000000001011110001",
			184 => "0000001011000100000100",
			185 => "0000000000001011110001",
			186 => "0000000000001011110001",
			187 => "1111111000001011110001",
			188 => "0010011100110100011100",
			189 => "0011010110100100001100",
			190 => "0000110011111100001000",
			191 => "0010111010111100000100",
			192 => "0000000000001100101101",
			193 => "0000000000001100101101",
			194 => "0000000000001100101101",
			195 => "0000101010001000000100",
			196 => "0000000000001100101101",
			197 => "0001000101101000001000",
			198 => "0010011100100000000100",
			199 => "0000000000001100101101",
			200 => "0000001000001100101101",
			201 => "0000000000001100101101",
			202 => "1111111000001100101101",
			203 => "0000010110000000011100",
			204 => "0011000100001000010000",
			205 => "0000111100110000001100",
			206 => "0001110111001000001000",
			207 => "0010111110110000000100",
			208 => "0000000000001101101001",
			209 => "0000000000001101101001",
			210 => "0000000000001101101001",
			211 => "0000000000001101101001",
			212 => "0000100011001000000100",
			213 => "0000000000001101101001",
			214 => "0001000011100100000100",
			215 => "0000000000001101101001",
			216 => "0000000000001101101001",
			217 => "1111111000001101101001",
			218 => "0001001111111100011000",
			219 => "0001000100100100001100",
			220 => "0010011100110100001000",
			221 => "0010010110000000000100",
			222 => "1111111000001111001101",
			223 => "1111111000001111001101",
			224 => "1111111000001111001101",
			225 => "0001011000011000000100",
			226 => "1111111000001111001101",
			227 => "0000100101100000000100",
			228 => "0000010000001111001101",
			229 => "1111111000001111001101",
			230 => "0011110000001100001100",
			231 => "0010011100100000000100",
			232 => "1111111000001111001101",
			233 => "0011001110001100000100",
			234 => "1111111000001111001101",
			235 => "0000010000001111001101",
			236 => "0010011100100000001000",
			237 => "0000001001010000000100",
			238 => "0000000000001111001101",
			239 => "1111111000001111001101",
			240 => "0000110010011000000100",
			241 => "0000001000001111001101",
			242 => "0000010000001111001101",
			243 => "0001000101001100000100",
			244 => "1111111000010000000001",
			245 => "0000101010001000000100",
			246 => "0000000000010000000001",
			247 => "0001000101101000010000",
			248 => "0011111001010100001100",
			249 => "0010011100100000000100",
			250 => "0000000000010000000001",
			251 => "0001011010111000000100",
			252 => "0000000000010000000001",
			253 => "0000001000010000000001",
			254 => "0000000000010000000001",
			255 => "0000000000010000000001",
			256 => "0001000010010000000100",
			257 => "1111111000010001000101",
			258 => "0011000100001000001100",
			259 => "0000001011000100000100",
			260 => "0000000000010001000101",
			261 => "0001100100110100000100",
			262 => "0000000000010001000101",
			263 => "0000000000010001000101",
			264 => "0001101101011000010000",
			265 => "0000000101001000001100",
			266 => "0011110000001100000100",
			267 => "0000000000010001000101",
			268 => "0000101000101000000100",
			269 => "0000001000010001000101",
			270 => "0000000000010001000101",
			271 => "0000000000010001000101",
			272 => "0000000000010001000101",
			273 => "0001001111111100011000",
			274 => "0001000010010000000100",
			275 => "1111111000010010101001",
			276 => "0010101100000100001100",
			277 => "0011000110000100000100",
			278 => "1111111000010010101001",
			279 => "0011111111010000000100",
			280 => "0000001000010010101001",
			281 => "0000000000010010101001",
			282 => "0001001101100100000100",
			283 => "1111111000010010101001",
			284 => "0000000000010010101001",
			285 => "0000000111100000001100",
			286 => "0000111111000100000100",
			287 => "0000000000010010101001",
			288 => "0011110000001100000100",
			289 => "0000000000010010101001",
			290 => "0000001000010010101001",
			291 => "0001101100011000000100",
			292 => "1111111000010010101001",
			293 => "0010100010111100001000",
			294 => "0000101100010100000100",
			295 => "0000000000010010101001",
			296 => "0000001000010010101001",
			297 => "1111111000010010101001",
			298 => "0001001111111100011000",
			299 => "0000010000011000010100",
			300 => "0000011110011100001000",
			301 => "0010101100000100000100",
			302 => "0000000000010100010101",
			303 => "1111111000010100010101",
			304 => "0010101001101000000100",
			305 => "0000000000010100010101",
			306 => "0000011110011100000100",
			307 => "0000000000010100010101",
			308 => "0000000000010100010101",
			309 => "1111111000010100010101",
			310 => "0000100011001000010000",
			311 => "0000001101000100001100",
			312 => "0010100001110100001000",
			313 => "0010100111000100000100",
			314 => "0000000000010100010101",
			315 => "0000000000010100010101",
			316 => "0000000000010100010101",
			317 => "1111111000010100010101",
			318 => "0000111111000100000100",
			319 => "0000000000010100010101",
			320 => "0001000101101000000100",
			321 => "0000001000010100010101",
			322 => "0011111010111100000100",
			323 => "0000000000010100010101",
			324 => "0000000000010100010101",
			325 => "0010010000011000101000",
			326 => "0000101010001000001100",
			327 => "0010011100100000001000",
			328 => "0000011110011100000100",
			329 => "1111111000010101111001",
			330 => "0000000000010101111001",
			331 => "0000000000010101111001",
			332 => "0000011110011100010100",
			333 => "0001101100011000001000",
			334 => "0000001100100100000100",
			335 => "0000000000010101111001",
			336 => "1111111000010101111001",
			337 => "0001110001111100000100",
			338 => "0000000000010101111001",
			339 => "0000001111010000000100",
			340 => "0000001000010101111001",
			341 => "0000000000010101111001",
			342 => "0001011010111000000100",
			343 => "0000000000010101111001",
			344 => "0000001000010101111001",
			345 => "0000000110110100001000",
			346 => "0000011100100000000100",
			347 => "0000000000010101111001",
			348 => "1111111000010101111001",
			349 => "0000000000010101111001",
			350 => "0001000010010000000100",
			351 => "1111111000010111000101",
			352 => "0001111110001100001000",
			353 => "0001001101001100000100",
			354 => "1111111000010111000101",
			355 => "0000000000010111000101",
			356 => "0001101101011000010100",
			357 => "0000001100100100001000",
			358 => "0000100101110000000100",
			359 => "0000000000010111000101",
			360 => "0000001000010111000101",
			361 => "0001101100011000000100",
			362 => "1111111000010111000101",
			363 => "0000101100010100000100",
			364 => "0000000000010111000101",
			365 => "0000001000010111000101",
			366 => "0001001111111000000100",
			367 => "0000000000010111000101",
			368 => "0000000000010111000101",
			369 => "0001000010010000000100",
			370 => "1111111000011000001001",
			371 => "0011010011100000000100",
			372 => "0000000000011000001001",
			373 => "0010011100100000010100",
			374 => "0001101100011000001000",
			375 => "0000000010110100000100",
			376 => "0000000000011000001001",
			377 => "1111111000011000001001",
			378 => "0000101010001000000100",
			379 => "0000000000011000001001",
			380 => "0000000010011100000100",
			381 => "0000000000011000001001",
			382 => "0000000000011000001001",
			383 => "0010010111100100000100",
			384 => "0000001000011000001001",
			385 => "0000000000011000001001",
			386 => "0001001111111100010000",
			387 => "0000010000011000001100",
			388 => "0001010100011000000100",
			389 => "1111111000011001011101",
			390 => "0000001001001000000100",
			391 => "0000010000011001011101",
			392 => "0000001000011001011101",
			393 => "1111111000011001011101",
			394 => "0000111111000100000100",
			395 => "1111111000011001011101",
			396 => "0010100010111100010100",
			397 => "0010011100100000000100",
			398 => "1111111000011001011101",
			399 => "0000100100101000000100",
			400 => "0000000000011001011101",
			401 => "0001000011100100001000",
			402 => "0000011100100000000100",
			403 => "0000001000011001011101",
			404 => "0000001000011001011101",
			405 => "0000000000011001011101",
			406 => "1111111000011001011101",
			407 => "0000001010001100010000",
			408 => "0000010110000000001100",
			409 => "0001010100011000000100",
			410 => "1111111000011011000001",
			411 => "0011101111000100000100",
			412 => "0000001000011011000001",
			413 => "0000001000011011000001",
			414 => "1111111000011011000001",
			415 => "0000111111000100000100",
			416 => "1111111000011011000001",
			417 => "0010011100100000001100",
			418 => "0001101100011000000100",
			419 => "1111111000011011000001",
			420 => "0010100010011000000100",
			421 => "0000001000011011000001",
			422 => "0000000000011011000001",
			423 => "0000000101001000001100",
			424 => "0000011011101000001000",
			425 => "0000100111111100000100",
			426 => "0000000000011011000001",
			427 => "0000001000011011000001",
			428 => "0000000000011011000001",
			429 => "0001101010011000000100",
			430 => "1111111000011011000001",
			431 => "0000001000011011000001",
			432 => "0010010000011000100100",
			433 => "0011110111001000011100",
			434 => "0001101100011000001000",
			435 => "0010011100100000000100",
			436 => "0000000000011100100101",
			437 => "0000000000011100100101",
			438 => "0001101101011000010000",
			439 => "0000001111010000001100",
			440 => "0000101010001000000100",
			441 => "0000000000011100100101",
			442 => "0000110000111000000100",
			443 => "0000000000011100100101",
			444 => "0000000000011100100101",
			445 => "0000000000011100100101",
			446 => "0000000000011100100101",
			447 => "0001011010111000000100",
			448 => "0000000000011100100101",
			449 => "0000001000011100100101",
			450 => "0001101110010100000100",
			451 => "0000000000011100100101",
			452 => "0010001000111000001000",
			453 => "0000011100100000000100",
			454 => "0000000000011100100101",
			455 => "1111111000011100100101",
			456 => "0000000000011100100101",
			457 => "0000011100100000101000",
			458 => "0011111010111000100000",
			459 => "0001101100011000001100",
			460 => "0011110111001000001000",
			461 => "0011000001111100000100",
			462 => "0000000000011110001001",
			463 => "0000000000011110001001",
			464 => "0000000000011110001001",
			465 => "0001101101011000010000",
			466 => "0000101010001000000100",
			467 => "0000000000011110001001",
			468 => "0001000011100100001000",
			469 => "0001010100000100000100",
			470 => "0000000000011110001001",
			471 => "0000000000011110001001",
			472 => "0000000000011110001001",
			473 => "0000000000011110001001",
			474 => "0001011010111000000100",
			475 => "0000000000011110001001",
			476 => "0000000000011110001001",
			477 => "0001001101001100001000",
			478 => "0001101110010100000100",
			479 => "0000000000011110001001",
			480 => "1111111000011110001001",
			481 => "0000000000011110001001",
			482 => "0001000010010000000100",
			483 => "1111111000011111001101",
			484 => "0011010100011000000100",
			485 => "1111111000011111001101",
			486 => "0001101001100100011000",
			487 => "0000001100100100001100",
			488 => "0000100101110000000100",
			489 => "0000000000011111001101",
			490 => "0000010010001100000100",
			491 => "0000001000011111001101",
			492 => "0000000000011111001101",
			493 => "0001101100011000000100",
			494 => "1111111000011111001101",
			495 => "0000101100010100000100",
			496 => "0000000000011111001101",
			497 => "0000001000011111001101",
			498 => "1111111000011111001101",
			499 => "0001001111111100010100",
			500 => "0001000010010000000100",
			501 => "1111111000100000110001",
			502 => "0010101100000100001100",
			503 => "0011000110000100000100",
			504 => "1111111000100000110001",
			505 => "0011101010111000000100",
			506 => "0000001000100000110001",
			507 => "0000000000100000110001",
			508 => "1111111000100000110001",
			509 => "0000111111000100000100",
			510 => "1111111000100000110001",
			511 => "0001101011001100011000",
			512 => "0010011100100000010000",
			513 => "0001101100011000001000",
			514 => "0001101100011000000100",
			515 => "1111111000100000110001",
			516 => "0000000000100000110001",
			517 => "0010100010111100000100",
			518 => "0000001000100000110001",
			519 => "0000000000100000110001",
			520 => "0010001101111000000100",
			521 => "0000001000100000110001",
			522 => "0000000000100000110001",
			523 => "0000000000100000110001",
			524 => "0000001010001100001100",
			525 => "0010011110100000001000",
			526 => "0001111110001100000100",
			527 => "1111111000100010011101",
			528 => "0000001000100010011101",
			529 => "1111111000100010011101",
			530 => "0000110010011000001100",
			531 => "0000001100100100001000",
			532 => "0000111111000100000100",
			533 => "0000000000100010011101",
			534 => "0000001000100010011101",
			535 => "1111111000100010011101",
			536 => "0001101000010000011100",
			537 => "0010011100100000001000",
			538 => "0010100010011000000100",
			539 => "0000000000100010011101",
			540 => "0000000000100010011101",
			541 => "0000101010001000001000",
			542 => "0000011110011100000100",
			543 => "0000000000100010011101",
			544 => "0000000000100010011101",
			545 => "0000000111100000000100",
			546 => "0000001000100010011101",
			547 => "0010011100100000000100",
			548 => "0000000000100010011101",
			549 => "0000001000100010011101",
			550 => "1111111000100010011101",
			551 => "0001001111111100100000",
			552 => "0001000100100100010100",
			553 => "0000010000011000010000",
			554 => "0010011110100000001100",
			555 => "0010010000011000000100",
			556 => "1111111000100100010001",
			557 => "0010010000011000000100",
			558 => "0000000000100100010001",
			559 => "1111111000100100010001",
			560 => "0000000000100100010001",
			561 => "1111111000100100010001",
			562 => "0001011000011000000100",
			563 => "1111111000100100010001",
			564 => "0000011011101000000100",
			565 => "0000001000100100010001",
			566 => "1111111000100100010001",
			567 => "0000111111000100000100",
			568 => "1111111000100100010001",
			569 => "0000001111010000010100",
			570 => "0010011100100000000100",
			571 => "0000000000100100010001",
			572 => "0011110000001100000100",
			573 => "0000001000100100010001",
			574 => "0001111110001100000100",
			575 => "0000010000100100010001",
			576 => "0011110100001000000100",
			577 => "0000010000100100010001",
			578 => "0000001000100100010001",
			579 => "1111111000100100010001",
			580 => "0001001111111100010100",
			581 => "0010011110100000010000",
			582 => "0011101000110000001000",
			583 => "0011100111000100000100",
			584 => "1111111000100110001101",
			585 => "0000000000100110001101",
			586 => "0000001011000100000100",
			587 => "0000000000100110001101",
			588 => "0000001000100110001101",
			589 => "1111111000100110001101",
			590 => "0000110010011000001100",
			591 => "0000001100100100001000",
			592 => "0000111111000100000100",
			593 => "0000000000100110001101",
			594 => "0000001000100110001101",
			595 => "1111111000100110001101",
			596 => "0000011100100000011100",
			597 => "0010011100100000001000",
			598 => "0010100010011000000100",
			599 => "0000000000100110001101",
			600 => "0000000000100110001101",
			601 => "0000101010001000001000",
			602 => "0000011110011100000100",
			603 => "0000000000100110001101",
			604 => "0000000000100110001101",
			605 => "0001000011100100001000",
			606 => "0001000001100000000100",
			607 => "0000001000100110001101",
			608 => "0000000000100110001101",
			609 => "0000000000100110001101",
			610 => "0000000000100110001101",
			611 => "0001000010010000000100",
			612 => "1111111000100111111011",
			613 => "0011000100001000011100",
			614 => "0000110011111100001100",
			615 => "0001110111001000001000",
			616 => "0000011110011100000100",
			617 => "0000000000100111111011",
			618 => "1111111000100111111011",
			619 => "0000000000100111111011",
			620 => "0010010000011000001100",
			621 => "0001011010111000000100",
			622 => "0000000000100111111011",
			623 => "0001010100000100000100",
			624 => "0000000000100111111011",
			625 => "0000000000100111111011",
			626 => "0000000000100111111011",
			627 => "0000010010001100010100",
			628 => "0000011110011100010000",
			629 => "0001101100011000000100",
			630 => "0000000000100111111011",
			631 => "0001101101011000001000",
			632 => "0000111111000100000100",
			633 => "0000000000100111111011",
			634 => "0000000000100111111011",
			635 => "0000000000100111111011",
			636 => "0000001000100111111011",
			637 => "0000000000100111111011",
			638 => "0000000000100111111101",
			639 => "0000000000101000000001",
			640 => "0000000000101000000101",
			641 => "0000000000101000001001",
			642 => "0000000000101000001101",
			643 => "0000000000101000010001",
			644 => "0000000000101000010101",
			645 => "0000000000101000011001",
			646 => "0000000000101000011101",
			647 => "0000000000101000100001",
			648 => "0000000000101000100101",
			649 => "0000000000101000101001",
			650 => "0000000000101000101101",
			651 => "0000000000101000110001",
			652 => "0000000000101000110101",
			653 => "0000000000101000111001",
			654 => "0000000000101000111101",
			655 => "0000000000101001000001",
			656 => "0000000000101001000101",
			657 => "0000000000101001001001",
			658 => "0000000000101001001101",
			659 => "0000000000101001010001",
			660 => "0000000000101001010101",
			661 => "0000000000101001011001",
			662 => "0000000000101001011101",
			663 => "0000000000101001100001",
			664 => "0000000000101001100101",
			665 => "0000000000101001101001",
			666 => "0000000000101001101101",
			667 => "0000000000101001110001",
			668 => "0000000000101001110101",
			669 => "0000000000101001111001",
			670 => "0000000000101001111101",
			671 => "0000000000101010000001",
			672 => "0000000000101010000101",
			673 => "0000000000101010001001",
			674 => "0000000000101010001101",
			675 => "0000000000101010010001",
			676 => "0001110001111100000100",
			677 => "0000000000101010011101",
			678 => "0000000000101010011101",
			679 => "0001000010010000000100",
			680 => "0000000000101010101001",
			681 => "0000000000101010101001",
			682 => "0000010110000000000100",
			683 => "0000000000101010110101",
			684 => "0000000000101010110101",
			685 => "0010011110100000000100",
			686 => "0000000000101011000001",
			687 => "0000000000101011000001",
			688 => "0000011100100000000100",
			689 => "0000000000101011001101",
			690 => "0000000000101011001101",
			691 => "0001110001111100000100",
			692 => "0000000000101011011001",
			693 => "0000000000101011011001",
			694 => "0001000010010000000100",
			695 => "0000000000101011101101",
			696 => "0000001100100100000100",
			697 => "0000000000101011101101",
			698 => "0000000000101011101101",
			699 => "0001000010010000000100",
			700 => "0000000000101100000001",
			701 => "0001101001100100000100",
			702 => "0000000000101100000001",
			703 => "0000000000101100000001",
			704 => "0011000100001000001000",
			705 => "0011011010001100000100",
			706 => "0000000000101100010101",
			707 => "0000000000101100010101",
			708 => "0000000000101100010101",
			709 => "0010011110100000001000",
			710 => "0000000111100000000100",
			711 => "0000000000101100110001",
			712 => "0000000000101100110001",
			713 => "0001000101001100000100",
			714 => "0000000000101100110001",
			715 => "0000000000101100110001",
			716 => "0000010110000000001100",
			717 => "0000001100100100001000",
			718 => "0000001011000100000100",
			719 => "0000000000101101001101",
			720 => "0000000000101101001101",
			721 => "0000000000101101001101",
			722 => "0000000000101101001101",
			723 => "0001110001111100001100",
			724 => "0001100001111000000100",
			725 => "0000000000101101101001",
			726 => "0001000000100100000100",
			727 => "0000000000101101101001",
			728 => "0000000000101101101001",
			729 => "0000000000101101101001",
			730 => "0011011010011100001100",
			731 => "0011000100001000001000",
			732 => "0010111010111000000100",
			733 => "0000000000101110000101",
			734 => "0000000000101110000101",
			735 => "0000000000101110000101",
			736 => "0000000000101110000101",
			737 => "0001110111001000001100",
			738 => "0011101001101000000100",
			739 => "0000000000101110100001",
			740 => "0000101111010100000100",
			741 => "0000000000101110100001",
			742 => "0000000000101110100001",
			743 => "0000000000101110100001",
			744 => "0001110001111100001100",
			745 => "0001100001111000000100",
			746 => "0000000000101111001101",
			747 => "0001000000100100000100",
			748 => "0000000000101111001101",
			749 => "0000000000101111001101",
			750 => "0000101010001000000100",
			751 => "0000000000101111001101",
			752 => "0000101000101000000100",
			753 => "0000000000101111001101",
			754 => "0000000000101111001101",
			755 => "0000010110000000010000",
			756 => "0011111101010100000100",
			757 => "0000000000101111110001",
			758 => "0011000011011100000100",
			759 => "0000000000101111110001",
			760 => "0010011100100000000100",
			761 => "0000000000101111110001",
			762 => "0000000000101111110001",
			763 => "0000000000101111110001",
			764 => "0000100011001000000100",
			765 => "0000000000110000010101",
			766 => "0000010110000000001100",
			767 => "0000011110011100000100",
			768 => "0000000000110000010101",
			769 => "0011100001110000000100",
			770 => "0000000000110000010101",
			771 => "0000000000110000010101",
			772 => "0000000000110000010101",
			773 => "0001110111001000010000",
			774 => "0011101001101000000100",
			775 => "0000000000110000111001",
			776 => "0001100101011100000100",
			777 => "0000000000110000111001",
			778 => "0011001101010100000100",
			779 => "0000000000110000111001",
			780 => "0000000000110000111001",
			781 => "0000000000110000111001",
			782 => "0001111110001100001000",
			783 => "0001001101001100000100",
			784 => "1111111000110001100101",
			785 => "0000000000110001100101",
			786 => "0001101101011000001100",
			787 => "0010011100100000000100",
			788 => "0000000000110001100101",
			789 => "0010010111100100000100",
			790 => "0000000000110001100101",
			791 => "0000000000110001100101",
			792 => "0000000000110001100101",
			793 => "0010010000011000010100",
			794 => "0011110000001100000100",
			795 => "0000000000110010011001",
			796 => "0010001101111000001100",
			797 => "0010111000000000001000",
			798 => "0001011010111000000100",
			799 => "0000000000110010011001",
			800 => "0000000000110010011001",
			801 => "0000000000110010011001",
			802 => "0000000000110010011001",
			803 => "0001110111001000000100",
			804 => "1111111000110010011001",
			805 => "0000000000110010011001",
			806 => "0001000101001100000100",
			807 => "1111111000110011000101",
			808 => "0001101100011000000100",
			809 => "0000000000110011000101",
			810 => "0010100010111100001100",
			811 => "0011110100010000001000",
			812 => "0011111101111000000100",
			813 => "0000000000110011000101",
			814 => "0000000000110011000101",
			815 => "0000000000110011000101",
			816 => "0000000000110011000101",
			817 => "0001001101001100001100",
			818 => "0000011100100000001000",
			819 => "0011000000001100000100",
			820 => "0000000000110100001001",
			821 => "0000000000110100001001",
			822 => "1111111000110100001001",
			823 => "0000101110010000001000",
			824 => "0010011100100000000100",
			825 => "1111111000110100001001",
			826 => "0000000000110100001001",
			827 => "0000111111000100000100",
			828 => "0000000000110100001001",
			829 => "0001000011100100001000",
			830 => "0010011100100000000100",
			831 => "0000000000110100001001",
			832 => "0000001000110100001001",
			833 => "0000000000110100001001",
			834 => "0001110001111100001000",
			835 => "0001000000100100000100",
			836 => "1111111000110101000101",
			837 => "0000000000110101000101",
			838 => "0000010010001100010100",
			839 => "0010011100100000010000",
			840 => "0011101001101000001000",
			841 => "0000111111000100000100",
			842 => "0000000000110101000101",
			843 => "0000000000110101000101",
			844 => "0000110010111100000100",
			845 => "0000000000110101000101",
			846 => "0000000000110101000101",
			847 => "0000000000110101000101",
			848 => "0000000000110101000101",
			849 => "0011001100110000000100",
			850 => "1111111000110110000001",
			851 => "0001101101011000010000",
			852 => "0011110000001100000100",
			853 => "0000000000110110000001",
			854 => "0001000001100000001000",
			855 => "0000011100110100000100",
			856 => "0000000000110110000001",
			857 => "0000000000110110000001",
			858 => "0000000000110110000001",
			859 => "0001010011100000000100",
			860 => "0000000000110110000001",
			861 => "0001000000100100000100",
			862 => "0000000000110110000001",
			863 => "0000000000110110000001",
			864 => "0001001111111100001100",
			865 => "0000010110000000001000",
			866 => "0001010100011000000100",
			867 => "1111111000110111001101",
			868 => "0000001000110111001101",
			869 => "1111111000110111001101",
			870 => "0000111111000100000100",
			871 => "1111111000110111001101",
			872 => "0010011100100000001100",
			873 => "0001101100011000000100",
			874 => "1111111000110111001101",
			875 => "0010100010011000000100",
			876 => "0000001000110111001101",
			877 => "0000000000110111001101",
			878 => "0001000011100100001000",
			879 => "0000001001010000000100",
			880 => "0000001000110111001101",
			881 => "0000000000110111001101",
			882 => "0000000000110111001101",
			883 => "0001000010010000000100",
			884 => "1111111000111000010001",
			885 => "0011000100001000010000",
			886 => "0000001011000100000100",
			887 => "0000000000111000010001",
			888 => "0001000000100100001000",
			889 => "0001110111001000000100",
			890 => "0000000000111000010001",
			891 => "0000000000111000010001",
			892 => "0000000000111000010001",
			893 => "0000110111110000001100",
			894 => "0000100011001000000100",
			895 => "0000000000111000010001",
			896 => "0001000011100100000100",
			897 => "0000001000111000010001",
			898 => "0000000000111000010001",
			899 => "0000000000111000010001",
			900 => "0001001111111100010100",
			901 => "0000010000011000001000",
			902 => "0001011000011000000100",
			903 => "1111111000111001101101",
			904 => "0000010000111001101101",
			905 => "0000010110000000001000",
			906 => "0000010110000000000100",
			907 => "1111111000111001101101",
			908 => "1111111000111001101101",
			909 => "1111111000111001101101",
			910 => "0011111101111000000100",
			911 => "1111111000111001101101",
			912 => "0001000011100100010000",
			913 => "0001010100011000000100",
			914 => "0000000000111001101101",
			915 => "0010011100100000000100",
			916 => "0000000000111001101101",
			917 => "0000001111010000000100",
			918 => "0000001000111001101101",
			919 => "0000000000111001101101",
			920 => "0001101100011000000100",
			921 => "1111111000111001101101",
			922 => "0000000000111001101101",
			923 => "0001001101001100010000",
			924 => "0001001011100100000100",
			925 => "1111111000111011001001",
			926 => "0001110001111100000100",
			927 => "1111111000111011001001",
			928 => "0010010111100100000100",
			929 => "0000001000111011001001",
			930 => "0000000000111011001001",
			931 => "0000101110010000001000",
			932 => "0010011100100000000100",
			933 => "1111111000111011001001",
			934 => "0000000000111011001001",
			935 => "0000011110011100010100",
			936 => "0001101100011000001000",
			937 => "0010101101010000000100",
			938 => "0000000000111011001001",
			939 => "1111111000111011001001",
			940 => "0001110001111100000100",
			941 => "0000000000111011001001",
			942 => "0000001111010000000100",
			943 => "0000001000111011001001",
			944 => "0000000000111011001001",
			945 => "0000001000111011001001",
			946 => "0010010000011000100100",
			947 => "0011110111001000011100",
			948 => "0001101100011000001100",
			949 => "0000011110011100001000",
			950 => "0010011100100000000100",
			951 => "1111111000111100110101",
			952 => "0000000000111100110101",
			953 => "0000000000111100110101",
			954 => "0010100010111100001100",
			955 => "0000101010001000000100",
			956 => "0000000000111100110101",
			957 => "0001010100000100000100",
			958 => "0000000000111100110101",
			959 => "0000000000111100110101",
			960 => "0000000000111100110101",
			961 => "0001011010111000000100",
			962 => "0000000000111100110101",
			963 => "0000001000111100110101",
			964 => "0000000110000100001000",
			965 => "0000010000011000000100",
			966 => "0000000000111100110101",
			967 => "1111111000111100110101",
			968 => "0011000100001000000100",
			969 => "0000000000111100110101",
			970 => "0000010010001100000100",
			971 => "0000000000111100110101",
			972 => "0000000000111100110101",
			973 => "0010010000011000100100",
			974 => "0011110111001000011100",
			975 => "0001101100011000001000",
			976 => "0010011100100000000100",
			977 => "0000000000111110011001",
			978 => "0000000000111110011001",
			979 => "0001101101011000001100",
			980 => "0000001111010000001000",
			981 => "0000101010001000000100",
			982 => "0000000000111110011001",
			983 => "0000000000111110011001",
			984 => "0000000000111110011001",
			985 => "0000011110011100000100",
			986 => "0000000000111110011001",
			987 => "0000000000111110011001",
			988 => "0001011010111000000100",
			989 => "0000000000111110011001",
			990 => "0000001000111110011001",
			991 => "0001101110010100000100",
			992 => "0000000000111110011001",
			993 => "0010001000111000001000",
			994 => "0000011100100000000100",
			995 => "0000000000111110011001",
			996 => "1111111000111110011001",
			997 => "0000000000111110011001",
			998 => "0001001111101100000100",
			999 => "1111111000111111100101",
			1000 => "0011000100001000010000",
			1001 => "0000110011111100001100",
			1002 => "0000011110011100000100",
			1003 => "0000000000111111100101",
			1004 => "0001110111001000000100",
			1005 => "0000000000111111100101",
			1006 => "0000000000111111100101",
			1007 => "0000000000111111100101",
			1008 => "0000101010001000000100",
			1009 => "0000000000111111100101",
			1010 => "0000011110011100000100",
			1011 => "0000000000111111100101",
			1012 => "0000010010001100001000",
			1013 => "0000000101001000000100",
			1014 => "0000000000111111100101",
			1015 => "0000000000111111100101",
			1016 => "0000000000111111100101",
			1017 => "0001001101001100010000",
			1018 => "0001000101001100000100",
			1019 => "1111111001000001000001",
			1020 => "0001110100001000000100",
			1021 => "1111111001000001000001",
			1022 => "0000011001111000000100",
			1023 => "0000000001000001000001",
			1024 => "0000000001000001000001",
			1025 => "0011110000001100001000",
			1026 => "0010011100100000000100",
			1027 => "0000000001000001000001",
			1028 => "0000000001000001000001",
			1029 => "0001000011100100010100",
			1030 => "0010111100101000000100",
			1031 => "0000000001000001000001",
			1032 => "0010111000000000001100",
			1033 => "0010100010111100001000",
			1034 => "0010011100100000000100",
			1035 => "0000000001000001000001",
			1036 => "0000001001000001000001",
			1037 => "0000000001000001000001",
			1038 => "0000000001000001000001",
			1039 => "0000000001000001000001",
			1040 => "0001001111111100100100",
			1041 => "0001000100100100011000",
			1042 => "0000010000011000010100",
			1043 => "0010011110100000001100",
			1044 => "0010010000011000000100",
			1045 => "1111111001000010101101",
			1046 => "0010010000011000000100",
			1047 => "0000000001000010101101",
			1048 => "1111111001000010101101",
			1049 => "0000000111111000000100",
			1050 => "1111111001000010101101",
			1051 => "0000001001000010101101",
			1052 => "1111111001000010101101",
			1053 => "0001011000011000000100",
			1054 => "1111111001000010101101",
			1055 => "0000011011101000000100",
			1056 => "0000001001000010101101",
			1057 => "1111111001000010101101",
			1058 => "0011111101111000000100",
			1059 => "1111111001000010101101",
			1060 => "0000001111010000001100",
			1061 => "0000111111000100000100",
			1062 => "1111111001000010101101",
			1063 => "0000011110011100000100",
			1064 => "0000001001000010101101",
			1065 => "0000001001000010101101",
			1066 => "1111111001000010101101",
			1067 => "0001001111111100010100",
			1068 => "0001000010010000000100",
			1069 => "1111111001000100010001",
			1070 => "0010101100000100001100",
			1071 => "0011000110000100000100",
			1072 => "1111111001000100010001",
			1073 => "0011101010111000000100",
			1074 => "0000010001000100010001",
			1075 => "1111111001000100010001",
			1076 => "1111111001000100010001",
			1077 => "0000111111000100000100",
			1078 => "1111111001000100010001",
			1079 => "0010011100100000010000",
			1080 => "0001101100011000000100",
			1081 => "1111111001000100010001",
			1082 => "0000100011001000001000",
			1083 => "0001001011010000000100",
			1084 => "0000000001000100010001",
			1085 => "0000000001000100010001",
			1086 => "0000001001000100010001",
			1087 => "0000101000101000001000",
			1088 => "0010001101111000000100",
			1089 => "0000001001000100010001",
			1090 => "0000000001000100010001",
			1091 => "0000000001000100010001",
			1092 => "0001001111111100010000",
			1093 => "0000010000011000001100",
			1094 => "0001010100011000000100",
			1095 => "1111111001000101101101",
			1096 => "0001001111110100000100",
			1097 => "0000010001000101101101",
			1098 => "0000001001000101101101",
			1099 => "1111111001000101101101",
			1100 => "0000111111000100000100",
			1101 => "1111111001000101101101",
			1102 => "0010011100100000001000",
			1103 => "0001101100011000000100",
			1104 => "1111111001000101101101",
			1105 => "0000001001000101101101",
			1106 => "0001000011100100010000",
			1107 => "0010100011111100001100",
			1108 => "0000100100101000000100",
			1109 => "0000000001000101101101",
			1110 => "0010010000011000000100",
			1111 => "0000001001000101101101",
			1112 => "0000001001000101101101",
			1113 => "1111111001000101101101",
			1114 => "0000000001000101101101",
			1115 => "0001000010010000000100",
			1116 => "1111111001000110111001",
			1117 => "0001111110001100001000",
			1118 => "0011010100011000000100",
			1119 => "1111111001000110111001",
			1120 => "0000000001000110111001",
			1121 => "0001101011001100011000",
			1122 => "0000001100100100001100",
			1123 => "0000100101110000000100",
			1124 => "0000000001000110111001",
			1125 => "0000010110101000000100",
			1126 => "0000001001000110111001",
			1127 => "0000000001000110111001",
			1128 => "0001101100011000000100",
			1129 => "1111111001000110111001",
			1130 => "0000101100010100000100",
			1131 => "0000000001000110111001",
			1132 => "0000001001000110111001",
			1133 => "1111111001000110111001",
			1134 => "0001000010010000000100",
			1135 => "1111111001000111111101",
			1136 => "0000100101110000000100",
			1137 => "0000000001000111111101",
			1138 => "0001101101011000010100",
			1139 => "0001000001100000010000",
			1140 => "0001110110000100000100",
			1141 => "0000000001000111111101",
			1142 => "0000011110100000001000",
			1143 => "0011110000001100000100",
			1144 => "0000000001000111111101",
			1145 => "0000001001000111111101",
			1146 => "0000000001000111111101",
			1147 => "0000000001000111111101",
			1148 => "0001001111111000000100",
			1149 => "0000000001000111111101",
			1150 => "0000000001000111111101",
			1151 => "0000000111010000011100",
			1152 => "0000001111011100010000",
			1153 => "0000010000011000001100",
			1154 => "0001010100011000000100",
			1155 => "1111111001001001110001",
			1156 => "0000001011000000000100",
			1157 => "0000101001001001110001",
			1158 => "0000011001001001110001",
			1159 => "1111111001001001110001",
			1160 => "0000110000111000000100",
			1161 => "1111111001001001110001",
			1162 => "0000011101101000000100",
			1163 => "0000011001001001110001",
			1164 => "1111111001001001110001",
			1165 => "0000111111000100000100",
			1166 => "1111111001001001110001",
			1167 => "0010100010111100010100",
			1168 => "0011111101111000000100",
			1169 => "1111111001001001110001",
			1170 => "0000001111010000001100",
			1171 => "0001101001100100001000",
			1172 => "0011011001001000000100",
			1173 => "0000100001001001110001",
			1174 => "0000011001001001110001",
			1175 => "0000000001001001110001",
			1176 => "1111111001001001110001",
			1177 => "0011101001101000000100",
			1178 => "0000000001001001110001",
			1179 => "1111111001001001110001",
			1180 => "0001000010010000000100",
			1181 => "1111111001001011001101",
			1182 => "0000100101110000001000",
			1183 => "0011000001111100000100",
			1184 => "1111111001001011001101",
			1185 => "0000000001001011001101",
			1186 => "0001101101011000011000",
			1187 => "0000001100100100001100",
			1188 => "0001110101101100000100",
			1189 => "0000000001001011001101",
			1190 => "0010010111100100000100",
			1191 => "0000001001001011001101",
			1192 => "0000000001001011001101",
			1193 => "0001101100011000000100",
			1194 => "0000000001001011001101",
			1195 => "0000101100010100000100",
			1196 => "0000000001001011001101",
			1197 => "0000001001001011001101",
			1198 => "0001101001100100000100",
			1199 => "0000000001001011001101",
			1200 => "0001111110001100000100",
			1201 => "0000000001001011001101",
			1202 => "0000000001001011001101",
			1203 => "0001001111111100100100",
			1204 => "0000010000011000100000",
			1205 => "0010010000011000001000",
			1206 => "0010101100000100000100",
			1207 => "0000000001001101011001",
			1208 => "1111111001001101011001",
			1209 => "0010000011111100001100",
			1210 => "0010100110011100001000",
			1211 => "0010101010110000000100",
			1212 => "0000000001001101011001",
			1213 => "0000000001001101011001",
			1214 => "0000000001001101011001",
			1215 => "0010000100010100001000",
			1216 => "0010101001101000000100",
			1217 => "0000000001001101011001",
			1218 => "0000000001001101011001",
			1219 => "0000000001001101011001",
			1220 => "1111111001001101011001",
			1221 => "0000100011001000001100",
			1222 => "0010011100100000000100",
			1223 => "1111111001001101011001",
			1224 => "0010100111000100000100",
			1225 => "0000000001001101011001",
			1226 => "0000000001001101011001",
			1227 => "0001000101101000001100",
			1228 => "0001101101011000001000",
			1229 => "0010011100100000000100",
			1230 => "0000000001001101011001",
			1231 => "0000001001001101011001",
			1232 => "0000000001001101011001",
			1233 => "0001101100011000000100",
			1234 => "0000000001001101011001",
			1235 => "0000100110010000000100",
			1236 => "0000000001001101011001",
			1237 => "0000000001001101011001",
			1238 => "0001001111101100000100",
			1239 => "1111111001001110110101",
			1240 => "0011000100001000010100",
			1241 => "0011100110001000010000",
			1242 => "0011101001101000000100",
			1243 => "0000000001001110110101",
			1244 => "0011011010001100001000",
			1245 => "0001111110110000000100",
			1246 => "0000000001001110110101",
			1247 => "0000000001001110110101",
			1248 => "0000000001001110110101",
			1249 => "0000000001001110110101",
			1250 => "0001101100011000000100",
			1251 => "0000000001001110110101",
			1252 => "0001101101011000010000",
			1253 => "0010011100100000000100",
			1254 => "0000000001001110110101",
			1255 => "0011111101111000000100",
			1256 => "0000000001001110110101",
			1257 => "0011110110110100000100",
			1258 => "0000000001001110110101",
			1259 => "0000000001001110110101",
			1260 => "0000000001001110110101",
			1261 => "0001000010010000000100",
			1262 => "1111111001010000010011",
			1263 => "0000100101110000001000",
			1264 => "0011000001111100000100",
			1265 => "1111111001010000010011",
			1266 => "0000000001010000010011",
			1267 => "0000010110000000100000",
			1268 => "0000011110011100010100",
			1269 => "0000001100100100001000",
			1270 => "0011101001101000000100",
			1271 => "0000000001010000010011",
			1272 => "0000000001010000010011",
			1273 => "0011100110001000001000",
			1274 => "0011011000011000000100",
			1275 => "0000000001010000010011",
			1276 => "0000000001010000010011",
			1277 => "0000000001010000010011",
			1278 => "0001011010111000000100",
			1279 => "0000000001010000010011",
			1280 => "0000000100101000000100",
			1281 => "0000001001010000010011",
			1282 => "0000000001010000010011",
			1283 => "0000000001010000010011",
			1284 => "0000000001010000010101",
			1285 => "0000000001010000011001",
			1286 => "0000000001010000011101",
			1287 => "0000000001010000100001",
			1288 => "0000000001010000100101",
			1289 => "0000000001010000101001",
			1290 => "0000000001010000101101",
			1291 => "0000000001010000110001",
			1292 => "0000000001010000110101",
			1293 => "0000000001010000111001",
			1294 => "0000000001010000111101",
			1295 => "0000000001010001000001",
			1296 => "0000000001010001000101",
			1297 => "0000000001010001001001",
			1298 => "0000000001010001001101",
			1299 => "0000000001010001010001",
			1300 => "0000000001010001010101",
			1301 => "0000000001010001011001",
			1302 => "0000000001010001011101",
			1303 => "0000000001010001100001",
			1304 => "0000000001010001100101",
			1305 => "0000000001010001101001",
			1306 => "0000000001010001101101",
			1307 => "0000000001010001110001",
			1308 => "0000000001010001110101",
			1309 => "0000000001010001111001",
			1310 => "0000000001010001111101",
			1311 => "0000000001010010000001",
			1312 => "0000000001010010000101",
			1313 => "0000000001010010001001",
			1314 => "0000000001010010001101",
			1315 => "0000000001010010010001",
			1316 => "0000000001010010010101",
			1317 => "0000000001010010011001",
			1318 => "0000000001010010011101",
			1319 => "0000000001010010100001",
			1320 => "0000000001010010100101",
			1321 => "0000000001010010101001",
			1322 => "0001000010010000000100",
			1323 => "0000000001010010110101",
			1324 => "0000000001010010110101",
			1325 => "0001110110000100000100",
			1326 => "0000000001010011000001",
			1327 => "0000000001010011000001",
			1328 => "0001110001111100000100",
			1329 => "0000000001010011001101",
			1330 => "0000000001010011001101",
			1331 => "0010011110100000000100",
			1332 => "0000000001010011011001",
			1333 => "0000000001010011011001",
			1334 => "0010010000011000000100",
			1335 => "0000000001010011100101",
			1336 => "0000000001010011100101",
			1337 => "0001110001111100000100",
			1338 => "0000000001010011110001",
			1339 => "0000000001010011110001",
			1340 => "0000010000011000001000",
			1341 => "0000101010001000000100",
			1342 => "0000000001010100000101",
			1343 => "0000000001010100000101",
			1344 => "0000000001010100000101",
			1345 => "0010011110100000000100",
			1346 => "0000000001010100011001",
			1347 => "0001000101001100000100",
			1348 => "0000000001010100011001",
			1349 => "0000000001010100011001",
			1350 => "0010111110001100001000",
			1351 => "0011101001101000000100",
			1352 => "0000000001010100110101",
			1353 => "0000000001010100110101",
			1354 => "0001101101011000000100",
			1355 => "0000000001010100110101",
			1356 => "0000000001010100110101",
			1357 => "0010011110100000001000",
			1358 => "0000000111100000000100",
			1359 => "0000000001010101010001",
			1360 => "0000000001010101010001",
			1361 => "0001000101001100000100",
			1362 => "0000000001010101010001",
			1363 => "0000000001010101010001",
			1364 => "0000010000011000001100",
			1365 => "0001101100011000000100",
			1366 => "0000000001010101101101",
			1367 => "0000101010001000000100",
			1368 => "0000000001010101101101",
			1369 => "0000000001010101101101",
			1370 => "0000000001010101101101",
			1371 => "0001110001111100000100",
			1372 => "0000000001010110001001",
			1373 => "0000101010001000000100",
			1374 => "0000000001010110001001",
			1375 => "0000101100111000000100",
			1376 => "0000000001010110001001",
			1377 => "0000000001010110001001",
			1378 => "0011011010011100001100",
			1379 => "0011000100001000001000",
			1380 => "0010111010111000000100",
			1381 => "0000000001010110100101",
			1382 => "0000000001010110100101",
			1383 => "0000000001010110100101",
			1384 => "0000000001010110100101",
			1385 => "0011000100001000001100",
			1386 => "0011011010001100001000",
			1387 => "0001110111001000000100",
			1388 => "0000000001010111000001",
			1389 => "0000000001010111000001",
			1390 => "0000000001010111000001",
			1391 => "0000000001010111000001",
			1392 => "0001110110000100000100",
			1393 => "1111111001010111100101",
			1394 => "0000011100110100001100",
			1395 => "0011110000001100000100",
			1396 => "0000000001010111100101",
			1397 => "0000001100100100000100",
			1398 => "0000000001010111100101",
			1399 => "0000000001010111100101",
			1400 => "0000000001010111100101",
			1401 => "0000100011001000000100",
			1402 => "0000000001011000001001",
			1403 => "0000010110000000001100",
			1404 => "0010011100100000000100",
			1405 => "0000000001011000001001",
			1406 => "0011100001110000000100",
			1407 => "0000000001011000001001",
			1408 => "0000000001011000001001",
			1409 => "0000000001011000001001",
			1410 => "0001110001111100000100",
			1411 => "0000000001011000101101",
			1412 => "0000011001111000001100",
			1413 => "0010011100100000000100",
			1414 => "0000000001011000101101",
			1415 => "0011010001101000000100",
			1416 => "0000000001011000101101",
			1417 => "0000000001011000101101",
			1418 => "0000000001011000101101",
			1419 => "0011000100001000010000",
			1420 => "0011101100000100000100",
			1421 => "0000000001011001010001",
			1422 => "0011011010001100001000",
			1423 => "0001110111001000000100",
			1424 => "0000000001011001010001",
			1425 => "0000000001011001010001",
			1426 => "0000000001011001010001",
			1427 => "0000000001011001010001",
			1428 => "0001111110001100001000",
			1429 => "0001001111111000000100",
			1430 => "0000000001011001111101",
			1431 => "0000000001011001111101",
			1432 => "0001101101011000001100",
			1433 => "0001101100011000000100",
			1434 => "0000000001011001111101",
			1435 => "0001101101011000000100",
			1436 => "0000000001011001111101",
			1437 => "0000000001011001111101",
			1438 => "0000000001011001111101",
			1439 => "0001111110001100001000",
			1440 => "0001001111111000000100",
			1441 => "0000000001011010110001",
			1442 => "0000000001011010110001",
			1443 => "0001101101011000010000",
			1444 => "0010011100100000000100",
			1445 => "0000000001011010110001",
			1446 => "0000010010001100001000",
			1447 => "0011101100000100000100",
			1448 => "0000000001011010110001",
			1449 => "0000000001011010110001",
			1450 => "0000000001011010110001",
			1451 => "0000000001011010110001",
			1452 => "0001110001111100000100",
			1453 => "0000000001011011011101",
			1454 => "0000011001111000010000",
			1455 => "0000101010001000000100",
			1456 => "0000000001011011011101",
			1457 => "0001000101101000001000",
			1458 => "0010011100100000000100",
			1459 => "0000000001011011011101",
			1460 => "0000000001011011011101",
			1461 => "0000000001011011011101",
			1462 => "0000000001011011011101",
			1463 => "0000010000011000011100",
			1464 => "0011010110100100001100",
			1465 => "0000110011111100001000",
			1466 => "0010111010111100000100",
			1467 => "0000000001011100100001",
			1468 => "0000000001011100100001",
			1469 => "0000000001011100100001",
			1470 => "0000101010001000001000",
			1471 => "0010011100100000000100",
			1472 => "0000000001011100100001",
			1473 => "0000000001011100100001",
			1474 => "0000000001000000000100",
			1475 => "0000000001011100100001",
			1476 => "0000000001011100100001",
			1477 => "0000001010001100000100",
			1478 => "1111111001011100100001",
			1479 => "0000000001011100100001",
			1480 => "0001000010010000000100",
			1481 => "1111111001011101011101",
			1482 => "0011000100001000001100",
			1483 => "0000110011111100001000",
			1484 => "0001111110110000000100",
			1485 => "0000000001011101011101",
			1486 => "0000000001011101011101",
			1487 => "0000000001011101011101",
			1488 => "0000010010001100001100",
			1489 => "0000100011001000000100",
			1490 => "0000000001011101011101",
			1491 => "0001000011100100000100",
			1492 => "0000000001011101011101",
			1493 => "0000000001011101011101",
			1494 => "0000000001011101011101",
			1495 => "0001111110001100001000",
			1496 => "0011000110000100000100",
			1497 => "1111111001011110011001",
			1498 => "0000000001011110011001",
			1499 => "0000010010001100010100",
			1500 => "0000000110100000000100",
			1501 => "0000000001011110011001",
			1502 => "0001101100011000000100",
			1503 => "0000000001011110011001",
			1504 => "0001101011001100001000",
			1505 => "0011001110001100000100",
			1506 => "0000000001011110011001",
			1507 => "0000000001011110011001",
			1508 => "0000000001011110011001",
			1509 => "0000000001011110011001",
			1510 => "0001000010010000000100",
			1511 => "1111111001011111001101",
			1512 => "0001101001100100010100",
			1513 => "0000100101110000000100",
			1514 => "0000000001011111001101",
			1515 => "0000000111100000001100",
			1516 => "0001110110000100000100",
			1517 => "0000000001011111001101",
			1518 => "0000011110100000000100",
			1519 => "0000001001011111001101",
			1520 => "0000000001011111001101",
			1521 => "0000000001011111001101",
			1522 => "0000000001011111001101",
			1523 => "0001001101001100010000",
			1524 => "0001001011100100000100",
			1525 => "1111111001100000101001",
			1526 => "0001110001111100000100",
			1527 => "1111111001100000101001",
			1528 => "0010010111100100000100",
			1529 => "0000001001100000101001",
			1530 => "0000000001100000101001",
			1531 => "0011110111001000011000",
			1532 => "0001101100011000001000",
			1533 => "0010011100100000000100",
			1534 => "1111111001100000101001",
			1535 => "0000000001100000101001",
			1536 => "0001101101011000001000",
			1537 => "0011110000001100000100",
			1538 => "0000000001100000101001",
			1539 => "0000001001100000101001",
			1540 => "0001110111001000000100",
			1541 => "0000000001100000101001",
			1542 => "0000000001100000101001",
			1543 => "0010011100100000000100",
			1544 => "0000000001100000101001",
			1545 => "0000001001100000101001",
			1546 => "0001001111111100011000",
			1547 => "0001000010010000000100",
			1548 => "1111111001100010000101",
			1549 => "0010101100000100001100",
			1550 => "0011000110000100000100",
			1551 => "1111111001100010000101",
			1552 => "0011111111010000000100",
			1553 => "0000001001100010000101",
			1554 => "0000000001100010000101",
			1555 => "0001001101100100000100",
			1556 => "1111111001100010000101",
			1557 => "0000000001100010000101",
			1558 => "0011111101111000000100",
			1559 => "1111111001100010000101",
			1560 => "0000000111100000001000",
			1561 => "0010111110001100000100",
			1562 => "0000000001100010000101",
			1563 => "0000001001100010000101",
			1564 => "0001101100011000000100",
			1565 => "1111111001100010000101",
			1566 => "0010100010111100000100",
			1567 => "0000001001100010000101",
			1568 => "0000000001100010000101",
			1569 => "0001000010100000011100",
			1570 => "0001001111111100010100",
			1571 => "0001000100100100001000",
			1572 => "0000010110000000000100",
			1573 => "1101010001100011111001",
			1574 => "1101010001100011111001",
			1575 => "0001011000011000000100",
			1576 => "1101010001100011111001",
			1577 => "0000011101101000000100",
			1578 => "1110110001100011111001",
			1579 => "1101010001100011111001",
			1580 => "0000100011001000000100",
			1581 => "1101010001100011111001",
			1582 => "1110101001100011111001",
			1583 => "0011110000001100001100",
			1584 => "0000001101000100001000",
			1585 => "0000100101110000000100",
			1586 => "1101010001100011111001",
			1587 => "1110011001100011111001",
			1588 => "1101010001100011111001",
			1589 => "0000001111010000010000",
			1590 => "0011110100001000001000",
			1591 => "0000000111100000000100",
			1592 => "1110101001100011111001",
			1593 => "1101011001100011111001",
			1594 => "0001011001001000000100",
			1595 => "1110001001100011111001",
			1596 => "1110110001100011111001",
			1597 => "1101010001100011111001",
			1598 => "0000001010001100010000",
			1599 => "0001000010010000000100",
			1600 => "1111111001100101011101",
			1601 => "0001111110001100000100",
			1602 => "1111111001100101011101",
			1603 => "0000010010001100000100",
			1604 => "0000001001100101011101",
			1605 => "1111111001100101011101",
			1606 => "0010011100100000010000",
			1607 => "0001101100011000000100",
			1608 => "1111111001100101011101",
			1609 => "0000001111010000001000",
			1610 => "0000111111000100000100",
			1611 => "0000000001100101011101",
			1612 => "0000001001100101011101",
			1613 => "0000000001100101011101",
			1614 => "0010100010111100010000",
			1615 => "0001001111111100000100",
			1616 => "0000000001100101011101",
			1617 => "0000000101001000001000",
			1618 => "0000111111000100000100",
			1619 => "0000000001100101011101",
			1620 => "0000001001100101011101",
			1621 => "0000000001100101011101",
			1622 => "0000000001100101011101",
			1623 => "0001001111111100010000",
			1624 => "0000010110000000001100",
			1625 => "0001110001111100000100",
			1626 => "1111111001100110111001",
			1627 => "0000001000000000000100",
			1628 => "0000011001100110111001",
			1629 => "0000001001100110111001",
			1630 => "1111111001100110111001",
			1631 => "0000111111000100000100",
			1632 => "1111111001100110111001",
			1633 => "0001000011100100010100",
			1634 => "0011110000001100001000",
			1635 => "0001001111111000000100",
			1636 => "0000001001100110111001",
			1637 => "1111111001100110111001",
			1638 => "0000011110011100000100",
			1639 => "0000001001100110111001",
			1640 => "0000101000101000000100",
			1641 => "0000001001100110111001",
			1642 => "0000001001100110111001",
			1643 => "0001101100011000000100",
			1644 => "1111111001100110111001",
			1645 => "0000000001100110111001",
			1646 => "0001001111111100011000",
			1647 => "0000010000011000010100",
			1648 => "0000011100100000001000",
			1649 => "0010101111001000000100",
			1650 => "0000000001101000101101",
			1651 => "0000000001101000101101",
			1652 => "0010000001110100000100",
			1653 => "0000000001101000101101",
			1654 => "0010100110011100000100",
			1655 => "0000000001101000101101",
			1656 => "0000000001101000101101",
			1657 => "1111111001101000101101",
			1658 => "0000100011001000010000",
			1659 => "0000001101000100001100",
			1660 => "0010100001110100001000",
			1661 => "0010100111000100000100",
			1662 => "0000000001101000101101",
			1663 => "0000000001101000101101",
			1664 => "0000000001101000101101",
			1665 => "1111111001101000101101",
			1666 => "0001000101101000001000",
			1667 => "0001101101011000000100",
			1668 => "0000001001101000101101",
			1669 => "0000000001101000101101",
			1670 => "0001101100011000000100",
			1671 => "0000000001101000101101",
			1672 => "0000100110010000000100",
			1673 => "0000000001101000101101",
			1674 => "0000000001101000101101",
			1675 => "0010010000011000100000",
			1676 => "0011110000001100001000",
			1677 => "0000011110011100000100",
			1678 => "0000000001101010001001",
			1679 => "0000000001101010001001",
			1680 => "0000111111000100000100",
			1681 => "0000000001101010001001",
			1682 => "0010011100100000000100",
			1683 => "0000000001101010001001",
			1684 => "0010111000000000001100",
			1685 => "0000000101001000001000",
			1686 => "0010100010111100000100",
			1687 => "0000001001101010001001",
			1688 => "0000000001101010001001",
			1689 => "0000000001101010001001",
			1690 => "0000000001101010001001",
			1691 => "0000000110110100001100",
			1692 => "0001101110010100000100",
			1693 => "0000000001101010001001",
			1694 => "0000011100100000000100",
			1695 => "0000000001101010001001",
			1696 => "1111111001101010001001",
			1697 => "0000000001101010001001",
			1698 => "0001001111111100010100",
			1699 => "0000010000011000001000",
			1700 => "0001011000011000000100",
			1701 => "1111111001101011101101",
			1702 => "0000010001101011101101",
			1703 => "0000010110000000001000",
			1704 => "0000010110000000000100",
			1705 => "1111111001101011101101",
			1706 => "1111111001101011101101",
			1707 => "1111111001101011101101",
			1708 => "0000111111000100000100",
			1709 => "1111111001101011101101",
			1710 => "0001000011100100010100",
			1711 => "0011111101111000000100",
			1712 => "1111111001101011101101",
			1713 => "0010011100100000000100",
			1714 => "0000000001101011101101",
			1715 => "0011110000001100000100",
			1716 => "0000001001101011101101",
			1717 => "0011110100001000000100",
			1718 => "0000001001101011101101",
			1719 => "0000001001101011101101",
			1720 => "0001101100011000000100",
			1721 => "1111111001101011101101",
			1722 => "0000000001101011101101",
			1723 => "0000001010001100010100",
			1724 => "0010011100110100001000",
			1725 => "0001010100011000000100",
			1726 => "1111111001101101010001",
			1727 => "0000001001101101010001",
			1728 => "0000000110000100000100",
			1729 => "1111111001101101010001",
			1730 => "0011110100010000000100",
			1731 => "0000001001101101010001",
			1732 => "1111111001101101010001",
			1733 => "0000111111000100000100",
			1734 => "1111111001101101010001",
			1735 => "0001101000010000011000",
			1736 => "0010011100100000010000",
			1737 => "0001101100011000001000",
			1738 => "0001101100011000000100",
			1739 => "1111111001101101010001",
			1740 => "0000000001101101010001",
			1741 => "0010100010111100000100",
			1742 => "0000001001101101010001",
			1743 => "0000000001101101010001",
			1744 => "0010001101111000000100",
			1745 => "0000001001101101010001",
			1746 => "0000000001101101010001",
			1747 => "1111111001101101010001",
			1748 => "0001001111111100010000",
			1749 => "0000010110000000001100",
			1750 => "0001010100011000000100",
			1751 => "1111111001101110101101",
			1752 => "0011101111000100000100",
			1753 => "0000001001101110101101",
			1754 => "0000010001101110101101",
			1755 => "1111111001101110101101",
			1756 => "0000111111000100000100",
			1757 => "1111111001101110101101",
			1758 => "0010011100100000001000",
			1759 => "0001101100011000000100",
			1760 => "1111111001101110101101",
			1761 => "0000000001101110101101",
			1762 => "0001000011100100010000",
			1763 => "0011111101111000000100",
			1764 => "0000000001101110101101",
			1765 => "0001000101101000000100",
			1766 => "0000001001101110101101",
			1767 => "0011111010111000000100",
			1768 => "0000000001101110101101",
			1769 => "0000001001101110101101",
			1770 => "0000000001101110101101",
			1771 => "0001001111111100100000",
			1772 => "0010011110100000011100",
			1773 => "0010010000011000001000",
			1774 => "0010010000011000000100",
			1775 => "1111111001110000101001",
			1776 => "0000000001110000101001",
			1777 => "0000011100100000001000",
			1778 => "0000001100001000000100",
			1779 => "0000001001110000101001",
			1780 => "0000000001110000101001",
			1781 => "0001001110001000001000",
			1782 => "0000010000011000000100",
			1783 => "0000000001110000101001",
			1784 => "0000000001110000101001",
			1785 => "0000000001110000101001",
			1786 => "1111111001110000101001",
			1787 => "0000110010011000001100",
			1788 => "0000001100100100001000",
			1789 => "0000111111000100000100",
			1790 => "0000000001110000101001",
			1791 => "0000000001110000101001",
			1792 => "1111111001110000101001",
			1793 => "0000101000101000010000",
			1794 => "0001000001100000001000",
			1795 => "0000101010001000000100",
			1796 => "0000000001110000101001",
			1797 => "0000001001110000101001",
			1798 => "0001101100011000000100",
			1799 => "1111111001110000101001",
			1800 => "0000001001110000101001",
			1801 => "0000000001110000101001",
			1802 => "0000001010001100010000",
			1803 => "0000010000011000001100",
			1804 => "0001010100011000000100",
			1805 => "1111111001110010001101",
			1806 => "0000001001001000000100",
			1807 => "0000010001110010001101",
			1808 => "0000001001110010001101",
			1809 => "1111111001110010001101",
			1810 => "0000111111000100000100",
			1811 => "1111111001110010001101",
			1812 => "0001101001100100011000",
			1813 => "0010011100100000001000",
			1814 => "0001101100011000000100",
			1815 => "1111111001110010001101",
			1816 => "0000001001110010001101",
			1817 => "0000001111010000001100",
			1818 => "0000100100101000000100",
			1819 => "0000000001110010001101",
			1820 => "0000000101001000000100",
			1821 => "0000001001110010001101",
			1822 => "0000001001110010001101",
			1823 => "1111111001110010001101",
			1824 => "0010001100110000000100",
			1825 => "1111111001110010001101",
			1826 => "0000000001110010001101",
			1827 => "0001001111111100010000",
			1828 => "0000010110000000001100",
			1829 => "0001011000011000000100",
			1830 => "1111111001110011110001",
			1831 => "0001001111110000000100",
			1832 => "0000010001110011110001",
			1833 => "0000001001110011110001",
			1834 => "1111111001110011110001",
			1835 => "0000111111000100000100",
			1836 => "1111111001110011110001",
			1837 => "0010011100100000001000",
			1838 => "0011001010111100000100",
			1839 => "1111111001110011110001",
			1840 => "0000000001110011110001",
			1841 => "0010100010111100010100",
			1842 => "0001000001100000001100",
			1843 => "0000100111111100000100",
			1844 => "0000000001110011110001",
			1845 => "0000101000101000000100",
			1846 => "0000001001110011110001",
			1847 => "0000000001110011110001",
			1848 => "0001101100011000000100",
			1849 => "1111111001110011110001",
			1850 => "0000001001110011110001",
			1851 => "1111111001110011110001",
			1852 => "0001000010010000000100",
			1853 => "1111111001110101001101",
			1854 => "0000100101110000001000",
			1855 => "0000110000111000000100",
			1856 => "1111111001110101001101",
			1857 => "0000000001110101001101",
			1858 => "0001101101011000011000",
			1859 => "0000001100100100001100",
			1860 => "0001110101101100000100",
			1861 => "0000000001110101001101",
			1862 => "0000010010001100000100",
			1863 => "0000001001110101001101",
			1864 => "0000000001110101001101",
			1865 => "0001101100011000000100",
			1866 => "0000000001110101001101",
			1867 => "0000101100010100000100",
			1868 => "0000000001110101001101",
			1869 => "0000000001110101001101",
			1870 => "0001101001100100000100",
			1871 => "0000000001110101001101",
			1872 => "0001111110001100000100",
			1873 => "0000000001110101001101",
			1874 => "0000000001110101001101",
			1875 => "0001001111111100010000",
			1876 => "0000010110000000001100",
			1877 => "0001011000011000000100",
			1878 => "1111111001110110110001",
			1879 => "0010111000000000000100",
			1880 => "0000001001110110110001",
			1881 => "0000010001110110110001",
			1882 => "1111111001110110110001",
			1883 => "0000111111000100000100",
			1884 => "1111111001110110110001",
			1885 => "0010011100100000001000",
			1886 => "0011001010111100000100",
			1887 => "1111111001110110110001",
			1888 => "0000000001110110110001",
			1889 => "0010100010111100010100",
			1890 => "0011111101111000000100",
			1891 => "0000000001110110110001",
			1892 => "0001000001100000001000",
			1893 => "0000101000101000000100",
			1894 => "0000001001110110110001",
			1895 => "0000000001110110110001",
			1896 => "0001101100011000000100",
			1897 => "1111111001110110110001",
			1898 => "0000001001110110110001",
			1899 => "1111111001110110110001",
			1900 => "0001001111111100101000",
			1901 => "0001000100100100011100",
			1902 => "0000010110000000011000",
			1903 => "0010011001111000010100",
			1904 => "0001000010010000000100",
			1905 => "1111111001111000110101",
			1906 => "0010010110000000001000",
			1907 => "0001000110110000000100",
			1908 => "0000000001111000110101",
			1909 => "1111111001111000110101",
			1910 => "0001001011100100000100",
			1911 => "1111111001111000110101",
			1912 => "0000010001111000110101",
			1913 => "0000001001111000110101",
			1914 => "1111111001111000110101",
			1915 => "0001011000011000000100",
			1916 => "1111111001111000110101",
			1917 => "0000011101101000000100",
			1918 => "0000010001111000110101",
			1919 => "1111111001111000110101",
			1920 => "0011111101111000000100",
			1921 => "1111111001111000110101",
			1922 => "0010011100100000001000",
			1923 => "0001101100011000000100",
			1924 => "1111111001111000110101",
			1925 => "0000000001111000110101",
			1926 => "0000001111010000001100",
			1927 => "0000000101001000001000",
			1928 => "0010111110001100000100",
			1929 => "0000001001111000110101",
			1930 => "0000010001111000110101",
			1931 => "0000001001111000110101",
			1932 => "1111111001111000110101",
			1933 => "0001001111111100100100",
			1934 => "0001000101001100000100",
			1935 => "1111111001111010111011",
			1936 => "0010101100000100001000",
			1937 => "0001111101111000000100",
			1938 => "1111111001111010111011",
			1939 => "0000010001111010111011",
			1940 => "0001001101100100010000",
			1941 => "0010000011010000001100",
			1942 => "0010101001101000000100",
			1943 => "1111111001111010111011",
			1944 => "0010101001101000000100",
			1945 => "0000001001111010111011",
			1946 => "0000000001111010111011",
			1947 => "1111111001111010111011",
			1948 => "0000111010000000000100",
			1949 => "1111111001111010111011",
			1950 => "0000001001111010111011",
			1951 => "0000111111000100000100",
			1952 => "1111111001111010111011",
			1953 => "0010100010111100011000",
			1954 => "0011111101111000000100",
			1955 => "0000000001111010111011",
			1956 => "0001000001100000001100",
			1957 => "0000101000101000001000",
			1958 => "0000101110010000000100",
			1959 => "0000001001111010111011",
			1960 => "0000001001111010111011",
			1961 => "0000000001111010111011",
			1962 => "0001101100011000000100",
			1963 => "1111111001111010111011",
			1964 => "0000001001111010111011",
			1965 => "1111111001111010111011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(638, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1284, initial_addr_3'length));
	end generate gen_rom_1;

	gen_rom_2: if SELECT_ROM = 2 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0011001011000000000100",
			4 => "0000000000000000100001",
			5 => "0011000110100100000100",
			6 => "0000000000000000100001",
			7 => "0000000000000000100001",
			8 => "0010110100010000001000",
			9 => "0010110000011100000100",
			10 => "0000000000000000110101",
			11 => "0000000000000000110101",
			12 => "0000000000000000110101",
			13 => "0010111011011100000100",
			14 => "0000000000000001001001",
			15 => "0010110001001000000100",
			16 => "0000000000000001001001",
			17 => "0000000000000001001001",
			18 => "0000001001101000001000",
			19 => "0011001010111000000100",
			20 => "0000000000000001100101",
			21 => "0000000000000001100101",
			22 => "0011001001110100000100",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0001011100100100001000",
			26 => "0001010110110100000100",
			27 => "0000000000000010000001",
			28 => "0000000000000010000001",
			29 => "0001011111010000000100",
			30 => "0000000000000010000001",
			31 => "0000000000000010000001",
			32 => "0010111011011100000100",
			33 => "0000000000000010011101",
			34 => "0000101100000000001000",
			35 => "0000100010000000000100",
			36 => "0000000000000010011101",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0000101100010000001100",
			40 => "0000001100000100001000",
			41 => "0000101101000100000100",
			42 => "0000000000000011000001",
			43 => "0000000000000011000001",
			44 => "0000000000000011000001",
			45 => "0000101010000100000100",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0000001001101000001100",
			49 => "0000101101000100000100",
			50 => "0000000000000011100101",
			51 => "0000101010000100000100",
			52 => "0000000000000011100101",
			53 => "0000000000000011100101",
			54 => "0000101000101000000100",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0000001100000100001100",
			58 => "0000101100000000001000",
			59 => "0000101101000100000100",
			60 => "0000000000000100010001",
			61 => "0000000000000100010001",
			62 => "0000000000000100010001",
			63 => "0000101000001100000100",
			64 => "0000000000000100010001",
			65 => "0000101101101100000100",
			66 => "0000000000000100010001",
			67 => "0000000000000100010001",
			68 => "0000000001110100010000",
			69 => "0010011111000000000100",
			70 => "0000000000000100110101",
			71 => "0001001110000000001000",
			72 => "0001000111011000000100",
			73 => "0000000000000100110101",
			74 => "0000000000000100110101",
			75 => "0000000000000100110101",
			76 => "0000000000000100110101",
			77 => "0001001101101100010000",
			78 => "0001110110100100000100",
			79 => "0000000000000101100001",
			80 => "0001000111011000000100",
			81 => "0000000000000101100001",
			82 => "0011000100011000000100",
			83 => "0000000000000101100001",
			84 => "0000000000000101100001",
			85 => "0011001001110100000100",
			86 => "0000000000000101100001",
			87 => "0000000000000101100001",
			88 => "0001101101111100001000",
			89 => "0011000100011000000100",
			90 => "0000000000000110001101",
			91 => "0000000000000110001101",
			92 => "0011001001110100001100",
			93 => "0001001010000100000100",
			94 => "0000000000000110001101",
			95 => "0001101011001100000100",
			96 => "0000000000000110001101",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0000001100000100001000",
			100 => "0010111001110100000100",
			101 => "0000000000000111000001",
			102 => "0000000000000111000001",
			103 => "0010110101100100001000",
			104 => "0010110000011100000100",
			105 => "0000000000000111000001",
			106 => "0000000000000111000001",
			107 => "0010110101110100001000",
			108 => "0010111011011100000100",
			109 => "0000000000000111000001",
			110 => "0000000000000111000001",
			111 => "0000000000000111000001",
			112 => "0000001100000100001000",
			113 => "0010111001110100000100",
			114 => "0000000000000111111101",
			115 => "0000000000000111111101",
			116 => "0010110101100100001000",
			117 => "0010110000011100000100",
			118 => "0000000000000111111101",
			119 => "0000000000000111111101",
			120 => "0010110101110100001000",
			121 => "0010111011011100000100",
			122 => "0000000000000111111101",
			123 => "0000000000000111111101",
			124 => "0010111011110100000100",
			125 => "0000000000000111111101",
			126 => "0000000000000111111101",
			127 => "0010111011011100001000",
			128 => "0010010111101100000100",
			129 => "0000000000001000110001",
			130 => "0000000000001000110001",
			131 => "0001110110100100000100",
			132 => "0000000000001000110001",
			133 => "0001111000011000001100",
			134 => "0010011111000000000100",
			135 => "0000000000001000110001",
			136 => "0010010010101100000100",
			137 => "0000000000001000110001",
			138 => "0000000000001000110001",
			139 => "0000000000001000110001",
			140 => "0011100111010100010100",
			141 => "0010110101110100010000",
			142 => "0001000110010000000100",
			143 => "0000000000001001011101",
			144 => "0001101101011000001000",
			145 => "0001111111011100000100",
			146 => "0000000000001001011101",
			147 => "0000000000001001011101",
			148 => "0000000000001001011101",
			149 => "0000000000001001011101",
			150 => "0000000000001001011101",
			151 => "0001000001011100010100",
			152 => "0010001000100100000100",
			153 => "0000000000001010011001",
			154 => "0011000100011000000100",
			155 => "0000000000001010011001",
			156 => "0011000001101000001000",
			157 => "0000001111001000000100",
			158 => "0000000000001010011001",
			159 => "0000000000001010011001",
			160 => "0000000000001010011001",
			161 => "0000011100011000001000",
			162 => "0011001011011100000100",
			163 => "0000000000001010011001",
			164 => "0000000000001010011001",
			165 => "0000000000001010011001",
			166 => "0011101100000000010000",
			167 => "0001001100010000000100",
			168 => "0000000000001011011101",
			169 => "0010100000001000000100",
			170 => "0000000000001011011101",
			171 => "0010101010100000000100",
			172 => "0000000000001011011101",
			173 => "0000000000001011011101",
			174 => "0001000001011100010000",
			175 => "0000011101111100001100",
			176 => "0000111000100000001000",
			177 => "0000111010000100000100",
			178 => "0000000000001011011101",
			179 => "0000000000001011011101",
			180 => "0000000000001011011101",
			181 => "0000000000001011011101",
			182 => "0000000000001011011101",
			183 => "0001001101101100011100",
			184 => "0011100111011000010100",
			185 => "0000001100000100001100",
			186 => "0000000001010100000100",
			187 => "0000000000001100110001",
			188 => "0000011001011000000100",
			189 => "0000000000001100110001",
			190 => "0000000000001100110001",
			191 => "0010110101100100000100",
			192 => "0000000000001100110001",
			193 => "0000000000001100110001",
			194 => "0000111010000100000100",
			195 => "0000000000001100110001",
			196 => "0000000000001100110001",
			197 => "0010011010100000001100",
			198 => "0001110101110100001000",
			199 => "0010000001010000000100",
			200 => "0000000000001100110001",
			201 => "0000000000001100110001",
			202 => "0000000000001100110001",
			203 => "0000000000001100110001",
			204 => "0001000001011100011000",
			205 => "0010010100111100000100",
			206 => "0000000000001101101101",
			207 => "0000011101111100010000",
			208 => "0001110110100100000100",
			209 => "0000000000001101101101",
			210 => "0000001111001000001000",
			211 => "0010110100000100000100",
			212 => "0000000000001101101101",
			213 => "0000000000001101101101",
			214 => "0000000000001101101101",
			215 => "0000000000001101101101",
			216 => "0001100100111100000100",
			217 => "0000000000001101101101",
			218 => "0000000000001101101101",
			219 => "0011101100000000001000",
			220 => "0011011001010100000100",
			221 => "0000000000001110101001",
			222 => "0000000000001110101001",
			223 => "0011010011001000010100",
			224 => "0010010100111100000100",
			225 => "0000000000001110101001",
			226 => "0011100010010100001100",
			227 => "0011011110000100000100",
			228 => "0000000000001110101001",
			229 => "0010010010101100000100",
			230 => "0000000000001110101001",
			231 => "0000000000001110101001",
			232 => "0000000000001110101001",
			233 => "0000000000001110101001",
			234 => "0000010000111100001000",
			235 => "0010000100101100000100",
			236 => "0000000000001111100101",
			237 => "0000000000001111100101",
			238 => "0011111011110000010100",
			239 => "0011101100010000000100",
			240 => "0000000000001111100101",
			241 => "0010010100111100000100",
			242 => "0000000000001111100101",
			243 => "0000011100011000001000",
			244 => "0010000001110000000100",
			245 => "0000000000001111100101",
			246 => "0000000000001111100101",
			247 => "0000000000001111100101",
			248 => "0000000000001111100101",
			249 => "0001001101101100011000",
			250 => "0000011001011000000100",
			251 => "0000000000010000101001",
			252 => "0000111000100000010000",
			253 => "0000001111001000001100",
			254 => "0011110010000100000100",
			255 => "0000000000010000101001",
			256 => "0000110010000100000100",
			257 => "0000000000010000101001",
			258 => "0000000000010000101001",
			259 => "0000000000010000101001",
			260 => "0000000000010000101001",
			261 => "0000010001111000001000",
			262 => "0000111111101000000100",
			263 => "0000000000010000101001",
			264 => "0000000000010000101001",
			265 => "0000000000010000101001",
			266 => "0011001010111000000100",
			267 => "0000000000010001011101",
			268 => "0001011111010000010100",
			269 => "0000000001110100010000",
			270 => "0011011010001000001100",
			271 => "0011011110000100000100",
			272 => "0000000000010001011101",
			273 => "0001111111011100000100",
			274 => "0000000000010001011101",
			275 => "0000000000010001011101",
			276 => "0000000000010001011101",
			277 => "0000000000010001011101",
			278 => "0000000000010001011101",
			279 => "0011001001110100011000",
			280 => "0001001100010000000100",
			281 => "0000000000010010010001",
			282 => "0010010111101100010000",
			283 => "0011001010111000000100",
			284 => "0000000000010010010001",
			285 => "0001111001001000000100",
			286 => "0000000000010010010001",
			287 => "0000010001111000000100",
			288 => "0000000000010010010001",
			289 => "0000000000010010010001",
			290 => "0000000000010010010001",
			291 => "0000000000010010010001",
			292 => "0001001011101100010000",
			293 => "0010100000001000000100",
			294 => "0000000000010011100101",
			295 => "0011010101001000000100",
			296 => "0000000000010011100101",
			297 => "0000111111100100000100",
			298 => "0000000000010011100101",
			299 => "0000000000010011100101",
			300 => "0010010111101100001000",
			301 => "0011001001110100000100",
			302 => "0000000000010011100101",
			303 => "0000000000010011100101",
			304 => "0011000110100100010000",
			305 => "0011100111010100000100",
			306 => "0000000000010011100101",
			307 => "0000011010011000001000",
			308 => "0000001010101100000100",
			309 => "0000000000010011100101",
			310 => "0000000000010011100101",
			311 => "0000000000010011100101",
			312 => "0000000000010011100101",
			313 => "0000001100000100001100",
			314 => "0010001000100100000100",
			315 => "0000000000010101000001",
			316 => "0010011111000000000100",
			317 => "0000000000010101000001",
			318 => "0000000000010101000001",
			319 => "0001100100111100010000",
			320 => "0010111011110100001100",
			321 => "0000100111011000000100",
			322 => "0000000000010101000001",
			323 => "0010001000010100000100",
			324 => "0000000000010101000001",
			325 => "0000000000010101000001",
			326 => "0000000000010101000001",
			327 => "0000001010101100010000",
			328 => "0010011010100000000100",
			329 => "0000000000010101000001",
			330 => "0010010011101000001000",
			331 => "0010110001001000000100",
			332 => "0000000000010101000001",
			333 => "0000000000010101000001",
			334 => "0000000000010101000001",
			335 => "0000000000010101000001",
			336 => "0001101001100100011000",
			337 => "0010111011110100010100",
			338 => "0000101010000100001100",
			339 => "0011101100000000001000",
			340 => "0011101110010000000100",
			341 => "0000000000010110011101",
			342 => "0000000000010110011101",
			343 => "0000000000010110011101",
			344 => "0010110000011100000100",
			345 => "0000000000010110011101",
			346 => "0000000000010110011101",
			347 => "0000000000010110011101",
			348 => "0010111010010100010100",
			349 => "0010010111101100000100",
			350 => "0000000000010110011101",
			351 => "0010101001000100001100",
			352 => "0011101000001100000100",
			353 => "0000000000010110011101",
			354 => "0011111110000000000100",
			355 => "0000000000010110011101",
			356 => "0000000000010110011101",
			357 => "0000000000010110011101",
			358 => "0000000000010110011101",
			359 => "0010111011011100010000",
			360 => "0011100111011000001000",
			361 => "0000111010000100000100",
			362 => "0000000000010111110001",
			363 => "0000000000010111110001",
			364 => "0010010000001000000100",
			365 => "0000000000010111110001",
			366 => "0000000000010111110001",
			367 => "0001110110100100000100",
			368 => "0000000000010111110001",
			369 => "0001001101101100010100",
			370 => "0000000101000100000100",
			371 => "0000000000010111110001",
			372 => "0001000111011000000100",
			373 => "0000000000010111110001",
			374 => "0000011001011000000100",
			375 => "0000000000010111110001",
			376 => "0011111100010000000100",
			377 => "0000000000010111110001",
			378 => "0000000000010111110001",
			379 => "0000000000010111110001",
			380 => "0000000111000100011100",
			381 => "0011001010111000000100",
			382 => "0000000000011000110101",
			383 => "0011011010001000010100",
			384 => "0011011110000100000100",
			385 => "0000000000011000110101",
			386 => "0010100000001000000100",
			387 => "0000000000011000110101",
			388 => "0010110001011000000100",
			389 => "0000000000011000110101",
			390 => "0010110101110100000100",
			391 => "0000000000011000110101",
			392 => "0000000000011000110101",
			393 => "0000000000011000110101",
			394 => "0001101000010000000100",
			395 => "0000000000011000110101",
			396 => "0000000000011000110101",
			397 => "0001001101101100100100",
			398 => "0011100111011000011100",
			399 => "0000001100000100010100",
			400 => "0010001000100100010000",
			401 => "0011010111111100001100",
			402 => "0011110010000000000100",
			403 => "0000000000011010010001",
			404 => "0011011110000100000100",
			405 => "0000000000011010010001",
			406 => "0000000000011010010001",
			407 => "0000000000011010010001",
			408 => "0000000000011010010001",
			409 => "0010110101100100000100",
			410 => "0000000000011010010001",
			411 => "0000000000011010010001",
			412 => "0000111010000100000100",
			413 => "0000000000011010010001",
			414 => "0000000000011010010001",
			415 => "0001100100111100001000",
			416 => "0011001111011100000100",
			417 => "0000000000011010010001",
			418 => "0000000000011010010001",
			419 => "0000000000011010010001",
			420 => "0001011111010000100100",
			421 => "0001011101000100001100",
			422 => "0000000001010100000100",
			423 => "0000000000011011110101",
			424 => "0000101000001100000100",
			425 => "0000000000011011110101",
			426 => "0000000000011011110101",
			427 => "0011001001001000010100",
			428 => "0001100100110100000100",
			429 => "0000000000011011110101",
			430 => "0000101101101100001100",
			431 => "0000010100110100001000",
			432 => "0000000001110100000100",
			433 => "0000000000011011110101",
			434 => "0000000000011011110101",
			435 => "0000000000011011110101",
			436 => "0000000000011011110101",
			437 => "0000000000011011110101",
			438 => "0010111011110100001100",
			439 => "0011100001011100001000",
			440 => "0010110010001000000100",
			441 => "0000000000011011110101",
			442 => "0000000000011011110101",
			443 => "0000000000011011110101",
			444 => "0000000000011011110101",
			445 => "0001000111010100010000",
			446 => "0010001000100100000100",
			447 => "0000000000011101011001",
			448 => "0011111111010100001000",
			449 => "0011100011001000000100",
			450 => "0000000000011101011001",
			451 => "0000000000011101011001",
			452 => "0000000000011101011001",
			453 => "0001100100111100011000",
			454 => "0010111011110100010100",
			455 => "0000001100000100000100",
			456 => "0000000000011101011001",
			457 => "0001101111000000001100",
			458 => "0010110000011100000100",
			459 => "0000000000011101011001",
			460 => "0010001000010100000100",
			461 => "0000000000011101011001",
			462 => "0000000000011101011001",
			463 => "0000000000011101011001",
			464 => "0000000000011101011001",
			465 => "0000001010101100001000",
			466 => "0000011010011000000100",
			467 => "0000000000011101011001",
			468 => "0000000000011101011001",
			469 => "0000000000011101011001",
			470 => "0001001100010000000100",
			471 => "0000000000011110010101",
			472 => "0001011111010000011000",
			473 => "0011100111010100010100",
			474 => "0010110100010000010000",
			475 => "0011001010111000000100",
			476 => "0000000000011110010101",
			477 => "0010110000011100000100",
			478 => "0000000000011110010101",
			479 => "0000110000010000000100",
			480 => "0000000000011110010101",
			481 => "0000000000011110010101",
			482 => "0000000000011110010101",
			483 => "0000000000011110010101",
			484 => "0000000000011110010101",
			485 => "0011100111010100011100",
			486 => "0010110101110100011000",
			487 => "0001011100100100000100",
			488 => "0000000000011111010001",
			489 => "0000011001011000000100",
			490 => "0000000000011111010001",
			491 => "0001011111010000001100",
			492 => "0010100010101100001000",
			493 => "0001111111011100000100",
			494 => "0000000000011111010001",
			495 => "0000000000011111010001",
			496 => "0000000000011111010001",
			497 => "0000000000011111010001",
			498 => "0000000000011111010001",
			499 => "0000000000011111010001",
			500 => "0010011111000000000100",
			501 => "0000000000100000001101",
			502 => "0000000111000100011000",
			503 => "0011011010001000010100",
			504 => "0011011110000100000100",
			505 => "0000000000100000001101",
			506 => "0010110000011100000100",
			507 => "0000000000100000001101",
			508 => "0010100000001000000100",
			509 => "0000000000100000001101",
			510 => "0011001010111000000100",
			511 => "0000000000100000001101",
			512 => "0000000000100000001101",
			513 => "0000000000100000001101",
			514 => "0000000000100000001101",
			515 => "0000000010101000011100",
			516 => "0010011111000000000100",
			517 => "0000000000100001001001",
			518 => "0001110110100100000100",
			519 => "0000000000100001001001",
			520 => "0000000001010100000100",
			521 => "0000000000100001001001",
			522 => "0000011010011000001100",
			523 => "0011001010111000000100",
			524 => "0000000000100001001001",
			525 => "0001000111011000000100",
			526 => "0000000000100001001001",
			527 => "0000000000100001001001",
			528 => "0000000000100001001001",
			529 => "0000000000100001001001",
			530 => "0000010000111100010100",
			531 => "0000101100010000000100",
			532 => "0000000000100010100101",
			533 => "0011010111111100000100",
			534 => "0000000000100010100101",
			535 => "0001010101110000001000",
			536 => "0011101100010000000100",
			537 => "0000000000100010100101",
			538 => "0000000000100010100101",
			539 => "0000000000100010100101",
			540 => "0000000001110100011000",
			541 => "0011000100011000000100",
			542 => "0000000000100010100101",
			543 => "0011101100000000000100",
			544 => "0000000000100010100101",
			545 => "0000011101111100001100",
			546 => "0000101101101100001000",
			547 => "0001010110100000000100",
			548 => "0000000000100010100101",
			549 => "0000000000100010100101",
			550 => "0000000000100010100101",
			551 => "0000000000100010100101",
			552 => "0000000000100010100101",
			553 => "0001001111100100011000",
			554 => "0011111110110100000100",
			555 => "0000000000100100011001",
			556 => "0000110000010000010000",
			557 => "0010101010100000000100",
			558 => "0000000000100100011001",
			559 => "0001110110100100000100",
			560 => "0000000000100100011001",
			561 => "0010100011101000000100",
			562 => "0000000000100100011001",
			563 => "0000000000100100011001",
			564 => "0000000000100100011001",
			565 => "0000111111100100010000",
			566 => "0011001010111000000100",
			567 => "0000000000100100011001",
			568 => "0001010010110100000100",
			569 => "0000000000100100011001",
			570 => "0001010111100000000100",
			571 => "0000000000100100011001",
			572 => "0000000000100100011001",
			573 => "0000011110010100000100",
			574 => "0000000000100100011001",
			575 => "0000101011110000001100",
			576 => "0000011010011000001000",
			577 => "0011111011110000000100",
			578 => "0000000000100100011001",
			579 => "0000000000100100011001",
			580 => "0000000000100100011001",
			581 => "0000000000100100011001",
			582 => "0010111011011100010000",
			583 => "0001001010000100000100",
			584 => "0000000000100110010101",
			585 => "0011100111010100001000",
			586 => "0001010111100000000100",
			587 => "0000000000100110010101",
			588 => "0000000000100110010101",
			589 => "0000000000100110010101",
			590 => "0001100100110100010000",
			591 => "0010110010001000000100",
			592 => "0000000000100110010101",
			593 => "0001011001010000001000",
			594 => "0011001011000000000100",
			595 => "0000000000100110010101",
			596 => "0000000000100110010101",
			597 => "0000000000100110010101",
			598 => "0001000001011100001000",
			599 => "0001110110100100000100",
			600 => "0000000000100110010101",
			601 => "0000000000100110010101",
			602 => "0010011010100000001000",
			603 => "0010110001001000000100",
			604 => "0000000000100110010101",
			605 => "0000000000100110010101",
			606 => "0000011010011000001100",
			607 => "0011011100010100001000",
			608 => "0000111000100000000100",
			609 => "0000000000100110010101",
			610 => "0000000000100110010101",
			611 => "0000000000100110010101",
			612 => "0000000000100110010101",
			613 => "0011001011000000101100",
			614 => "0001000110111100010000",
			615 => "0011001010111000000100",
			616 => "0000000000101000011001",
			617 => "0001111000011000001000",
			618 => "0001111011000000000100",
			619 => "0000000000101000011001",
			620 => "0000000000101000011001",
			621 => "0000000000101000011001",
			622 => "0010010111101100001100",
			623 => "0001011110101000000100",
			624 => "0000000000101000011001",
			625 => "0011101100010000000100",
			626 => "0000000000101000011001",
			627 => "0000000000101000011001",
			628 => "0000011101111100001100",
			629 => "0011101111010100000100",
			630 => "0000000000101000011001",
			631 => "0010101000100100000100",
			632 => "0000000000101000011001",
			633 => "0000000000101000011001",
			634 => "0000000000101000011001",
			635 => "0010110100010000000100",
			636 => "0000000000101000011001",
			637 => "0000011100011000010000",
			638 => "0001111000011000000100",
			639 => "0000000000101000011001",
			640 => "0011111011110000001000",
			641 => "0000000111000000000100",
			642 => "0000000000101000011001",
			643 => "0000000000101000011001",
			644 => "0000000000101000011001",
			645 => "0000000000101000011001",
			646 => "0001101101111100010000",
			647 => "0001111011000000000100",
			648 => "0000000000101010010101",
			649 => "0001111111011100001000",
			650 => "0000101100000000000100",
			651 => "0000000000101010010101",
			652 => "0000000000101010010101",
			653 => "0000000000101010010101",
			654 => "0001111000011000100100",
			655 => "0010010100101100010000",
			656 => "0001011100100100000100",
			657 => "0000000000101010010101",
			658 => "0011011001011100001000",
			659 => "0011010010011100000100",
			660 => "0000000000101010010101",
			661 => "0000000000101010010101",
			662 => "0000000000101010010101",
			663 => "0010101000100100010000",
			664 => "0010100010101100000100",
			665 => "0000000000101010010101",
			666 => "0000101101101100001000",
			667 => "0000100010000100000100",
			668 => "0000000000101010010101",
			669 => "0000000000101010010101",
			670 => "0000000000101010010101",
			671 => "0000000000101010010101",
			672 => "0000111000100000001000",
			673 => "0010000110011100000100",
			674 => "0000000000101010010101",
			675 => "0000000000101010010101",
			676 => "0000000000101010010101",
			677 => "0011001001110100110000",
			678 => "0001100100111100100100",
			679 => "0001001111100100011000",
			680 => "0000100110111100010000",
			681 => "0000101110110100000100",
			682 => "0000000000101100011001",
			683 => "0010100010101100001000",
			684 => "0011110010000100000100",
			685 => "0000000000101100011001",
			686 => "0000000000101100011001",
			687 => "0000000000101100011001",
			688 => "0001101100011000000100",
			689 => "0000000000101100011001",
			690 => "0000000000101100011001",
			691 => "0001110110100100000100",
			692 => "0000000000101100011001",
			693 => "0001101101011000000100",
			694 => "0000000000101100011001",
			695 => "0000000000101100011001",
			696 => "0000000010101000001000",
			697 => "0000111100111000000100",
			698 => "0000000000101100011001",
			699 => "0000000000101100011001",
			700 => "0000000000101100011001",
			701 => "0000100010010100010000",
			702 => "0010001000100100000100",
			703 => "0000000000101100011001",
			704 => "0001110101100100001000",
			705 => "0000011100011000000100",
			706 => "0000000000101100011001",
			707 => "0000000000101100011001",
			708 => "0000000000101100011001",
			709 => "0000000000101100011001",
			710 => "0001001011101100111000",
			711 => "0011001011000000100100",
			712 => "0001110110100100010000",
			713 => "0001111001001000000100",
			714 => "0000000000101110110101",
			715 => "0010100010101100001000",
			716 => "0001001001100000000100",
			717 => "0000000000101110110101",
			718 => "0000000000101110110101",
			719 => "0000000000101110110101",
			720 => "0001101101111100000100",
			721 => "0000000000101110110101",
			722 => "0001001000100000001100",
			723 => "0001011111010000001000",
			724 => "0010100000001000000100",
			725 => "0000000000101110110101",
			726 => "0000000000101110110101",
			727 => "0000000000101110110101",
			728 => "0000000000101110110101",
			729 => "0001010111100000001100",
			730 => "0010010100101100001000",
			731 => "0001000010000100000100",
			732 => "0000000000101110110101",
			733 => "0000000000101110110101",
			734 => "0000000000101110110101",
			735 => "0000101110110100000100",
			736 => "0000000000101110110101",
			737 => "0000000000101110110101",
			738 => "0001101001100100001100",
			739 => "0011001001110100001000",
			740 => "0000001011010100000100",
			741 => "0000000000101110110101",
			742 => "0000000000101110110101",
			743 => "0000000000101110110101",
			744 => "0000000111000100001000",
			745 => "0001110111010000000100",
			746 => "0000000000101110110101",
			747 => "0000000000101110110101",
			748 => "0000000000101110110101",
			749 => "0001000001011100110000",
			750 => "0010110100010000101000",
			751 => "0011010101110000010100",
			752 => "0011011110000100000100",
			753 => "0000000000110000101001",
			754 => "0010011111000000000100",
			755 => "0000000000110000101001",
			756 => "0010010111101100001000",
			757 => "0010100000001000000100",
			758 => "0000000000110000101001",
			759 => "0000000000110000101001",
			760 => "0000000000110000101001",
			761 => "0010000001010000010000",
			762 => "0011010111111100001100",
			763 => "0010011111000000000100",
			764 => "0000000000110000101001",
			765 => "0000100110010000000100",
			766 => "0000000000110000101001",
			767 => "0000000000110000101001",
			768 => "0000000000110000101001",
			769 => "0000000000110000101001",
			770 => "0000111000100000000100",
			771 => "0000000000110000101001",
			772 => "0000000000110000101001",
			773 => "0011001001110100001000",
			774 => "0000110010010100000100",
			775 => "0000000000110000101001",
			776 => "0000000000110000101001",
			777 => "0000000000110000101001",
			778 => "0010111011011100010100",
			779 => "0000001100000100001100",
			780 => "0011001011000000001000",
			781 => "0011001101010100000100",
			782 => "0000000000110011000101",
			783 => "0000000000110011000101",
			784 => "0000000000110011000101",
			785 => "0011100111010100000100",
			786 => "0000000000110011000101",
			787 => "0000000000110011000101",
			788 => "0001100100110100010100",
			789 => "0011101100010000010000",
			790 => "0011010010011100000100",
			791 => "0000000000110011000101",
			792 => "0011000100011000000100",
			793 => "0000000000110011000101",
			794 => "0011100010000000000100",
			795 => "0000000000110011000101",
			796 => "0000000000110011000101",
			797 => "0000000000110011000101",
			798 => "0001000001011100001100",
			799 => "0010011111000000000100",
			800 => "0000000000110011000101",
			801 => "0001110110100100000100",
			802 => "0000000000110011000101",
			803 => "0000000000110011000101",
			804 => "0010011010100000001100",
			805 => "0010110001001000001000",
			806 => "0010011010100000000100",
			807 => "0000000000110011000101",
			808 => "0000000000110011000101",
			809 => "0000000000110011000101",
			810 => "0000011010011000001100",
			811 => "0011011100010100001000",
			812 => "0000001010101100000100",
			813 => "0000000000110011000101",
			814 => "0000000000110011000101",
			815 => "0000000000110011000101",
			816 => "0000000000110011000101",
			817 => "0000001001101000101100",
			818 => "0011101010000100100100",
			819 => "0011001010111000000100",
			820 => "0000000000110101100001",
			821 => "0010101010100000010000",
			822 => "0010011111000000001000",
			823 => "0000111111010100000100",
			824 => "0000000000110101100001",
			825 => "0000000000110101100001",
			826 => "0000100010000000000100",
			827 => "0000000000110101100001",
			828 => "0000000000110101100001",
			829 => "0001010110100000000100",
			830 => "0000000000110101100001",
			831 => "0001110110100100000100",
			832 => "0000000000110101100001",
			833 => "0000111011111000000100",
			834 => "0000000000110101100001",
			835 => "0000000000110101100001",
			836 => "0011001001001000000100",
			837 => "0000000000110101100001",
			838 => "0000000000110101100001",
			839 => "0001101001100100010000",
			840 => "0001001011101100001000",
			841 => "0001000110101100000100",
			842 => "0000000000110101100001",
			843 => "0000000000110101100001",
			844 => "0011001001110100000100",
			845 => "0000000000110101100001",
			846 => "0000000000110101100001",
			847 => "0011001001110100010000",
			848 => "0001000101000000001100",
			849 => "0011000100011000000100",
			850 => "0000000000110101100001",
			851 => "0010101001000100000100",
			852 => "0000000000110101100001",
			853 => "0000000000110101100001",
			854 => "0000000000110101100001",
			855 => "0000000000110101100001",
			856 => "0000001010101100101000",
			857 => "0011001101010100000100",
			858 => "1111111000110110110101",
			859 => "0001011110010000100000",
			860 => "0011101101101100010100",
			861 => "0010011111000000001000",
			862 => "0000100001000000000100",
			863 => "0000001000110110110101",
			864 => "1111111000110110110101",
			865 => "0000000001110100001000",
			866 => "0011001001110100000100",
			867 => "0000000000110110110101",
			868 => "0000001000110110110101",
			869 => "1111111000110110110101",
			870 => "0000001010101100001000",
			871 => "0010000001010100000100",
			872 => "0000000000110110110101",
			873 => "0000001000110110110101",
			874 => "0000010000110110110101",
			875 => "1111111000110110110101",
			876 => "1111111000110110110101",
			877 => "0001001000001100100000",
			878 => "0011001010111000000100",
			879 => "0000000000111001100001",
			880 => "0001111000011000001100",
			881 => "0000011011111100001000",
			882 => "0000011001011000000100",
			883 => "0000000000111001100001",
			884 => "0000000000111001100001",
			885 => "0000000000111001100001",
			886 => "0000000001010100001000",
			887 => "0000000101000100000100",
			888 => "0000000000111001100001",
			889 => "0000000000111001100001",
			890 => "0000000001010100000100",
			891 => "0000000000111001100001",
			892 => "0000000000111001100001",
			893 => "0000111010000100010000",
			894 => "0011001011000000001100",
			895 => "0001110001101000001000",
			896 => "0011101111010100000100",
			897 => "1111111000111001100001",
			898 => "0000000000111001100001",
			899 => "0000000000111001100001",
			900 => "0000000000111001100001",
			901 => "0000101000001100001000",
			902 => "0000010000111100000100",
			903 => "0000000000111001100001",
			904 => "0000000000111001100001",
			905 => "0011100111010100001100",
			906 => "0011001011000000001000",
			907 => "0001110110100100000100",
			908 => "0000000000111001100001",
			909 => "0000000000111001100001",
			910 => "0000000000111001100001",
			911 => "0000101011111000000100",
			912 => "0000000000111001100001",
			913 => "0000010001111000001000",
			914 => "0001110001011000000100",
			915 => "0000000000111001100001",
			916 => "0000000000111001100001",
			917 => "0000010100110100000100",
			918 => "0000000000111001100001",
			919 => "0000000000111001100001",
			920 => "0000001010101100101000",
			921 => "0011001101010100000100",
			922 => "1111111000111010110101",
			923 => "0011011001100000100000",
			924 => "0011101101101100011000",
			925 => "0010011111000000001000",
			926 => "0010101001111100000100",
			927 => "0000001000111010110101",
			928 => "1111111000111010110101",
			929 => "0011001001110100001000",
			930 => "0011011110010000000100",
			931 => "0000000000111010110101",
			932 => "1111111000111010110101",
			933 => "0000010100110100000100",
			934 => "0000001000111010110101",
			935 => "0000000000111010110101",
			936 => "0000001010101100000100",
			937 => "0000001000111010110101",
			938 => "0000010000111010110101",
			939 => "1111111000111010110101",
			940 => "1111111000111010110101",
			941 => "0001001011110000111100",
			942 => "0010011111000000010000",
			943 => "0010110010001000001100",
			944 => "0001100000111100001000",
			945 => "0010001001111100000100",
			946 => "1111111000111101010001",
			947 => "0000001000111101010001",
			948 => "1111111000111101010001",
			949 => "0000000000111101010001",
			950 => "0011010001000000001000",
			951 => "0001101010011000000100",
			952 => "0000000000111101010001",
			953 => "1111111000111101010001",
			954 => "0011010110010000011100",
			955 => "0011101011101100010000",
			956 => "0001000001011100001000",
			957 => "0010100000001000000100",
			958 => "0000000000111101010001",
			959 => "0000001000111101010001",
			960 => "0011101000001100000100",
			961 => "1111111000111101010001",
			962 => "0000001000111101010001",
			963 => "0001111000011000001000",
			964 => "0010000101000100000100",
			965 => "0000001000111101010001",
			966 => "0000000000111101010001",
			967 => "0000010000111101010001",
			968 => "0011000100000100000100",
			969 => "1111111000111101010001",
			970 => "0000000000111101010001",
			971 => "0001000101000000010000",
			972 => "0001101000010000000100",
			973 => "1111111000111101010001",
			974 => "0001011111010000000100",
			975 => "1111111000111101010001",
			976 => "0000011010011000000100",
			977 => "0000010000111101010001",
			978 => "1111111000111101010001",
			979 => "1111111000111101010001",
			980 => "0000000111000101000000",
			981 => "0001101101011000110000",
			982 => "0000011011111100100100",
			983 => "0000110110111100010000",
			984 => "0001101101111100000100",
			985 => "0000000000111111011101",
			986 => "0001000111010100001000",
			987 => "0010100000001000000100",
			988 => "0000000000111111011101",
			989 => "0000000000111111011101",
			990 => "0000000000111111011101",
			991 => "0011001001110100001100",
			992 => "0001101101111100000100",
			993 => "0000000000111111011101",
			994 => "0000010001000100000100",
			995 => "0000000000111111011101",
			996 => "0000000000111111011101",
			997 => "0011110111011000000100",
			998 => "0000000000111111011101",
			999 => "0000000000111111011101",
			1000 => "0010100010101100001000",
			1001 => "0001111001001000000100",
			1002 => "0000000000111111011101",
			1003 => "0000000000111111011101",
			1004 => "0000000000111111011101",
			1005 => "0010011001111100000100",
			1006 => "0000000000111111011101",
			1007 => "0011000100011000000100",
			1008 => "0000000000111111011101",
			1009 => "0000110110111100000100",
			1010 => "0000000000111111011101",
			1011 => "0000001000111111011101",
			1012 => "0001100100111100000100",
			1013 => "0000000000111111011101",
			1014 => "0000000000111111011101",
			1015 => "0011111100000000001100",
			1016 => "0001001100010000000100",
			1017 => "0000000001000010001001",
			1018 => "0010001000100100000100",
			1019 => "0000000001000010001001",
			1020 => "0000000001000010001001",
			1021 => "0001000001011100100000",
			1022 => "0010100010101100010100",
			1023 => "0001011111010000001100",
			1024 => "0000101100010000000100",
			1025 => "0000000001000010001001",
			1026 => "0001011100100100000100",
			1027 => "0000000001000010001001",
			1028 => "0000000001000010001001",
			1029 => "0000011001011000000100",
			1030 => "0000000001000010001001",
			1031 => "0000000001000010001001",
			1032 => "0000001111001000001000",
			1033 => "0011011110000100000100",
			1034 => "0000000001000010001001",
			1035 => "0000001001000010001001",
			1036 => "0000000001000010001001",
			1037 => "0000101000100000001100",
			1038 => "0001101111000000001000",
			1039 => "0001111001001000000100",
			1040 => "0000000001000010001001",
			1041 => "0000000001000010001001",
			1042 => "0000000001000010001001",
			1043 => "0000000001110100010000",
			1044 => "0001110110100100000100",
			1045 => "0000000001000010001001",
			1046 => "0001001110000000001000",
			1047 => "0000011100011000000100",
			1048 => "0000000001000010001001",
			1049 => "0000000001000010001001",
			1050 => "0000000001000010001001",
			1051 => "0001101000010000000100",
			1052 => "0000000001000010001001",
			1053 => "0001000101000000001000",
			1054 => "0010011010100100000100",
			1055 => "0000000001000010001001",
			1056 => "0000000001000010001001",
			1057 => "0000000001000010001001",
			1058 => "0001001000001100110000",
			1059 => "0000011011111100100100",
			1060 => "0000110111010100100000",
			1061 => "0010100000001000010000",
			1062 => "0000111100010000001100",
			1063 => "0000110111100000000100",
			1064 => "0000000001000101001101",
			1065 => "0001011100100100000100",
			1066 => "0000000001000101001101",
			1067 => "0000000001000101001101",
			1068 => "0000000001000101001101",
			1069 => "0001111001001000000100",
			1070 => "0000000001000101001101",
			1071 => "0000011001011000000100",
			1072 => "0000000001000101001101",
			1073 => "0000000101000100000100",
			1074 => "0000000001000101001101",
			1075 => "0000000001000101001101",
			1076 => "0000000001000101001101",
			1077 => "0010110101100100001000",
			1078 => "0010100010101100000100",
			1079 => "0000000001000101001101",
			1080 => "0000000001000101001101",
			1081 => "0000000001000101001101",
			1082 => "0001100100111100100000",
			1083 => "0001001011101100010100",
			1084 => "0010100010101100001100",
			1085 => "0010110100010000001000",
			1086 => "0001011110101000000100",
			1087 => "0000000001000101001101",
			1088 => "0000000001000101001101",
			1089 => "0000000001000101001101",
			1090 => "0000110110111100000100",
			1091 => "0000000001000101001101",
			1092 => "0000000001000101001101",
			1093 => "0010111010010100001000",
			1094 => "0001101001100100000100",
			1095 => "1111111001000101001101",
			1096 => "0000000001000101001101",
			1097 => "0000000001000101001101",
			1098 => "0010011010100000000100",
			1099 => "0000000001000101001101",
			1100 => "0000001010101100001100",
			1101 => "0010111010010100001000",
			1102 => "0010111011011100000100",
			1103 => "0000000001000101001101",
			1104 => "0000000001000101001101",
			1105 => "0000000001000101001101",
			1106 => "0000000001000101001101",
			1107 => "0011000100011000011100",
			1108 => "0011100111010100010000",
			1109 => "0000001001101000001100",
			1110 => "0010100010101100001000",
			1111 => "0010001000010100000100",
			1112 => "0000000001000111111001",
			1113 => "0000000001000111111001",
			1114 => "0000000001000111111001",
			1115 => "1111111001000111111001",
			1116 => "0000000001110100001000",
			1117 => "0010010111101100000100",
			1118 => "0000000001000111111001",
			1119 => "0000000001000111111001",
			1120 => "0000000001000111111001",
			1121 => "0000000010101000111000",
			1122 => "0011101100000000011100",
			1123 => "0001010111100000010000",
			1124 => "0001001100010000000100",
			1125 => "0000000001000111111001",
			1126 => "0010110000011100000100",
			1127 => "0000000001000111111001",
			1128 => "0001010111100000000100",
			1129 => "0000000001000111111001",
			1130 => "0000000001000111111001",
			1131 => "0010100000001000000100",
			1132 => "0000000001000111111001",
			1133 => "0000101100000000000100",
			1134 => "0000000001000111111001",
			1135 => "0000000001000111111001",
			1136 => "0000010000111100001000",
			1137 => "0000111011111000000100",
			1138 => "0000000001000111111001",
			1139 => "0000000001000111111001",
			1140 => "0000011101111100001000",
			1141 => "0000000111000100000100",
			1142 => "0000001001000111111001",
			1143 => "0000000001000111111001",
			1144 => "0001011100100100000100",
			1145 => "0000000001000111111001",
			1146 => "0001010101110000000100",
			1147 => "0000000001000111111001",
			1148 => "0000000001000111111001",
			1149 => "0000000001000111111001",
			1150 => "0011111100000000001100",
			1151 => "0001001100010000000100",
			1152 => "0000000001001010101101",
			1153 => "0010001000100100000100",
			1154 => "0000000001001010101101",
			1155 => "0000000001001010101101",
			1156 => "0001000001011100100000",
			1157 => "0001101101011000010100",
			1158 => "0010110110110100001000",
			1159 => "0001011100100100000100",
			1160 => "0000000001001010101101",
			1161 => "0000000001001010101101",
			1162 => "0000000001010100000100",
			1163 => "0000000001001010101101",
			1164 => "0011010100101000000100",
			1165 => "0000000001001010101101",
			1166 => "0000000001001010101101",
			1167 => "0000001111001000001000",
			1168 => "0011011110000100000100",
			1169 => "0000000001001010101101",
			1170 => "0000000001001010101101",
			1171 => "0000000001001010101101",
			1172 => "0000101000100000010000",
			1173 => "0001101111000000001100",
			1174 => "0001111001001000000100",
			1175 => "0000000001001010101101",
			1176 => "0010110101100100000100",
			1177 => "0000000001001010101101",
			1178 => "0000000001001010101101",
			1179 => "0000000001001010101101",
			1180 => "0000000001110100010000",
			1181 => "0001110110100100000100",
			1182 => "0000000001001010101101",
			1183 => "0001001110000000001000",
			1184 => "0000011100011000000100",
			1185 => "0000000001001010101101",
			1186 => "0000000001001010101101",
			1187 => "0000000001001010101101",
			1188 => "0001101000010000000100",
			1189 => "0000000001001010101101",
			1190 => "0000101011110000001000",
			1191 => "0000011100011000000100",
			1192 => "0000000001001010101101",
			1193 => "0000000001001010101101",
			1194 => "0000000001001010101101",
			1195 => "0000000010101001000100",
			1196 => "0000011001011000010000",
			1197 => "0001100000111100001000",
			1198 => "0010010001000100000100",
			1199 => "1111111001001101001001",
			1200 => "0000001001001101001001",
			1201 => "0010011111000000000100",
			1202 => "1111111001001101001001",
			1203 => "0000000001001101001001",
			1204 => "0011010110010000101100",
			1205 => "0001110110100100010100",
			1206 => "0000001111001000010000",
			1207 => "0011000100011000001000",
			1208 => "0000101100010000000100",
			1209 => "0000000001001101001001",
			1210 => "1111111001001101001001",
			1211 => "0010110100000100000100",
			1212 => "0000000001001101001001",
			1213 => "0000001001001101001001",
			1214 => "1111111001001101001001",
			1215 => "0000111100111000010000",
			1216 => "0000000111000100001000",
			1217 => "0000011101111100000100",
			1218 => "0000001001001101001001",
			1219 => "0000000001001101001001",
			1220 => "0010111011011100000100",
			1221 => "1111111001001101001001",
			1222 => "0000000001001101001001",
			1223 => "0001101000010000000100",
			1224 => "0000001001001101001001",
			1225 => "0000001001001101001001",
			1226 => "0001110101110100000100",
			1227 => "1111111001001101001001",
			1228 => "0000000001001101001001",
			1229 => "0000001010101100001000",
			1230 => "0001101000010000000100",
			1231 => "1111111001001101001001",
			1232 => "0000001001001101001001",
			1233 => "1111111001001101001001",
			1234 => "0000000010101001000000",
			1235 => "0000111100111000110000",
			1236 => "0000001111001000101000",
			1237 => "0001101011001100100000",
			1238 => "0000100111011000010000",
			1239 => "0000011001011000001000",
			1240 => "0000000110011100000100",
			1241 => "0000000001001111010101",
			1242 => "0000000001001111010101",
			1243 => "0010110100010000000100",
			1244 => "0000000001001111010101",
			1245 => "0000000001001111010101",
			1246 => "0011001011000000001000",
			1247 => "0011001010111000000100",
			1248 => "0000000001001111010101",
			1249 => "0000000001001111010101",
			1250 => "0000010001000100000100",
			1251 => "0000000001001111010101",
			1252 => "0000000001001111010101",
			1253 => "0000111010000100000100",
			1254 => "0000000001001111010101",
			1255 => "0000001001001111010101",
			1256 => "0000111000100000000100",
			1257 => "1111111001001111010101",
			1258 => "0000000001001111010101",
			1259 => "0000101101101100000100",
			1260 => "0000001001001111010101",
			1261 => "0011011110010000000100",
			1262 => "0000000001001111010101",
			1263 => "0000100011000000000100",
			1264 => "0000000001001111010101",
			1265 => "0000000001001111010101",
			1266 => "0010010010101100000100",
			1267 => "1111111001001111010101",
			1268 => "0000000001001111010101",
			1269 => "0001001011110000111100",
			1270 => "0010011111000000010000",
			1271 => "0011100010000100001100",
			1272 => "0001100000111100001000",
			1273 => "0001100000111100000100",
			1274 => "1111111001010010111001",
			1275 => "0000001001010010111001",
			1276 => "1111111001010010111001",
			1277 => "0000001001010010111001",
			1278 => "0011011110000100001100",
			1279 => "0000011011111100001000",
			1280 => "0001000111010100000100",
			1281 => "0000010001010010111001",
			1282 => "1111111001010010111001",
			1283 => "1111111001010010111001",
			1284 => "0000010100110100011000",
			1285 => "0010100000001000001000",
			1286 => "0001011100100100000100",
			1287 => "0000001001010010111001",
			1288 => "1111111001010010111001",
			1289 => "0001000110111000001000",
			1290 => "0000011001011000000100",
			1291 => "0000000001010010111001",
			1292 => "0000010001010010111001",
			1293 => "0000111100111000000100",
			1294 => "1111111001010010111001",
			1295 => "0000100001010010111001",
			1296 => "0011001011000000000100",
			1297 => "0000000001010010111001",
			1298 => "1111111001010010111001",
			1299 => "0001001000110100011000",
			1300 => "0001101000010000010000",
			1301 => "0001101000010000001000",
			1302 => "0001001110000000000100",
			1303 => "1111111001010010111001",
			1304 => "1111111001010010111001",
			1305 => "0001001000000100000100",
			1306 => "0000000001010010111001",
			1307 => "1111111001010010111001",
			1308 => "0000111000101000000100",
			1309 => "1111111001010010111001",
			1310 => "0000011001010010111001",
			1311 => "0001000101000000011100",
			1312 => "0001000101000000010000",
			1313 => "0010000001110000000100",
			1314 => "1111111001010010111001",
			1315 => "0010001100000100001000",
			1316 => "0010000001110000000100",
			1317 => "0000000001010010111001",
			1318 => "0000000001010010111001",
			1319 => "1111111001010010111001",
			1320 => "0010000001110000000100",
			1321 => "1111111001010010111001",
			1322 => "0000011101111100000100",
			1323 => "1111111001010010111001",
			1324 => "0000010001010010111001",
			1325 => "1111111001010010111001",
			1326 => "0000000111000101000100",
			1327 => "0000110110111100011100",
			1328 => "0010011111000000001100",
			1329 => "0010011111000000000100",
			1330 => "1100101001010110101101",
			1331 => "0010100000001000000100",
			1332 => "1100101001010110101101",
			1333 => "1101010001010110101101",
			1334 => "0000001100000100001000",
			1335 => "0011001000000000000100",
			1336 => "1111011001010110101101",
			1337 => "1110011001010110101101",
			1338 => "0011010101001000000100",
			1339 => "1100101001010110101101",
			1340 => "1101111001010110101101",
			1341 => "0011010101001000001000",
			1342 => "0011011110000100000100",
			1343 => "1100101001010110101101",
			1344 => "1101011001010110101101",
			1345 => "0010011111000000010000",
			1346 => "0001100100110100001000",
			1347 => "0010001000100100000100",
			1348 => "1100101001010110101101",
			1349 => "1101010001010110101101",
			1350 => "0001111000011000000100",
			1351 => "1101000001010110101101",
			1352 => "1110100001010110101101",
			1353 => "0000010100110100001100",
			1354 => "0001000110111000001000",
			1355 => "0010001000100100000100",
			1356 => "1110100001010110101101",
			1357 => "1111010001010110101101",
			1358 => "1110000001010110101101",
			1359 => "1100101001010110101101",
			1360 => "0000000001110100011000",
			1361 => "0010000101000100010100",
			1362 => "0001100100111100001100",
			1363 => "0001100100111100000100",
			1364 => "1100101001010110101101",
			1365 => "0001001011110000000100",
			1366 => "1100111001010110101101",
			1367 => "1100101001010110101101",
			1368 => "0000011010011000000100",
			1369 => "1101011001010110101101",
			1370 => "1100101001010110101101",
			1371 => "1110101001010110101101",
			1372 => "0000001010101100011000",
			1373 => "0001101000010000010100",
			1374 => "0010000001010100001100",
			1375 => "0010000001010100000100",
			1376 => "1100101001010110101101",
			1377 => "0001001000000100000100",
			1378 => "1100111001010110101101",
			1379 => "1100101001010110101101",
			1380 => "0000011010011000000100",
			1381 => "1101101001010110101101",
			1382 => "1100101001010110101101",
			1383 => "1110111001010110101101",
			1384 => "0000001010101100000100",
			1385 => "1100101001010110101101",
			1386 => "1100101001010110101101",
			1387 => "0010010111101101010000",
			1388 => "0000001001101000111100",
			1389 => "0001011100100100011000",
			1390 => "0010001000100100010000",
			1391 => "0010011000010000001100",
			1392 => "0011000100011000000100",
			1393 => "0000000001011010101001",
			1394 => "0000111100000000000100",
			1395 => "0000000001011010101001",
			1396 => "0000000001011010101001",
			1397 => "0000000001011010101001",
			1398 => "0001010110100000000100",
			1399 => "0000000001011010101001",
			1400 => "0000000001011010101001",
			1401 => "0001010111100000001100",
			1402 => "0011111111010100001000",
			1403 => "0001100100110100000100",
			1404 => "0000000001011010101001",
			1405 => "0000000001011010101001",
			1406 => "0000000001011010101001",
			1407 => "0000010000111100010000",
			1408 => "0000111111010100001000",
			1409 => "0010011111000000000100",
			1410 => "0000000001011010101001",
			1411 => "0000000001011010101001",
			1412 => "0001111111011100000100",
			1413 => "0000000001011010101001",
			1414 => "0000000001011010101001",
			1415 => "0010000110011000000100",
			1416 => "0000000001011010101001",
			1417 => "0000000001011010101001",
			1418 => "0011000100011000001000",
			1419 => "0000010001111000000100",
			1420 => "1111111001011010101001",
			1421 => "0000000001011010101001",
			1422 => "0000010001000100000100",
			1423 => "0000000001011010101001",
			1424 => "0010010100101100000100",
			1425 => "0000000001011010101001",
			1426 => "0000000001011010101001",
			1427 => "0000000111000100010000",
			1428 => "0001101011001100000100",
			1429 => "0000000001011010101001",
			1430 => "0000110111010100000100",
			1431 => "0000000001011010101001",
			1432 => "0001011001010000000100",
			1433 => "0000001001011010101001",
			1434 => "0000000001011010101001",
			1435 => "0011101100111000001100",
			1436 => "0011000100011000000100",
			1437 => "0000000001011010101001",
			1438 => "0000110011000000000100",
			1439 => "0000000001011010101001",
			1440 => "0000000001011010101001",
			1441 => "0011111110000000010000",
			1442 => "0001101000010000000100",
			1443 => "0000000001011010101001",
			1444 => "0001010001000000000100",
			1445 => "0000000001011010101001",
			1446 => "0010101001000100000100",
			1447 => "0000000001011010101001",
			1448 => "0000000001011010101001",
			1449 => "0000000001011010101001",
			1450 => "0011001010111000001100",
			1451 => "0011100111010100001000",
			1452 => "0001011101000100000100",
			1453 => "0000000001011101110101",
			1454 => "0000000001011101110101",
			1455 => "0000000001011101110101",
			1456 => "0011001000000000110000",
			1457 => "0001010101001000100000",
			1458 => "0010010111101100001100",
			1459 => "0000000110001000001000",
			1460 => "0001111111011100000100",
			1461 => "0000000001011101110101",
			1462 => "0000000001011101110101",
			1463 => "0000000001011101110101",
			1464 => "0001101011001100001000",
			1465 => "0010010000001000000100",
			1466 => "0000000001011101110101",
			1467 => "0000000001011101110101",
			1468 => "0000000001110100001000",
			1469 => "0001100100111100000100",
			1470 => "0000000001011101110101",
			1471 => "0000000001011101110101",
			1472 => "0000000001011101110101",
			1473 => "0010010101010000001000",
			1474 => "0000111010000100000100",
			1475 => "0000000001011101110101",
			1476 => "0000000001011101110101",
			1477 => "0000001010101100000100",
			1478 => "0000000001011101110101",
			1479 => "0000000001011101110101",
			1480 => "0001011110000100001000",
			1481 => "0001111000011000000100",
			1482 => "0000000001011101110101",
			1483 => "0000000001011101110101",
			1484 => "0011001001110100010100",
			1485 => "0011001001001000001100",
			1486 => "0001010010011100001000",
			1487 => "0011011010001000000100",
			1488 => "0000000001011101110101",
			1489 => "0000000001011101110101",
			1490 => "0000000001011101110101",
			1491 => "0000101000101000000100",
			1492 => "0000000001011101110101",
			1493 => "0000000001011101110101",
			1494 => "0000100010010100001100",
			1495 => "0011110111011000000100",
			1496 => "0000000001011101110101",
			1497 => "0001001000110100000100",
			1498 => "0000000001011101110101",
			1499 => "0000000001011101110101",
			1500 => "0000000001011101110101",
			1501 => "0011000100011000100100",
			1502 => "0001001010000100001100",
			1503 => "0011101110101100000100",
			1504 => "0000000001100001110001",
			1505 => "0000101110110100000100",
			1506 => "0000000001100001110001",
			1507 => "0000000001100001110001",
			1508 => "0010010000001000001100",
			1509 => "0000001001101000001000",
			1510 => "0000001100000100000100",
			1511 => "0000000001100001110001",
			1512 => "0000000001100001110001",
			1513 => "1111111001100001110001",
			1514 => "0000000001110100001000",
			1515 => "0011100111010100000100",
			1516 => "0000000001100001110001",
			1517 => "0000000001100001110001",
			1518 => "0000000001100001110001",
			1519 => "0001101101111100011000",
			1520 => "0000101110110100010000",
			1521 => "0000111100000000001100",
			1522 => "0000110010000000000100",
			1523 => "0000000001100001110001",
			1524 => "0011010010011100000100",
			1525 => "0000000001100001110001",
			1526 => "0000000001100001110001",
			1527 => "0000000001100001110001",
			1528 => "0011010111111100000100",
			1529 => "0000000001100001110001",
			1530 => "0000000001100001110001",
			1531 => "0011000100011000010000",
			1532 => "0001100100111100001100",
			1533 => "0000000001110100001000",
			1534 => "0011010001000000000100",
			1535 => "0000000001100001110001",
			1536 => "0000000001100001110001",
			1537 => "0000000001100001110001",
			1538 => "0000000001100001110001",
			1539 => "0001010111100000010100",
			1540 => "0010010101010000001000",
			1541 => "0010011111000000000100",
			1542 => "0000000001100001110001",
			1543 => "0000000001100001110001",
			1544 => "0010100010101100000100",
			1545 => "1111111001100001110001",
			1546 => "0010010000001000000100",
			1547 => "0000000001100001110001",
			1548 => "0000000001100001110001",
			1549 => "0000010101011100010000",
			1550 => "0001101010011000001000",
			1551 => "0011001001110100000100",
			1552 => "0000000001100001110001",
			1553 => "0000000001100001110001",
			1554 => "0000111000100000000100",
			1555 => "0000000001100001110001",
			1556 => "0000000001100001110001",
			1557 => "0000000001110100001000",
			1558 => "0000110010010100000100",
			1559 => "0000000001100001110001",
			1560 => "0000000001100001110001",
			1561 => "0011101101101100000100",
			1562 => "0000000001100001110001",
			1563 => "0000000001100001110001",
			1564 => "0011001010111000011000",
			1565 => "0000000110001000010100",
			1566 => "0000100111011000001100",
			1567 => "0011001010111000001000",
			1568 => "0001110110100100000100",
			1569 => "0000000001100101011101",
			1570 => "0000000001100101011101",
			1571 => "0000000001100101011101",
			1572 => "0011010101001000000100",
			1573 => "0000000001100101011101",
			1574 => "0000000001100101011101",
			1575 => "1111111001100101011101",
			1576 => "0011001011000000111000",
			1577 => "0001010101001000101100",
			1578 => "0000011101111100100000",
			1579 => "0011011111010000010000",
			1580 => "0001010010110100001000",
			1581 => "0000001011010100000100",
			1582 => "0000000001100101011101",
			1583 => "0000000001100101011101",
			1584 => "0001010110100000000100",
			1585 => "1111111001100101011101",
			1586 => "0000000001100101011101",
			1587 => "0011010100101000001000",
			1588 => "0001101101111100000100",
			1589 => "0000000001100101011101",
			1590 => "0000001001100101011101",
			1591 => "0001010111100000000100",
			1592 => "0000000001100101011101",
			1593 => "0000000001100101011101",
			1594 => "0011010100101000001000",
			1595 => "0011000100011000000100",
			1596 => "0000000001100101011101",
			1597 => "0000000001100101011101",
			1598 => "0000000001100101011101",
			1599 => "0000111010000100000100",
			1600 => "0000000001100101011101",
			1601 => "0010010101010000000100",
			1602 => "1111111001100101011101",
			1603 => "0000000001100101011101",
			1604 => "0000101110110100001100",
			1605 => "0000010000111100001000",
			1606 => "0001000010000100000100",
			1607 => "0000000001100101011101",
			1608 => "0000000001100101011101",
			1609 => "0000000001100101011101",
			1610 => "0011000110100100010000",
			1611 => "0010010011101000001100",
			1612 => "0000011001011000000100",
			1613 => "0000000001100101011101",
			1614 => "0000001010101100000100",
			1615 => "0000001001100101011101",
			1616 => "0000000001100101011101",
			1617 => "0000000001100101011101",
			1618 => "0010001100011100001000",
			1619 => "0001111111011100000100",
			1620 => "0000000001100101011101",
			1621 => "0000000001100101011101",
			1622 => "0000000001100101011101",
			1623 => "0010010111101101010000",
			1624 => "0001001111100101000000",
			1625 => "0001011100100100100000",
			1626 => "0011011111010000010100",
			1627 => "0000011011111100001000",
			1628 => "0011001010111000000100",
			1629 => "0000000001101001101001",
			1630 => "0000000001101001101001",
			1631 => "0010100010101100001000",
			1632 => "0011001010111000000100",
			1633 => "0000000001101001101001",
			1634 => "0000000001101001101001",
			1635 => "0000000001101001101001",
			1636 => "0001101101111100000100",
			1637 => "0000000001101001101001",
			1638 => "0000100010000000000100",
			1639 => "0000000001101001101001",
			1640 => "0000000001101001101001",
			1641 => "0001110001101000001100",
			1642 => "0001101010011000001000",
			1643 => "0000111100000000000100",
			1644 => "0000000001101001101001",
			1645 => "0000000001101001101001",
			1646 => "0000000001101001101001",
			1647 => "0001111000011000001000",
			1648 => "0000100010000100000100",
			1649 => "0000000001101001101001",
			1650 => "0000000001101001101001",
			1651 => "0000110110111100000100",
			1652 => "0000000001101001101001",
			1653 => "0001111111011100000100",
			1654 => "0000000001101001101001",
			1655 => "0000000001101001101001",
			1656 => "0011000110100100001100",
			1657 => "0010010111101100001000",
			1658 => "0010000110011000000100",
			1659 => "0000000001101001101001",
			1660 => "1111111001101001101001",
			1661 => "0000000001101001101001",
			1662 => "0000000001101001101001",
			1663 => "0001110001101000011000",
			1664 => "0001101011001100000100",
			1665 => "0000000001101001101001",
			1666 => "0000101101101100010000",
			1667 => "0000111000001100000100",
			1668 => "0000000001101001101001",
			1669 => "0010101000100100001000",
			1670 => "0011010101001000000100",
			1671 => "0000000001101001101001",
			1672 => "0000000001101001101001",
			1673 => "0000000001101001101001",
			1674 => "0000000001101001101001",
			1675 => "0011101100111000001100",
			1676 => "0001001011101100000100",
			1677 => "0000000001101001101001",
			1678 => "0000110011000000000100",
			1679 => "0000000001101001101001",
			1680 => "0000000001101001101001",
			1681 => "0011111110000000010000",
			1682 => "0001011110000100000100",
			1683 => "0000000001101001101001",
			1684 => "0001110000011100001000",
			1685 => "0011000110100100000100",
			1686 => "0000000001101001101001",
			1687 => "0000000001101001101001",
			1688 => "0000000001101001101001",
			1689 => "0000000001101001101001",
			1690 => "0000001010101101000000",
			1691 => "0011000111001000001100",
			1692 => "0001110110100100000100",
			1693 => "1111111001101011101101",
			1694 => "0001101101111100000100",
			1695 => "0000000001101011101101",
			1696 => "0000000001101011101101",
			1697 => "0010101000010100110000",
			1698 => "0000001111001000011100",
			1699 => "0001101101011000010000",
			1700 => "0000001001101000001000",
			1701 => "0010110100010000000100",
			1702 => "0000000001101011101101",
			1703 => "0000001001101011101101",
			1704 => "0011001011000000000100",
			1705 => "1111111001101011101101",
			1706 => "0000000001101011101101",
			1707 => "0011101111010100001000",
			1708 => "0000010111101000000100",
			1709 => "0000001001101011101101",
			1710 => "1111111001101011101101",
			1711 => "0000001001101011101101",
			1712 => "0000111111100100000100",
			1713 => "1111111001101011101101",
			1714 => "0000010100110100001000",
			1715 => "0000000010101000000100",
			1716 => "0000001001101011101101",
			1717 => "0000000001101011101101",
			1718 => "0010101000010100000100",
			1719 => "1111111001101011101101",
			1720 => "0000000001101011101101",
			1721 => "0000010001101011101101",
			1722 => "1111111001101011101101",
			1723 => "0011001010111000001000",
			1724 => "0000000110001000000100",
			1725 => "0000000001101110111001",
			1726 => "0000000001101110111001",
			1727 => "0011001000000000110000",
			1728 => "0010110101110100101000",
			1729 => "0001110110100100011000",
			1730 => "0001111001001000001100",
			1731 => "0000001111001000001000",
			1732 => "0001111011000000000100",
			1733 => "0000000001101110111001",
			1734 => "0000000001101110111001",
			1735 => "0000000001101110111001",
			1736 => "0010100010101100001000",
			1737 => "0011111100010000000100",
			1738 => "0000000001101110111001",
			1739 => "0000000001101110111001",
			1740 => "0000000001101110111001",
			1741 => "0000000010101000001100",
			1742 => "0001101101111100000100",
			1743 => "0000000001101110111001",
			1744 => "0000011001011000000100",
			1745 => "0000000001101110111001",
			1746 => "0000001001101110111001",
			1747 => "0000000001101110111001",
			1748 => "0010010101010000000100",
			1749 => "0000000001101110111001",
			1750 => "0000000001101110111001",
			1751 => "0010110100010000001100",
			1752 => "0001101000010000001000",
			1753 => "0011001001110100000100",
			1754 => "0000000001101110111001",
			1755 => "0000000001101110111001",
			1756 => "0000000001101110111001",
			1757 => "0011011100010100010000",
			1758 => "0001111000011000000100",
			1759 => "0000000001101110111001",
			1760 => "0011000001101000001000",
			1761 => "0000001000101100000100",
			1762 => "0000000001101110111001",
			1763 => "0000000001101110111001",
			1764 => "0000000001101110111001",
			1765 => "0001110000011100001000",
			1766 => "0010010010101100000100",
			1767 => "0000000001101110111001",
			1768 => "0000000001101110111001",
			1769 => "0000010111101000001000",
			1770 => "0010111110101100000100",
			1771 => "0000000001101110111001",
			1772 => "0000000001101110111001",
			1773 => "0000000001101110111001",
			1774 => "0000001010101101000100",
			1775 => "0011000111001000001100",
			1776 => "0001110110100100000100",
			1777 => "1111111001110001000101",
			1778 => "0001101101111100000100",
			1779 => "0000000001110001000101",
			1780 => "0000000001110001000101",
			1781 => "0010101000010100110100",
			1782 => "0011010011001000100000",
			1783 => "0010110110110100010000",
			1784 => "0000001111001000001000",
			1785 => "0011010101110000000100",
			1786 => "0000001001110001000101",
			1787 => "0000000001110001000101",
			1788 => "0011010101110000000100",
			1789 => "1111111001110001000101",
			1790 => "0000001001110001000101",
			1791 => "0000000101000100001000",
			1792 => "0001100100110100000100",
			1793 => "1111111001110001000101",
			1794 => "0000000001110001000101",
			1795 => "0000111010000100000100",
			1796 => "0000001001110001000101",
			1797 => "0000000001110001000101",
			1798 => "0001001101101100001000",
			1799 => "0001111111011100000100",
			1800 => "0000000001110001000101",
			1801 => "0000001001110001000101",
			1802 => "0001110101110100001000",
			1803 => "0010101000010100000100",
			1804 => "1111111001110001000101",
			1805 => "0000000001110001000101",
			1806 => "0000000001110001000101",
			1807 => "0000010001110001000101",
			1808 => "1111111001110001000101",
			1809 => "0001110110100100010000",
			1810 => "0000000001010100000100",
			1811 => "0000000001110100111001",
			1812 => "0000110111010100001000",
			1813 => "0011001011000000000100",
			1814 => "1111111001110100111001",
			1815 => "0000000001110100111001",
			1816 => "0000000001110100111001",
			1817 => "0001111000011001001000",
			1818 => "0001011100100100100100",
			1819 => "0011100110010000001000",
			1820 => "0000011011111100000100",
			1821 => "0000000001110100111001",
			1822 => "0000000001110100111001",
			1823 => "0000010111101000001100",
			1824 => "0000000110001000001000",
			1825 => "0010100000001000000100",
			1826 => "0000000001110100111001",
			1827 => "0000000001110100111001",
			1828 => "0000000001110100111001",
			1829 => "0000110000010000001000",
			1830 => "0001001011101100000100",
			1831 => "0000000001110100111001",
			1832 => "0000000001110100111001",
			1833 => "0010101000100100000100",
			1834 => "0000000001110100111001",
			1835 => "0000000001110100111001",
			1836 => "0011110111011000010100",
			1837 => "0011100010000100001100",
			1838 => "0010100000001000001000",
			1839 => "0000111100010000000100",
			1840 => "0000000001110100111001",
			1841 => "0000000001110100111001",
			1842 => "0000000001110100111001",
			1843 => "0000111010000100000100",
			1844 => "0000000001110100111001",
			1845 => "0000000001110100111001",
			1846 => "0011001001110100001100",
			1847 => "0011001010111000000100",
			1848 => "0000000001110100111001",
			1849 => "0001110110100100000100",
			1850 => "0000000001110100111001",
			1851 => "0000000001110100111001",
			1852 => "0000000001110100111001",
			1853 => "0000111000100000010000",
			1854 => "0000000101000100000100",
			1855 => "0000000001110100111001",
			1856 => "0001000011000000001000",
			1857 => "0001111000011000000100",
			1858 => "0000000001110100111001",
			1859 => "0000001001110100111001",
			1860 => "0000000001110100111001",
			1861 => "0000010001000100000100",
			1862 => "0000000001110100111001",
			1863 => "0000100010010100001100",
			1864 => "0000011010011000001000",
			1865 => "0000110001011100000100",
			1866 => "0000000001110100111001",
			1867 => "0000000001110100111001",
			1868 => "0000000001110100111001",
			1869 => "0000000001110100111001",
			1870 => "0001110110100100010000",
			1871 => "0001001010000100000100",
			1872 => "0000000001111000110101",
			1873 => "0000100110111100001000",
			1874 => "0011000100011000000100",
			1875 => "1111111001111000110101",
			1876 => "0000000001111000110101",
			1877 => "0000000001111000110101",
			1878 => "0001101101011001000000",
			1879 => "0001000110101100110000",
			1880 => "0010101010100000011100",
			1881 => "0000011001011000001100",
			1882 => "0001101101111100001000",
			1883 => "0011001011000000000100",
			1884 => "0000000001111000110101",
			1885 => "0000000001111000110101",
			1886 => "0000000001111000110101",
			1887 => "0001100100110100001000",
			1888 => "0011100010000000000100",
			1889 => "0000000001111000110101",
			1890 => "0000000001111000110101",
			1891 => "0000111100010000000100",
			1892 => "0000000001111000110101",
			1893 => "0000000001111000110101",
			1894 => "0010110101100100001100",
			1895 => "0011110110111100001000",
			1896 => "0000010101011100000100",
			1897 => "0000000001111000110101",
			1898 => "0000000001111000110101",
			1899 => "0000000001111000110101",
			1900 => "0000010000111100000100",
			1901 => "0000000001111000110101",
			1902 => "0000000001111000110101",
			1903 => "0001110111010000001100",
			1904 => "0001011100100100000100",
			1905 => "0000000001111000110101",
			1906 => "0011001001110100000100",
			1907 => "1111111001111000110101",
			1908 => "0000000001111000110101",
			1909 => "0000000001111000110101",
			1910 => "0000001111001000010000",
			1911 => "0000011101111100001100",
			1912 => "0011000100011000000100",
			1913 => "0000000001111000110101",
			1914 => "0000110110111100000100",
			1915 => "0000000001111000110101",
			1916 => "0000001001111000110101",
			1917 => "0000000001111000110101",
			1918 => "0000011101111100001000",
			1919 => "0011001011011100000100",
			1920 => "0000000001111000110101",
			1921 => "0000000001111000110101",
			1922 => "0000010100110100001100",
			1923 => "0010101000010100001000",
			1924 => "0001011110101000000100",
			1925 => "0000000001111000110101",
			1926 => "0000000001111000110101",
			1927 => "0000000001111000110101",
			1928 => "0010101000010100000100",
			1929 => "0000000001111000110101",
			1930 => "0001000101000000000100",
			1931 => "0000000001111000110101",
			1932 => "0000000001111000110101",
			1933 => "0010011111000000010000",
			1934 => "0010000100101100001100",
			1935 => "0001000111010000000100",
			1936 => "0000000001111100010001",
			1937 => "0010101001100100000100",
			1938 => "0000000001111100010001",
			1939 => "0000000001111100010001",
			1940 => "1111111001111100010001",
			1941 => "0011000001101001010100",
			1942 => "0011000100011000110000",
			1943 => "0001010111100000011100",
			1944 => "0010011010100000010000",
			1945 => "0001110110100100001000",
			1946 => "0010101010100100000100",
			1947 => "0000000001111100010001",
			1948 => "1111111001111100010001",
			1949 => "0010110110110100000100",
			1950 => "0000001001111100010001",
			1951 => "0000000001111100010001",
			1952 => "0010111011011100000100",
			1953 => "1111111001111100010001",
			1954 => "0000010100110100000100",
			1955 => "0000000001111100010001",
			1956 => "0000000001111100010001",
			1957 => "0010110010001000010000",
			1958 => "0001101001100100001000",
			1959 => "0011100010000100000100",
			1960 => "0000000001111100010001",
			1961 => "1111111001111100010001",
			1962 => "0000010100110100000100",
			1963 => "0000000001111100010001",
			1964 => "0000000001111100010001",
			1965 => "0000000001111100010001",
			1966 => "0000011001011000001000",
			1967 => "0000110110111100000100",
			1968 => "0000001001111100010001",
			1969 => "0000000001111100010001",
			1970 => "0001100100110100001100",
			1971 => "0010011111000000000100",
			1972 => "0000000001111100010001",
			1973 => "0010010100111100000100",
			1974 => "1111111001111100010001",
			1975 => "0000000001111100010001",
			1976 => "0000101100010000001000",
			1977 => "0000011110010100000100",
			1978 => "0000001001111100010001",
			1979 => "0000000001111100010001",
			1980 => "0011101100000000000100",
			1981 => "1111111001111100010001",
			1982 => "0000000001111100010001",
			1983 => "0010011000010000000100",
			1984 => "1111101001111100010001",
			1985 => "0000101101101100000100",
			1986 => "0000000001111100010001",
			1987 => "1111111001111100010001",
			1988 => "0011001010111000010000",
			1989 => "0000000110001000001100",
			1990 => "0010110000011100000100",
			1991 => "0000000010000000010101",
			1992 => "0010000111110100000100",
			1993 => "0000000010000000010101",
			1994 => "0000000010000000010101",
			1995 => "1111111010000000010101",
			1996 => "0000100111011000110000",
			1997 => "0000011011111100100100",
			1998 => "0000111111010100011000",
			1999 => "0000000101000100001100",
			2000 => "0010110110110100001000",
			2001 => "0001001100010000000100",
			2002 => "0000000010000000010101",
			2003 => "0000000010000000010101",
			2004 => "0000000010000000010101",
			2005 => "0010100000001000000100",
			2006 => "0000000010000000010101",
			2007 => "0010011001100100000100",
			2008 => "0000000010000000010101",
			2009 => "0000001010000000010101",
			2010 => "0010001000100100001000",
			2011 => "0000000001010100000100",
			2012 => "0000000010000000010101",
			2013 => "0000000010000000010101",
			2014 => "0000000010000000010101",
			2015 => "0011100110010000000100",
			2016 => "1111111010000000010101",
			2017 => "0000110111011000000100",
			2018 => "0000000010000000010101",
			2019 => "0000000010000000010101",
			2020 => "0011100111010100101100",
			2021 => "0001001111100100011000",
			2022 => "0010100010101100010000",
			2023 => "0001111111011100001000",
			2024 => "0011111111010100000100",
			2025 => "0000000010000000010101",
			2026 => "1111111010000000010101",
			2027 => "0010110100010000000100",
			2028 => "0000000010000000010101",
			2029 => "0000000010000000010101",
			2030 => "0010010111101100000100",
			2031 => "0000001010000000010101",
			2032 => "0000000010000000010101",
			2033 => "0000110000010000001100",
			2034 => "0011001010111000000100",
			2035 => "0000000010000000010101",
			2036 => "0001101001100100000100",
			2037 => "1111111010000000010101",
			2038 => "0000000010000000010101",
			2039 => "0001101001100100000100",
			2040 => "0000000010000000010101",
			2041 => "0000000010000000010101",
			2042 => "0001000001011100000100",
			2043 => "0000001010000000010101",
			2044 => "0000111000100000000100",
			2045 => "1111111010000000010101",
			2046 => "0010110101110100001000",
			2047 => "0000010100110100000100",
			2048 => "0000001010000000010101",
			2049 => "0000000010000000010101",
			2050 => "0001110101110100000100",
			2051 => "0000000010000000010101",
			2052 => "0000000010000000010101",
			2053 => "0010011111000000001000",
			2054 => "0001100000111100000100",
			2055 => "0000000010000100001001",
			2056 => "1111111010000100001001",
			2057 => "0010010111101101001000",
			2058 => "0000001100000100101000",
			2059 => "0000000001010100011000",
			2060 => "0011010101110000001000",
			2061 => "0011010010011100000100",
			2062 => "0000001010000100001001",
			2063 => "0000000010000100001001",
			2064 => "0011111100000000001000",
			2065 => "0010001000100100000100",
			2066 => "1111111010000100001001",
			2067 => "0000000010000100001001",
			2068 => "0000101100010000000100",
			2069 => "0000000010000100001001",
			2070 => "0000000010000100001001",
			2071 => "0000100010000000000100",
			2072 => "0000000010000100001001",
			2073 => "0011111000001100001000",
			2074 => "0001110110100100000100",
			2075 => "0000000010000100001001",
			2076 => "0000001010000100001001",
			2077 => "0000000010000100001001",
			2078 => "0011001000011000011000",
			2079 => "0001001101101100010000",
			2080 => "0010111011011100001000",
			2081 => "0010100010101100000100",
			2082 => "1111111010000100001001",
			2083 => "0000000010000100001001",
			2084 => "0000010101011100000100",
			2085 => "0000000010000100001001",
			2086 => "0000000010000100001001",
			2087 => "0011000110100100000100",
			2088 => "1111111010000100001001",
			2089 => "0000000010000100001001",
			2090 => "0001000110001100000100",
			2091 => "0000000010000100001001",
			2092 => "0000000010000100001001",
			2093 => "0000000001110100010100",
			2094 => "0001101011001100001000",
			2095 => "0010010111101100000100",
			2096 => "0000000010000100001001",
			2097 => "0000000010000100001001",
			2098 => "0011101111010100000100",
			2099 => "0000000010000100001001",
			2100 => "0001110000011100000100",
			2101 => "0000001010000100001001",
			2102 => "0000000010000100001001",
			2103 => "0011101100111000000100",
			2104 => "1111111010000100001001",
			2105 => "0001101000010000001000",
			2106 => "0010101000100100000100",
			2107 => "0000000010000100001001",
			2108 => "0000000010000100001001",
			2109 => "0011111110000000001000",
			2110 => "0010111011110100000100",
			2111 => "0000000010000100001001",
			2112 => "0000000010000100001001",
			2113 => "0000000010000100001001",
			2114 => "0000001010101101110000",
			2115 => "0001111000011001001100",
			2116 => "0001111000011000111000",
			2117 => "0001011100100100011000",
			2118 => "0000010111101000001100",
			2119 => "0000111010000100001000",
			2120 => "0000011011111100000100",
			2121 => "0000000010000111101101",
			2122 => "1111111010000111101101",
			2123 => "0000001010000111101101",
			2124 => "0001011101000100000100",
			2125 => "1111111010000111101101",
			2126 => "0011000100011000000100",
			2127 => "0000000010000111101101",
			2128 => "0000000010000111101101",
			2129 => "0011000100011000010000",
			2130 => "0001011100100100001000",
			2131 => "0000010000111100000100",
			2132 => "0000000010000111101101",
			2133 => "0000000010000111101101",
			2134 => "0011010010011100000100",
			2135 => "0000000010000111101101",
			2136 => "1111111010000111101101",
			2137 => "0000010000111100001000",
			2138 => "0001011111010000000100",
			2139 => "0000000010000111101101",
			2140 => "1111111010000111101101",
			2141 => "0000000001110100000100",
			2142 => "0000001010000111101101",
			2143 => "0000000010000111101101",
			2144 => "0001100100110100000100",
			2145 => "0000000010000111101101",
			2146 => "0001101011001100001000",
			2147 => "0000111111010100000100",
			2148 => "0000000010000111101101",
			2149 => "1111111010000111101101",
			2150 => "0010010000001000000100",
			2151 => "0000000010000111101101",
			2152 => "0000000010000111101101",
			2153 => "0011000001101000011000",
			2154 => "0011011100010100010000",
			2155 => "0000000101000100000100",
			2156 => "0000000010000111101101",
			2157 => "0010110100010000001000",
			2158 => "0010110010001000000100",
			2159 => "0000001010000111101101",
			2160 => "0000000010000111101101",
			2161 => "0000001010000111101101",
			2162 => "0001010011001000000100",
			2163 => "0000000010000111101101",
			2164 => "0000000010000111101101",
			2165 => "0010010101010000000100",
			2166 => "1111111010000111101101",
			2167 => "0000010100110100000100",
			2168 => "0000000010000111101101",
			2169 => "0000000010000111101101",
			2170 => "1111111010000111101101",
			2171 => "0011000111001000001000",
			2172 => "0001110110100100000100",
			2173 => "1111111010001011101001",
			2174 => "0000000010001011101001",
			2175 => "0001101101111100100000",
			2176 => "0011010111111100011100",
			2177 => "0010111011011100001100",
			2178 => "0011000100011000000100",
			2179 => "0000000010001011101001",
			2180 => "0011010010011100000100",
			2181 => "0000000010001011101001",
			2182 => "0000000010001011101001",
			2183 => "0001110001101000001000",
			2184 => "0011010010011100000100",
			2185 => "0000000010001011101001",
			2186 => "0000000010001011101001",
			2187 => "0000011001011000000100",
			2188 => "0000000010001011101001",
			2189 => "0000000010001011101001",
			2190 => "0000001010001011101001",
			2191 => "0001011100100100101000",
			2192 => "0000010111101000010100",
			2193 => "0011100111011000010000",
			2194 => "0000011011111100001000",
			2195 => "0010001100011100000100",
			2196 => "0000001010001011101001",
			2197 => "0000000010001011101001",
			2198 => "0011000100011000000100",
			2199 => "0000000010001011101001",
			2200 => "1111111010001011101001",
			2201 => "0000001010001011101001",
			2202 => "0011010010011100001100",
			2203 => "0001111001001000000100",
			2204 => "0000000010001011101001",
			2205 => "0010100011101000000100",
			2206 => "0000000010001011101001",
			2207 => "1111111010001011101001",
			2208 => "0010101000010100000100",
			2209 => "0000000010001011101001",
			2210 => "0000000010001011101001",
			2211 => "0001011100100100010100",
			2212 => "0000010100110100001100",
			2213 => "0011010100101000001000",
			2214 => "0000101101101100000100",
			2215 => "0000001010001011101001",
			2216 => "0000000010001011101001",
			2217 => "0000000010001011101001",
			2218 => "0001110001101000000100",
			2219 => "0000000010001011101001",
			2220 => "0000000010001011101001",
			2221 => "0011000110100100010000",
			2222 => "0001111000011000001000",
			2223 => "0001111000011000000100",
			2224 => "0000000010001011101001",
			2225 => "0000000010001011101001",
			2226 => "0011011100010100000100",
			2227 => "0000001010001011101001",
			2228 => "0000000010001011101001",
			2229 => "0010110101110100000100",
			2230 => "1111111010001011101001",
			2231 => "0001101001100100000100",
			2232 => "0000000010001011101001",
			2233 => "0000000010001011101001",
			2234 => "0011000111001000001000",
			2235 => "0001110110100100000100",
			2236 => "1111111010001111010101",
			2237 => "0000000010001111010101",
			2238 => "0011000001101001100000",
			2239 => "0011001011000000110100",
			2240 => "0001110001101000011100",
			2241 => "0001110110100100010000",
			2242 => "0001111001001000001000",
			2243 => "0000001111001000000100",
			2244 => "0000000010001111010101",
			2245 => "0000000010001111010101",
			2246 => "0010100010101100000100",
			2247 => "1111111010001111010101",
			2248 => "0000000010001111010101",
			2249 => "0010000111110100000100",
			2250 => "0000000010001111010101",
			2251 => "0000000001110100000100",
			2252 => "0000001010001111010101",
			2253 => "0000000010001111010101",
			2254 => "0011111100010000001000",
			2255 => "0010100000001000000100",
			2256 => "0000000010001111010101",
			2257 => "0000001010001111010101",
			2258 => "0011001010111000001000",
			2259 => "0011010101110000000100",
			2260 => "1111111010001111010101",
			2261 => "0000000010001111010101",
			2262 => "0001100100110100000100",
			2263 => "1111111010001111010101",
			2264 => "0000000010001111010101",
			2265 => "0011010010011100010000",
			2266 => "0011001000000000001100",
			2267 => "0000000110001000001000",
			2268 => "0000011001011000000100",
			2269 => "0000000010001111010101",
			2270 => "0000000010001111010101",
			2271 => "0000000010001111010101",
			2272 => "1111111010001111010101",
			2273 => "0011011110010000010000",
			2274 => "0001100100110100001000",
			2275 => "0001101101111100000100",
			2276 => "0000001010001111010101",
			2277 => "0000000010001111010101",
			2278 => "0000001010101100000100",
			2279 => "0000001010001111010101",
			2280 => "0000000010001111010101",
			2281 => "0001111000011000000100",
			2282 => "0000000010001111010101",
			2283 => "0011011100010100000100",
			2284 => "0000000010001111010101",
			2285 => "0000000010001111010101",
			2286 => "0010110101110100000100",
			2287 => "1111110010001111010101",
			2288 => "0001101001100100000100",
			2289 => "0000000010001111010101",
			2290 => "0001110111010000000100",
			2291 => "0000000010001111010101",
			2292 => "1111111010001111010101",
			2293 => "0000001010101110000000",
			2294 => "0000010000111101000000",
			2295 => "0001111000011000100100",
			2296 => "0001110001101000011000",
			2297 => "0000111100000000010000",
			2298 => "0011000100011000001000",
			2299 => "0001110110100100000100",
			2300 => "1111111010010011011011",
			2301 => "0000000010010011011011",
			2302 => "0010011111000000000100",
			2303 => "0000000010010011011011",
			2304 => "0000001010010011011011",
			2305 => "0001011100100100000100",
			2306 => "0000000010010011011011",
			2307 => "1111111010010011011011",
			2308 => "0000000101000100001000",
			2309 => "0000111100000000000100",
			2310 => "0000000010010011011011",
			2311 => "0000000010010011011011",
			2312 => "0000001010010011011011",
			2313 => "0000110110111100001100",
			2314 => "0001111000011000001000",
			2315 => "0000100110010000000100",
			2316 => "0000000010010011011011",
			2317 => "0000000010010011011011",
			2318 => "0000010010010011011011",
			2319 => "0000000001010100000100",
			2320 => "1111111010010011011011",
			2321 => "0001111000011000000100",
			2322 => "1111111010010011011011",
			2323 => "0000100110111100000100",
			2324 => "0000001010010011011011",
			2325 => "1111111010010011011011",
			2326 => "0001110001101000100000",
			2327 => "0011001001001000011100",
			2328 => "0000001111001000001100",
			2329 => "0000011101111100001000",
			2330 => "0001010110100000000100",
			2331 => "0000000010010011011011",
			2332 => "0000001010010011011011",
			2333 => "1111111010010011011011",
			2334 => "0001101111000000001000",
			2335 => "0011001011000000000100",
			2336 => "1111111010010011011011",
			2337 => "0000000010010011011011",
			2338 => "0001011100100100000100",
			2339 => "1111111010010011011011",
			2340 => "0000001010010011011011",
			2341 => "1111111010010011011011",
			2342 => "0011010110010000011000",
			2343 => "0010010100111100001000",
			2344 => "0000100111011000000100",
			2345 => "0000000010010011011011",
			2346 => "0000000010010011011011",
			2347 => "0010111011011100001000",
			2348 => "0000001111001000000100",
			2349 => "0000001010010011011011",
			2350 => "0000000010010011011011",
			2351 => "0000001010101100000100",
			2352 => "0000001010010011011011",
			2353 => "0000010010010011011011",
			2354 => "0001110101110100000100",
			2355 => "1111111010010011011011",
			2356 => "0000000010010011011011",
			2357 => "1111111010010011011011",
			2358 => "0000000010010011011101",
			2359 => "0000000010010011100001",
			2360 => "0000000010010011100101",
			2361 => "0011001011000000000100",
			2362 => "0000000010010011111001",
			2363 => "0011000110100100000100",
			2364 => "0000000010010011111001",
			2365 => "0000000010010011111001",
			2366 => "0011001010111000000100",
			2367 => "0000000010010100001101",
			2368 => "0000000001110100000100",
			2369 => "0000000010010100001101",
			2370 => "0000000010010100001101",
			2371 => "0000001100000100001000",
			2372 => "0000000011101000000100",
			2373 => "0000000010010100100001",
			2374 => "0000000010010100100001",
			2375 => "0000000010010100100001",
			2376 => "0001011100100100001000",
			2377 => "0001010110110100000100",
			2378 => "0000000010010100111101",
			2379 => "0000000010010100111101",
			2380 => "0001011111010000000100",
			2381 => "0000000010010100111101",
			2382 => "0000000010010100111101",
			2383 => "0001001101101100001000",
			2384 => "0000101101000100000100",
			2385 => "0000000010010101011001",
			2386 => "0000000010010101011001",
			2387 => "0000101000101000000100",
			2388 => "0000000010010101011001",
			2389 => "0000000010010101011001",
			2390 => "0011100111010100001100",
			2391 => "0001110001101000001000",
			2392 => "0010011001111100000100",
			2393 => "0000000010010101111101",
			2394 => "0000000010010101111101",
			2395 => "0000000010010101111101",
			2396 => "0000101101101100000100",
			2397 => "0000000010010101111101",
			2398 => "0000000010010101111101",
			2399 => "0011001001110100001100",
			2400 => "0011000100011000000100",
			2401 => "0000000010010110100001",
			2402 => "0011001011000000000100",
			2403 => "0000000010010110100001",
			2404 => "0000000010010110100001",
			2405 => "0011000110100100000100",
			2406 => "0000000010010110100001",
			2407 => "0000000010010110100001",
			2408 => "0000001001101000001100",
			2409 => "0000100010000100000100",
			2410 => "0000000010010111001101",
			2411 => "0011000100011000000100",
			2412 => "0000000010010111001101",
			2413 => "0000000010010111001101",
			2414 => "0011001001110100001000",
			2415 => "0000100010010100000100",
			2416 => "0000000010010111001101",
			2417 => "0000000010010111001101",
			2418 => "0000000010010111001101",
			2419 => "0001001100010000000100",
			2420 => "0000000010010111110001",
			2421 => "0010111011110100001100",
			2422 => "0011101100111000001000",
			2423 => "0000110001011100000100",
			2424 => "0000000010010111110001",
			2425 => "0000000010010111110001",
			2426 => "0000000010010111110001",
			2427 => "0000000010010111110001",
			2428 => "0001001101101100010000",
			2429 => "0001010110100000000100",
			2430 => "0000000010011000010101",
			2431 => "0001010101001000001000",
			2432 => "0001000010000000000100",
			2433 => "0000000010011000010101",
			2434 => "0000000010011000010101",
			2435 => "0000000010011000010101",
			2436 => "0000000010011000010101",
			2437 => "0011001001110100010000",
			2438 => "0001101101111100000100",
			2439 => "0000000010011001000001",
			2440 => "0001101001100100001000",
			2441 => "0010110000011100000100",
			2442 => "0000000010011001000001",
			2443 => "0000000010011001000001",
			2444 => "0000000010011001000001",
			2445 => "0011000110100100000100",
			2446 => "0000000010011001000001",
			2447 => "0000000010011001000001",
			2448 => "0001101101111100001000",
			2449 => "0011000100011000000100",
			2450 => "0000000010011001101101",
			2451 => "0000000010011001101101",
			2452 => "0011001001110100001100",
			2453 => "0001001010000100000100",
			2454 => "0000000010011001101101",
			2455 => "0001101011001100000100",
			2456 => "0000000010011001101101",
			2457 => "0000000010011001101101",
			2458 => "0000000010011001101101",
			2459 => "0000101100010000001100",
			2460 => "0000001100000100001000",
			2461 => "0000101101000100000100",
			2462 => "0000000010011010100001",
			2463 => "0000000010011010100001",
			2464 => "0000000010011010100001",
			2465 => "0000101010000100000100",
			2466 => "0000000010011010100001",
			2467 => "0000000111000100001000",
			2468 => "0000001001101000000100",
			2469 => "0000000010011010100001",
			2470 => "0000000010011010100001",
			2471 => "0000000010011010100001",
			2472 => "0001000001011100010100",
			2473 => "0010100000001000000100",
			2474 => "0000000010011011010101",
			2475 => "0000010111101000001100",
			2476 => "0010011111000000000100",
			2477 => "0000000010011011010101",
			2478 => "0011100010000000000100",
			2479 => "0000000010011011010101",
			2480 => "0000000010011011010101",
			2481 => "0000000010011011010101",
			2482 => "0010011010100100000100",
			2483 => "0000000010011011010101",
			2484 => "0000000010011011010101",
			2485 => "0000000111000100010100",
			2486 => "0011001010111000000100",
			2487 => "0000000010011100000001",
			2488 => "0011011010001000001100",
			2489 => "0011011110000100000100",
			2490 => "0000000010011100000001",
			2491 => "0010100000001000000100",
			2492 => "0000000010011100000001",
			2493 => "0000000010011100000001",
			2494 => "0000000010011100000001",
			2495 => "0000000010011100000001",
			2496 => "0001011111010000010100",
			2497 => "0011000100011000000100",
			2498 => "0000000010011100101101",
			2499 => "0000000010101000001100",
			2500 => "0011001001001000001000",
			2501 => "0011011001011100000100",
			2502 => "0000000010011100101101",
			2503 => "0000000010011100101101",
			2504 => "0000000010011100101101",
			2505 => "0000000010011100101101",
			2506 => "0000000010011100101101",
			2507 => "0000010000111100001100",
			2508 => "0000101100010000000100",
			2509 => "0000000010011101101001",
			2510 => "0011010111111100000100",
			2511 => "0000000010011101101001",
			2512 => "0000000010011101101001",
			2513 => "0011000100011000000100",
			2514 => "0000000010011101101001",
			2515 => "0000100110111000001100",
			2516 => "0000011010011000001000",
			2517 => "0011010010011100000100",
			2518 => "0000000010011101101001",
			2519 => "0000000010011101101001",
			2520 => "0000000010011101101001",
			2521 => "0000000010011101101001",
			2522 => "0001010110100000001000",
			2523 => "0011100111010100000100",
			2524 => "0000000010011110101101",
			2525 => "0000000010011110101101",
			2526 => "0001011100100100010000",
			2527 => "0000101101101100001100",
			2528 => "0011100010000000000100",
			2529 => "0000000010011110101101",
			2530 => "0000100110010000000100",
			2531 => "0000000010011110101101",
			2532 => "0000000010011110101101",
			2533 => "0000000010011110101101",
			2534 => "0001111000011000000100",
			2535 => "0000000010011110101101",
			2536 => "0001110101100100000100",
			2537 => "0000000010011110101101",
			2538 => "0000000010011110101101",
			2539 => "0000001100000100010000",
			2540 => "0010010101010000001100",
			2541 => "0001000110111100001000",
			2542 => "0010111001110100000100",
			2543 => "0000000010100000000001",
			2544 => "0000000010100000000001",
			2545 => "0000000010100000000001",
			2546 => "0000000010100000000001",
			2547 => "0010010111101100001100",
			2548 => "0010111011110100001000",
			2549 => "0010110000011100000100",
			2550 => "0000000010100000000001",
			2551 => "0000000010100000000001",
			2552 => "0000000010100000000001",
			2553 => "0000000001110100001100",
			2554 => "0010110101100100000100",
			2555 => "0000000010100000000001",
			2556 => "0010111011110100000100",
			2557 => "0000000010100000000001",
			2558 => "0000000010100000000001",
			2559 => "0000000010100000000001",
			2560 => "0001000001011100011000",
			2561 => "0010010100111100000100",
			2562 => "0000000010100000111101",
			2563 => "0000011101111100010000",
			2564 => "0001110110100100000100",
			2565 => "0000000010100000111101",
			2566 => "0010110100000100000100",
			2567 => "0000000010100000111101",
			2568 => "0010100111110100000100",
			2569 => "0000000010100000111101",
			2570 => "0000000010100000111101",
			2571 => "0000000010100000111101",
			2572 => "0010011010100000000100",
			2573 => "0000000010100000111101",
			2574 => "0000000010100000111101",
			2575 => "0011101100000000001000",
			2576 => "0011011001010100000100",
			2577 => "0000000010100001111001",
			2578 => "0000000010100001111001",
			2579 => "0011010011001000010100",
			2580 => "0010010100111100000100",
			2581 => "0000000010100001111001",
			2582 => "0011100010010100001100",
			2583 => "0011011110000100000100",
			2584 => "0000000010100001111001",
			2585 => "0010010010101100000100",
			2586 => "0000000010100001111001",
			2587 => "0000000010100001111001",
			2588 => "0000000010100001111001",
			2589 => "0000000010100001111001",
			2590 => "0000010000111100001000",
			2591 => "0010101001100100000100",
			2592 => "0000000010100010110101",
			2593 => "0000000010100010110101",
			2594 => "0011111011110000010100",
			2595 => "0000011100011000010000",
			2596 => "0010010100111100000100",
			2597 => "0000000010100010110101",
			2598 => "0010101010100000000100",
			2599 => "0000000010100010110101",
			2600 => "0010101001000100000100",
			2601 => "0000000010100010110101",
			2602 => "0000000010100010110101",
			2603 => "0000000010100010110101",
			2604 => "0000000010100010110101",
			2605 => "0001101001100100011100",
			2606 => "0001000110101100010000",
			2607 => "0011001011000000001000",
			2608 => "0011001010111000000100",
			2609 => "0000000010100100010001",
			2610 => "0000000010100100010001",
			2611 => "0011001001110100000100",
			2612 => "0000000010100100010001",
			2613 => "0000000010100100010001",
			2614 => "0010111011110100001000",
			2615 => "0010101010100000000100",
			2616 => "0000000010100100010001",
			2617 => "0000000010100100010001",
			2618 => "0000000010100100010001",
			2619 => "0000000001110100010000",
			2620 => "0001010101110000001100",
			2621 => "0011001010111000000100",
			2622 => "0000000010100100010001",
			2623 => "0011101010000100000100",
			2624 => "0000000010100100010001",
			2625 => "0000000010100100010001",
			2626 => "0000000010100100010001",
			2627 => "0000000010100100010001",
			2628 => "0001000001011100011000",
			2629 => "0000111000100000010100",
			2630 => "0011001010111000000100",
			2631 => "0000000010100101000101",
			2632 => "0011001001001000001100",
			2633 => "0001111000011000001000",
			2634 => "0000001001101000000100",
			2635 => "0000000010100101000101",
			2636 => "0000000010100101000101",
			2637 => "0000000010100101000101",
			2638 => "0000000010100101000101",
			2639 => "0000000010100101000101",
			2640 => "0000000010100101000101",
			2641 => "0000000010101000011100",
			2642 => "0011101100000000001000",
			2643 => "0001001100010000000100",
			2644 => "0000000010100110000001",
			2645 => "0000000010100110000001",
			2646 => "0011011001010000000100",
			2647 => "0000000010100110000001",
			2648 => "0001011001010000001100",
			2649 => "0011001010111000000100",
			2650 => "0000000010100110000001",
			2651 => "0010010100111100000100",
			2652 => "0000000010100110000001",
			2653 => "0000000010100110000001",
			2654 => "0000000010100110000001",
			2655 => "0000000010100110000001",
			2656 => "0011111100000000001100",
			2657 => "0010001000100100001000",
			2658 => "0001110110100100000100",
			2659 => "0000000010100111011101",
			2660 => "0000000010100111011101",
			2661 => "0000000010100111011101",
			2662 => "0011001000000000010000",
			2663 => "0010100010101100001000",
			2664 => "0001101101111100000100",
			2665 => "0000000010100111011101",
			2666 => "0000000010100111011101",
			2667 => "0010101000100100000100",
			2668 => "0000000010100111011101",
			2669 => "0000000010100111011101",
			2670 => "0011000110100100010000",
			2671 => "0011011100010100001100",
			2672 => "0011101110110100000100",
			2673 => "0000000010100111011101",
			2674 => "0010101001000100000100",
			2675 => "0000000010100111011101",
			2676 => "0000000010100111011101",
			2677 => "0000000010100111011101",
			2678 => "0000000010100111011101",
			2679 => "0001001011101100100100",
			2680 => "0011001011000000010000",
			2681 => "0011000100011000000100",
			2682 => "0000000010101001001001",
			2683 => "0010100111101100000100",
			2684 => "0000000010101001001001",
			2685 => "0010110100000100000100",
			2686 => "0000000010101001001001",
			2687 => "0000000010101001001001",
			2688 => "0010110100010000010000",
			2689 => "0000001001101000001100",
			2690 => "0011001001110100001000",
			2691 => "0000100010000000000100",
			2692 => "0000000010101001001001",
			2693 => "0000000010101001001001",
			2694 => "0000000010101001001001",
			2695 => "0000000010101001001001",
			2696 => "0000000010101001001001",
			2697 => "0000101000100000001100",
			2698 => "0000001011010100000100",
			2699 => "0000000010101001001001",
			2700 => "0010110101100100000100",
			2701 => "0000000010101001001001",
			2702 => "0000000010101001001001",
			2703 => "0000101101101100000100",
			2704 => "0000000010101001001001",
			2705 => "0000000010101001001001",
			2706 => "0001000001011100100000",
			2707 => "0010001000100100001000",
			2708 => "0000011001011000000100",
			2709 => "0000000010101010011101",
			2710 => "0000000010101010011101",
			2711 => "0001110110100100000100",
			2712 => "0000000010101010011101",
			2713 => "0001100100110100000100",
			2714 => "0000000010101010011101",
			2715 => "0011000001101000001100",
			2716 => "0001101101011000001000",
			2717 => "0000001001101000000100",
			2718 => "0000000010101010011101",
			2719 => "0000000010101010011101",
			2720 => "0000000010101010011101",
			2721 => "0000000010101010011101",
			2722 => "0001101000010000001000",
			2723 => "0011001000011000000100",
			2724 => "0000000010101010011101",
			2725 => "0000000010101010011101",
			2726 => "0000000010101010011101",
			2727 => "0001000001011100011100",
			2728 => "0010100000001000000100",
			2729 => "0000000010101011101001",
			2730 => "0011000100011000000100",
			2731 => "0000000010101011101001",
			2732 => "0011000001101000010000",
			2733 => "0011100010000000000100",
			2734 => "0000000010101011101001",
			2735 => "0010011111000000000100",
			2736 => "0000000010101011101001",
			2737 => "0011010001000000000100",
			2738 => "0000000010101011101001",
			2739 => "0000000010101011101001",
			2740 => "0000000010101011101001",
			2741 => "0001100100111100001000",
			2742 => "0011000001011000000100",
			2743 => "0000000010101011101001",
			2744 => "0000000010101011101001",
			2745 => "0000000010101011101001",
			2746 => "0011001001110100011100",
			2747 => "0010011010100000011000",
			2748 => "0010110000011100000100",
			2749 => "0000000010101100101101",
			2750 => "0000011001011000000100",
			2751 => "0000000010101100101101",
			2752 => "0011111001100000000100",
			2753 => "0000000010101100101101",
			2754 => "0010001100011100001000",
			2755 => "0001111001001000000100",
			2756 => "0000000010101100101101",
			2757 => "0000000010101100101101",
			2758 => "0000000010101100101101",
			2759 => "0000000010101100101101",
			2760 => "0011000110100100000100",
			2761 => "0000000010101100101101",
			2762 => "0000000010101100101101",
			2763 => "0010011010100000100100",
			2764 => "0010110101100100010100",
			2765 => "0010111001110100000100",
			2766 => "0000000010101110011001",
			2767 => "0000011101111100001100",
			2768 => "0011111011101100001000",
			2769 => "0011101110101100000100",
			2770 => "0000000010101110011001",
			2771 => "0000000010101110011001",
			2772 => "0000000010101110011001",
			2773 => "0000000010101110011001",
			2774 => "0010110110110100001100",
			2775 => "0011111001100000000100",
			2776 => "0000000010101110011001",
			2777 => "0011101000001100000100",
			2778 => "0000000010101110011001",
			2779 => "0000000010101110011001",
			2780 => "0000000010101110011001",
			2781 => "0010111010010100010000",
			2782 => "0001011110101000000100",
			2783 => "0000000010101110011001",
			2784 => "0011111110000000001000",
			2785 => "0000101011110000000100",
			2786 => "0000000010101110011001",
			2787 => "0000000010101110011001",
			2788 => "0000000010101110011001",
			2789 => "0000000010101110011001",
			2790 => "0001011111010000100100",
			2791 => "0001011101000100001100",
			2792 => "0000000001010100000100",
			2793 => "0000000010101111111101",
			2794 => "0001101011001100000100",
			2795 => "0000000010101111111101",
			2796 => "0000000010101111111101",
			2797 => "0011001001001000010100",
			2798 => "0001100100110100000100",
			2799 => "0000000010101111111101",
			2800 => "0000101101101100001100",
			2801 => "0010001000100100000100",
			2802 => "0000000010101111111101",
			2803 => "0010101000100100000100",
			2804 => "0000000010101111111101",
			2805 => "0000000010101111111101",
			2806 => "0000000010101111111101",
			2807 => "0000000010101111111101",
			2808 => "0010111011110100001100",
			2809 => "0011100001011100001000",
			2810 => "0000111000100000000100",
			2811 => "0000000010101111111101",
			2812 => "0000000010101111111101",
			2813 => "0000000010101111111101",
			2814 => "0000000010101111111101",
			2815 => "0011010101110000011100",
			2816 => "0000001111001000010100",
			2817 => "0010011111000000000100",
			2818 => "0000000010110001111001",
			2819 => "0001110110100100000100",
			2820 => "0000000010110001111001",
			2821 => "0010110110110100001000",
			2822 => "0011010001000000000100",
			2823 => "0000000010110001111001",
			2824 => "0000000010110001111001",
			2825 => "0000000010110001111001",
			2826 => "0011010101110000000100",
			2827 => "0000000010110001111001",
			2828 => "0000000010110001111001",
			2829 => "0001101100011000010000",
			2830 => "0010100000001000000100",
			2831 => "0000000010110001111001",
			2832 => "0010110110110100000100",
			2833 => "0000000010110001111001",
			2834 => "0000100110111100000100",
			2835 => "0000000010110001111001",
			2836 => "0000000010110001111001",
			2837 => "0010100011101000001000",
			2838 => "0001111111011100000100",
			2839 => "0000000010110001111001",
			2840 => "0000000010110001111001",
			2841 => "0000000001110100001000",
			2842 => "0000101000101000000100",
			2843 => "0000000010110001111001",
			2844 => "0000000010110001111001",
			2845 => "0000000010110001111001",
			2846 => "0001001100010000000100",
			2847 => "0000000010110010110101",
			2848 => "0010110110110100011000",
			2849 => "0011101100111000010100",
			2850 => "0010110101100100000100",
			2851 => "0000000010110010110101",
			2852 => "0001111001001000000100",
			2853 => "0000000010110010110101",
			2854 => "0001010101001000001000",
			2855 => "0001111000011000000100",
			2856 => "0000000010110010110101",
			2857 => "0000000010110010110101",
			2858 => "0000000010110010110101",
			2859 => "0000000010110010110101",
			2860 => "0000000010110010110101",
			2861 => "0010011111000000000100",
			2862 => "0000000010110011110001",
			2863 => "0000001010101100011000",
			2864 => "0011000100011000000100",
			2865 => "0000000010110011110001",
			2866 => "0001011110010000010000",
			2867 => "0010100000001000000100",
			2868 => "0000000010110011110001",
			2869 => "0000011010011000001000",
			2870 => "0010110100000100000100",
			2871 => "0000000010110011110001",
			2872 => "0000000010110011110001",
			2873 => "0000000010110011110001",
			2874 => "0000000010110011110001",
			2875 => "0000000010110011110001",
			2876 => "0000000010101000011100",
			2877 => "0011001101010100000100",
			2878 => "0000000010110100101101",
			2879 => "0010011111000000000100",
			2880 => "0000000010110100101101",
			2881 => "0001110110100100000100",
			2882 => "0000000010110100101101",
			2883 => "0000101110110100000100",
			2884 => "0000000010110100101101",
			2885 => "0000011010011000001000",
			2886 => "0000110010010100000100",
			2887 => "0000000010110100101101",
			2888 => "0000000010110100101101",
			2889 => "0000000010110100101101",
			2890 => "0000000010110100101101",
			2891 => "0001001100010000000100",
			2892 => "0000000010110101111001",
			2893 => "0001011111010000011100",
			2894 => "0011100111010100010100",
			2895 => "0010110100010000010000",
			2896 => "0010110000011100000100",
			2897 => "0000000010110101111001",
			2898 => "0011001010111000000100",
			2899 => "0000000010110101111001",
			2900 => "0000110000010000000100",
			2901 => "0000000010110101111001",
			2902 => "0000000010110101111001",
			2903 => "0000000010110101111001",
			2904 => "0010101000100100000100",
			2905 => "0000000010110101111001",
			2906 => "0000000010110101111001",
			2907 => "0000111000001100000100",
			2908 => "0000000010110101111001",
			2909 => "0000000010110101111001",
			2910 => "0000001001101000011100",
			2911 => "0000011011111100010000",
			2912 => "0001111011000000000100",
			2913 => "0000000010111000000101",
			2914 => "0011111111010100001000",
			2915 => "0000110111010100000100",
			2916 => "0000000010111000000101",
			2917 => "0000000010111000000101",
			2918 => "0000000010111000000101",
			2919 => "0010100010101100001000",
			2920 => "0001111001001000000100",
			2921 => "0000000010111000000101",
			2922 => "0000000010111000000101",
			2923 => "0000000010111000000101",
			2924 => "0010010111101100010000",
			2925 => "0001110110110100001100",
			2926 => "0001001000100000001000",
			2927 => "0001000110101100000100",
			2928 => "0000000010111000000101",
			2929 => "0000000010111000000101",
			2930 => "0000000010111000000101",
			2931 => "0000000010111000000101",
			2932 => "0011010010011100010000",
			2933 => "0001010110100000000100",
			2934 => "0000000010111000000101",
			2935 => "0011101010000100000100",
			2936 => "0000000010111000000101",
			2937 => "0001011100100100000100",
			2938 => "0000000010111000000101",
			2939 => "0000000010111000000101",
			2940 => "0011011100010100001000",
			2941 => "0011100110111000000100",
			2942 => "0000000010111000000101",
			2943 => "0000000010111000000101",
			2944 => "0000000010111000000101",
			2945 => "0011001011000000101000",
			2946 => "0001001100010000001000",
			2947 => "0000011101101000000100",
			2948 => "0000000010111010000001",
			2949 => "0000000010111010000001",
			2950 => "0010010100101100010000",
			2951 => "0001111000011000001100",
			2952 => "0001101101111100000100",
			2953 => "0000000010111010000001",
			2954 => "0010110101100100000100",
			2955 => "0000000010111010000001",
			2956 => "0000000010111010000001",
			2957 => "0000000010111010000001",
			2958 => "0000011101111100001100",
			2959 => "0001110001101000001000",
			2960 => "0001111000000000000100",
			2961 => "0000000010111010000001",
			2962 => "0000000010111010000001",
			2963 => "0000000010111010000001",
			2964 => "0000000010111010000001",
			2965 => "0000000101000100000100",
			2966 => "0000000010111010000001",
			2967 => "0001101100011000001000",
			2968 => "0011001000000000000100",
			2969 => "0000000010111010000001",
			2970 => "0000000010111010000001",
			2971 => "0000010001000100000100",
			2972 => "0000000010111010000001",
			2973 => "0000011010011000000100",
			2974 => "0000000010111010000001",
			2975 => "0000000010111010000001",
			2976 => "0011100111010100101100",
			2977 => "0000001100000100011100",
			2978 => "0000111010000100010100",
			2979 => "0010011111000000000100",
			2980 => "0000000010111011111101",
			2981 => "0001101100011000001100",
			2982 => "0000011001011000000100",
			2983 => "0000000010111011111101",
			2984 => "0000000101000100000100",
			2985 => "0000000010111011111101",
			2986 => "0000000010111011111101",
			2987 => "0000000010111011111101",
			2988 => "0010001000010100000100",
			2989 => "0000000010111011111101",
			2990 => "0000000010111011111101",
			2991 => "0001010010110100000100",
			2992 => "0000000010111011111101",
			2993 => "0011011110010000001000",
			2994 => "0010110000011100000100",
			2995 => "0000000010111011111101",
			2996 => "0000000010111011111101",
			2997 => "0000000010111011111101",
			2998 => "0000000001110100010000",
			2999 => "0001001110000000001100",
			3000 => "0010000001010000000100",
			3001 => "0000000010111011111101",
			3002 => "0000011100011000000100",
			3003 => "0000000010111011111101",
			3004 => "0000000010111011111101",
			3005 => "0000000010111011111101",
			3006 => "0000000010111011111101",
			3007 => "0011001011000000101100",
			3008 => "0001000110111100010000",
			3009 => "0011001010111000000100",
			3010 => "0000000010111110000001",
			3011 => "0001111000011000001000",
			3012 => "0001111011000000000100",
			3013 => "0000000010111110000001",
			3014 => "0000000010111110000001",
			3015 => "0000000010111110000001",
			3016 => "0010010111101100001100",
			3017 => "0010110000011100000100",
			3018 => "0000000010111110000001",
			3019 => "0011101100010000000100",
			3020 => "0000000010111110000001",
			3021 => "0000000010111110000001",
			3022 => "0000011101111100001100",
			3023 => "0011101111010100000100",
			3024 => "0000000010111110000001",
			3025 => "0010101000100100000100",
			3026 => "0000000010111110000001",
			3027 => "0000000010111110000001",
			3028 => "0000000010111110000001",
			3029 => "0011101100000000000100",
			3030 => "0000000010111110000001",
			3031 => "0000011100011000010000",
			3032 => "0000010000111100000100",
			3033 => "0000000010111110000001",
			3034 => "0000000111000000001000",
			3035 => "0011010010000100000100",
			3036 => "0000000010111110000001",
			3037 => "0000000010111110000001",
			3038 => "0000000010111110000001",
			3039 => "0000000010111110000001",
			3040 => "0001001011101100110100",
			3041 => "0011010101110000011000",
			3042 => "0001110110100100000100",
			3043 => "0000000011000000010101",
			3044 => "0010011111000000000100",
			3045 => "0000000011000000010101",
			3046 => "0010110110110100001100",
			3047 => "0010100000001000000100",
			3048 => "0000000011000000010101",
			3049 => "0011011110000100000100",
			3050 => "0000000011000000010101",
			3051 => "0000000011000000010101",
			3052 => "0000000011000000010101",
			3053 => "0010110110110100001100",
			3054 => "0000110000010000001000",
			3055 => "0011111001100000000100",
			3056 => "0000000011000000010101",
			3057 => "0000000011000000010101",
			3058 => "0000000011000000010101",
			3059 => "0000110111010100001000",
			3060 => "0011111100000000000100",
			3061 => "0000000011000000010101",
			3062 => "0000000011000000010101",
			3063 => "0000101010000100000100",
			3064 => "0000000011000000010101",
			3065 => "0000000011000000010101",
			3066 => "0000111111100100001100",
			3067 => "0011101000001100001000",
			3068 => "0000001011010100000100",
			3069 => "0000000011000000010101",
			3070 => "0000000011000000010101",
			3071 => "0000000011000000010101",
			3072 => "0000000111000100001000",
			3073 => "0000001011010100000100",
			3074 => "0000000011000000010101",
			3075 => "0000000011000000010101",
			3076 => "0000000011000000010101",
			3077 => "0000001001101000100000",
			3078 => "0011010101001000001100",
			3079 => "0000011011111100001000",
			3080 => "0000011101101000000100",
			3081 => "0000000011000010101001",
			3082 => "0000000011000010101001",
			3083 => "0000000011000010101001",
			3084 => "0001010101001000010000",
			3085 => "0011111110110100000100",
			3086 => "0000000011000010101001",
			3087 => "0010011111000000000100",
			3088 => "0000000011000010101001",
			3089 => "0011100110111100000100",
			3090 => "0000000011000010101001",
			3091 => "0000000011000010101001",
			3092 => "0000000011000010101001",
			3093 => "0000010111101000001100",
			3094 => "0010111010010100001000",
			3095 => "0001000000010000000100",
			3096 => "0000000011000010101001",
			3097 => "0000000011000010101001",
			3098 => "0000000011000010101001",
			3099 => "0001011100100100001100",
			3100 => "0000011101111100000100",
			3101 => "0000000011000010101001",
			3102 => "0001110001101000000100",
			3103 => "0000000011000010101001",
			3104 => "0000000011000010101001",
			3105 => "0011011100010100010000",
			3106 => "0000011010011000001100",
			3107 => "0010111011011100000100",
			3108 => "0000000011000010101001",
			3109 => "0000001010101100000100",
			3110 => "0000000011000010101001",
			3111 => "0000000011000010101001",
			3112 => "0000000011000010101001",
			3113 => "0000000011000010101001",
			3114 => "0000000111000100110100",
			3115 => "0010010111101100101000",
			3116 => "0000101010000100011100",
			3117 => "0010001001000100010100",
			3118 => "0000010101011100001100",
			3119 => "0010010100111100001000",
			3120 => "0001110001101000000100",
			3121 => "0000000011000100011101",
			3122 => "0000000011000100011101",
			3123 => "0000000011000100011101",
			3124 => "0001110001101000000100",
			3125 => "0000000011000100011101",
			3126 => "0000000011000100011101",
			3127 => "0011011111010000000100",
			3128 => "0000000011000100011101",
			3129 => "0000000011000100011101",
			3130 => "0010111011110100001000",
			3131 => "0010010100101100000100",
			3132 => "0000000011000100011101",
			3133 => "0000000011000100011101",
			3134 => "0000000011000100011101",
			3135 => "0000101000001100000100",
			3136 => "0000000011000100011101",
			3137 => "0000111000001100000100",
			3138 => "0000000011000100011101",
			3139 => "0000000011000100011101",
			3140 => "0011100001011100000100",
			3141 => "0000000011000100011101",
			3142 => "0000000011000100011101",
			3143 => "0011100111010100110100",
			3144 => "0000001100000100011100",
			3145 => "0000111010000100010100",
			3146 => "0010011111000000000100",
			3147 => "0000000011000110100001",
			3148 => "0001101100011000001100",
			3149 => "0000011001011000000100",
			3150 => "0000000011000110100001",
			3151 => "0000000101000100000100",
			3152 => "0000000011000110100001",
			3153 => "0000000011000110100001",
			3154 => "0000000011000110100001",
			3155 => "0010001000010100000100",
			3156 => "0000000011000110100001",
			3157 => "0000000011000110100001",
			3158 => "0001010010110100000100",
			3159 => "0000000011000110100001",
			3160 => "0001111001001000000100",
			3161 => "0000000011000110100001",
			3162 => "0010110101110100001100",
			3163 => "0010110000011100000100",
			3164 => "0000000011000110100001",
			3165 => "0001111111011100000100",
			3166 => "0000000011000110100001",
			3167 => "0000000011000110100001",
			3168 => "0000000011000110100001",
			3169 => "0000000001110100001100",
			3170 => "0000011110010100000100",
			3171 => "0000000011000110100001",
			3172 => "0000011100011000000100",
			3173 => "0000000011000110100001",
			3174 => "0000000011000110100001",
			3175 => "0000000011000110100001",
			3176 => "0001000110111000110000",
			3177 => "0010011111000000010000",
			3178 => "0001111000011000001100",
			3179 => "0010101001100100001000",
			3180 => "0011000000001100000100",
			3181 => "1111111011001001000101",
			3182 => "0000011011001001000101",
			3183 => "1111111011001001000101",
			3184 => "0000000011001001000101",
			3185 => "0011011110000100001000",
			3186 => "0010000110011000000100",
			3187 => "0000001011001001000101",
			3188 => "1111111011001001000101",
			3189 => "0000111000101000010000",
			3190 => "0000011001011000000100",
			3191 => "0000000011001001000101",
			3192 => "0010101000100100001000",
			3193 => "0010100000001000000100",
			3194 => "0000001011001001000101",
			3195 => "0000001011001001000101",
			3196 => "1111111011001001000101",
			3197 => "0001000010010100000100",
			3198 => "1111111011001001000101",
			3199 => "0000001011001001000101",
			3200 => "0001001000110100011000",
			3201 => "0001110001101000000100",
			3202 => "1111111011001001000101",
			3203 => "0011011100010100010000",
			3204 => "0001010101001000001000",
			3205 => "0011010100101000000100",
			3206 => "1111111011001001000101",
			3207 => "0000001011001001000101",
			3208 => "0011110010010100000100",
			3209 => "0000010011001001000101",
			3210 => "0000011011001001000101",
			3211 => "1111111011001001000101",
			3212 => "0001000101000000001000",
			3213 => "0001000101000000000100",
			3214 => "1111111011001001000101",
			3215 => "0000000011001001000101",
			3216 => "1111111011001001000101",
			3217 => "0000000010101000111000",
			3218 => "0010011001100100001100",
			3219 => "0001100000111100001000",
			3220 => "0000100111010000000100",
			3221 => "1111111011001011001001",
			3222 => "0000001011001011001001",
			3223 => "1111111011001011001001",
			3224 => "0011011100010100100100",
			3225 => "0001010110100000001100",
			3226 => "0000011011111100001000",
			3227 => "0011001010111000000100",
			3228 => "0000000011001011001001",
			3229 => "0000001011001011001001",
			3230 => "1111111011001011001001",
			3231 => "0001100100111100010000",
			3232 => "0000001111001000001000",
			3233 => "0000010000111100000100",
			3234 => "0000000011001011001001",
			3235 => "0000001011001011001001",
			3236 => "0000111111100100000100",
			3237 => "1111111011001011001001",
			3238 => "0000001011001011001001",
			3239 => "0000101000101000000100",
			3240 => "0000001011001011001001",
			3241 => "0000010011001011001001",
			3242 => "0000101100111000000100",
			3243 => "0000000011001011001001",
			3244 => "1111111011001011001001",
			3245 => "0000001010101100001000",
			3246 => "0001101000010000000100",
			3247 => "1111111011001011001001",
			3248 => "0000001011001011001001",
			3249 => "1111111011001011001001",
			3250 => "0000000010101000111100",
			3251 => "0000011001011000010000",
			3252 => "0010110010001000001100",
			3253 => "0001100000111100001000",
			3254 => "0000000011101000000100",
			3255 => "1111111011001101010101",
			3256 => "0000001011001101010101",
			3257 => "1111111011001101010101",
			3258 => "0000000011001101010101",
			3259 => "0011011100010100100100",
			3260 => "0001010110100000001100",
			3261 => "0000011011111100001000",
			3262 => "0011001010111000000100",
			3263 => "0000000011001101010101",
			3264 => "0000001011001101010101",
			3265 => "1111111011001101010101",
			3266 => "0001100100111100010000",
			3267 => "0010100000001000001000",
			3268 => "0000111110110100000100",
			3269 => "0000001011001101010101",
			3270 => "1111111011001101010101",
			3271 => "0000001111001000000100",
			3272 => "0000001011001101010101",
			3273 => "0000000011001101010101",
			3274 => "0001011001010000000100",
			3275 => "0000010011001101010101",
			3276 => "0000001011001101010101",
			3277 => "0000101100111000000100",
			3278 => "0000000011001101010101",
			3279 => "1111111011001101010101",
			3280 => "0000001010101100001000",
			3281 => "0001101000010000000100",
			3282 => "1111111011001101010101",
			3283 => "0000001011001101010101",
			3284 => "1111111011001101010101",
			3285 => "0011111100000000010000",
			3286 => "0010101001100100000100",
			3287 => "0000000011001111111001",
			3288 => "0010010100111100001000",
			3289 => "0000010000111100000100",
			3290 => "0000000011001111111001",
			3291 => "0000000011001111111001",
			3292 => "0000000011001111111001",
			3293 => "0000100000010000100100",
			3294 => "0010100010101100010100",
			3295 => "0010110110110100001000",
			3296 => "0001011100100100000100",
			3297 => "0000000011001111111001",
			3298 => "0000000011001111111001",
			3299 => "0010011111000000000100",
			3300 => "0000000011001111111001",
			3301 => "0000011001011000000100",
			3302 => "0000000011001111111001",
			3303 => "0000000011001111111001",
			3304 => "0000110110111100000100",
			3305 => "0000000011001111111001",
			3306 => "0011011110000100000100",
			3307 => "0000000011001111111001",
			3308 => "0010100111110100000100",
			3309 => "0000000011001111111001",
			3310 => "0000000011001111111001",
			3311 => "0011101000001100000100",
			3312 => "0000000011001111111001",
			3313 => "0011011100010100010100",
			3314 => "0000000001110100001000",
			3315 => "0001101001100100000100",
			3316 => "0000000011001111111001",
			3317 => "0000000011001111111001",
			3318 => "0010011010100100000100",
			3319 => "0000000011001111111001",
			3320 => "0000110001011100000100",
			3321 => "0000000011001111111001",
			3322 => "0000000011001111111001",
			3323 => "0010110001001000000100",
			3324 => "0000000011001111111001",
			3325 => "0000000011001111111001",
			3326 => "0000000001110100111100",
			3327 => "0010011111000000010000",
			3328 => "0001010101001000001100",
			3329 => "0001100000111100001000",
			3330 => "0010010001000100000100",
			3331 => "1111111011010010011101",
			3332 => "0000001011010010011101",
			3333 => "1111111011010010011101",
			3334 => "0000000011010010011101",
			3335 => "0011010001000000001000",
			3336 => "0010011001111100000100",
			3337 => "0000000011010010011101",
			3338 => "1111111011010010011101",
			3339 => "0011011100010100011100",
			3340 => "0010100000001000001100",
			3341 => "0000111100010000000100",
			3342 => "0000001011010010011101",
			3343 => "0001011100100100000100",
			3344 => "0000000011010010011101",
			3345 => "1111111011010010011101",
			3346 => "0011001010111000001000",
			3347 => "0000000110001000000100",
			3348 => "0000001011010010011101",
			3349 => "1111111011010010011101",
			3350 => "0000111100111000000100",
			3351 => "0000001011010010011101",
			3352 => "0000001011010010011101",
			3353 => "0000001111001000000100",
			3354 => "0000000011010010011101",
			3355 => "1111111011010010011101",
			3356 => "0000001010101100010100",
			3357 => "0010000001010100001100",
			3358 => "0000000001110100001000",
			3359 => "0010000101000100000100",
			3360 => "1111111011010010011101",
			3361 => "0000001011010010011101",
			3362 => "1111111011010010011101",
			3363 => "0001101000010000000100",
			3364 => "0000000011010010011101",
			3365 => "0000010011010010011101",
			3366 => "1111111011010010011101",
			3367 => "0001001011110000110100",
			3368 => "0000011001011000001100",
			3369 => "0001100000111100001000",
			3370 => "0011101011000000000100",
			3371 => "1111111011010100111001",
			3372 => "0000001011010100111001",
			3373 => "1111111011010100111001",
			3374 => "0011011110000100001100",
			3375 => "0001001100010000000100",
			3376 => "0000001011010100111001",
			3377 => "0001011101000100000100",
			3378 => "1111111011010100111001",
			3379 => "0000000011010100111001",
			3380 => "0000011100011000011000",
			3381 => "0010100000001000001000",
			3382 => "0000101100010100000100",
			3383 => "0000000011010100111001",
			3384 => "1111111011010100111001",
			3385 => "0000101100000000001000",
			3386 => "0001011111010000000100",
			3387 => "0000001011010100111001",
			3388 => "0000000011010100111001",
			3389 => "0010001000010100000100",
			3390 => "0000000011010100111001",
			3391 => "0000001011010100111001",
			3392 => "1111111011010100111001",
			3393 => "0000010100110100000100",
			3394 => "1111111011010100111001",
			3395 => "0000110110111000010100",
			3396 => "0011010111111100000100",
			3397 => "1111111011010100111001",
			3398 => "0001111000011000001000",
			3399 => "0001000101000000000100",
			3400 => "0000010011010100111001",
			3401 => "0000000011010100111001",
			3402 => "0001100101010000000100",
			3403 => "1111111011010100111001",
			3404 => "0000000011010100111001",
			3405 => "1111111011010100111001",
			3406 => "0000001001101000101000",
			3407 => "0011010101001000001100",
			3408 => "0000011011111100001000",
			3409 => "0000011101101000000100",
			3410 => "0000000011010111111101",
			3411 => "0000000011010111111101",
			3412 => "0000000011010111111101",
			3413 => "0001101100011000010100",
			3414 => "0011101100010000001100",
			3415 => "0011010111111100001000",
			3416 => "0011010010011100000100",
			3417 => "0000000011010111111101",
			3418 => "0000000011010111111101",
			3419 => "0000000011010111111101",
			3420 => "0011011001011100000100",
			3421 => "0000000011010111111101",
			3422 => "0000000011010111111101",
			3423 => "0000010101011100000100",
			3424 => "0000000011010111111101",
			3425 => "0000000011010111111101",
			3426 => "0001101011001100001100",
			3427 => "0011001001110100001000",
			3428 => "0001000000010000000100",
			3429 => "0000000011010111111101",
			3430 => "0000000011010111111101",
			3431 => "0000000011010111111101",
			3432 => "0001110001101000010000",
			3433 => "0010110000011100000100",
			3434 => "0000000011010111111101",
			3435 => "0010101000010100001000",
			3436 => "0000111010000100000100",
			3437 => "0000000011010111111101",
			3438 => "0000000011010111111101",
			3439 => "0000000011010111111101",
			3440 => "0000110001011100010000",
			3441 => "0010100011101000000100",
			3442 => "0000000011010111111101",
			3443 => "0011100001011100001000",
			3444 => "0001101001100100000100",
			3445 => "0000000011010111111101",
			3446 => "0000000011010111111101",
			3447 => "0000000011010111111101",
			3448 => "0001000101000000001100",
			3449 => "0011011100010100001000",
			3450 => "0001011110000100000100",
			3451 => "0000000011010111111101",
			3452 => "0000000011010111111101",
			3453 => "0000000011010111111101",
			3454 => "0000000011010111111101",
			3455 => "0011000100011000011100",
			3456 => "0011100111010100001000",
			3457 => "0000001001101000000100",
			3458 => "0000000011011010011001",
			3459 => "1111111011011010011001",
			3460 => "0001110001101000010000",
			3461 => "0011110011000000001100",
			3462 => "0001111001001000000100",
			3463 => "0000000011011010011001",
			3464 => "0000000010101000000100",
			3465 => "0000000011011010011001",
			3466 => "0000000011011010011001",
			3467 => "0000000011011010011001",
			3468 => "0000000011011010011001",
			3469 => "0000000010101000110000",
			3470 => "0011101100000000011000",
			3471 => "0011010111111100010000",
			3472 => "0001110110100100000100",
			3473 => "0000000011011010011001",
			3474 => "0010110000011100000100",
			3475 => "0000000011011010011001",
			3476 => "0001111000011000000100",
			3477 => "0000000011011010011001",
			3478 => "0000000011011010011001",
			3479 => "0000101100000000000100",
			3480 => "0000000011011010011001",
			3481 => "0000000011011010011001",
			3482 => "0000010000111100000100",
			3483 => "0000000011011010011001",
			3484 => "0011010010011100001000",
			3485 => "0000011101111100000100",
			3486 => "0000000011011010011001",
			3487 => "0000000011011010011001",
			3488 => "0001011110010000001000",
			3489 => "0000011100011000000100",
			3490 => "0000001011011010011001",
			3491 => "0000000011011010011001",
			3492 => "0000000011011010011001",
			3493 => "0000000011011010011001",
			3494 => "0000000010101001000000",
			3495 => "0000111100111000101100",
			3496 => "0000001111001000100100",
			3497 => "0001101011001100011100",
			3498 => "0011111111010100010000",
			3499 => "0000000001010100001000",
			3500 => "0001010111100000000100",
			3501 => "0000000011011100100101",
			3502 => "0000000011011100100101",
			3503 => "0011011111010000000100",
			3504 => "0000000011011100100101",
			3505 => "0000000011011100100101",
			3506 => "0010111011110100001000",
			3507 => "0000010001000100000100",
			3508 => "1111111011011100100101",
			3509 => "0000000011011100100101",
			3510 => "0000000011011100100101",
			3511 => "0000111010000100000100",
			3512 => "0000000011011100100101",
			3513 => "0000001011011100100101",
			3514 => "0000111000100000000100",
			3515 => "1111111011011100100101",
			3516 => "0000000011011100100101",
			3517 => "0000101101101100000100",
			3518 => "0000001011011100100101",
			3519 => "0010000101000100001000",
			3520 => "0001001110000000000100",
			3521 => "0000000011011100100101",
			3522 => "0000000011011100100101",
			3523 => "0000011010011000000100",
			3524 => "0000000011011100100101",
			3525 => "0000000011011100100101",
			3526 => "0000011100011000000100",
			3527 => "1111111011011100100101",
			3528 => "0000000011011100100101",
			3529 => "0000001001101000101100",
			3530 => "0011010101001000001100",
			3531 => "0000011011111100001000",
			3532 => "0000011101101000000100",
			3533 => "0000000011011111110001",
			3534 => "0000000011011111110001",
			3535 => "0000000011011111110001",
			3536 => "0001101100011000011000",
			3537 => "0011010111111100001100",
			3538 => "0000100110010000000100",
			3539 => "0000000011011111110001",
			3540 => "0011010010011100000100",
			3541 => "0000000011011111110001",
			3542 => "0000000011011111110001",
			3543 => "0010101010100000001000",
			3544 => "0000010000111100000100",
			3545 => "0000000011011111110001",
			3546 => "0000000011011111110001",
			3547 => "0000000011011111110001",
			3548 => "0000101000001100000100",
			3549 => "0000000011011111110001",
			3550 => "0000000011011111110001",
			3551 => "0001101011001100001100",
			3552 => "0011001001110100001000",
			3553 => "0001010010110100000100",
			3554 => "0000000011011111110001",
			3555 => "0000000011011111110001",
			3556 => "0000000011011111110001",
			3557 => "0001110001101000010000",
			3558 => "0010110000011100000100",
			3559 => "0000000011011111110001",
			3560 => "0010101000010100001000",
			3561 => "0000111010000100000100",
			3562 => "0000000011011111110001",
			3563 => "0000000011011111110001",
			3564 => "0000000011011111110001",
			3565 => "0001111000011000010000",
			3566 => "0010010000001000000100",
			3567 => "0000000011011111110001",
			3568 => "0011001001110100001000",
			3569 => "0000110010010100000100",
			3570 => "0000000011011111110001",
			3571 => "0000000011011111110001",
			3572 => "0000000011011111110001",
			3573 => "0011011100010100001100",
			3574 => "0010010111101100000100",
			3575 => "0000000011011111110001",
			3576 => "0011000100011000000100",
			3577 => "0000000011011111110001",
			3578 => "0000000011011111110001",
			3579 => "0000000011011111110001",
			3580 => "0001010001000000111000",
			3581 => "0000101000001100100100",
			3582 => "0000001001101000011000",
			3583 => "0010101010100100010000",
			3584 => "0010110101100100000100",
			3585 => "0000000011100010110101",
			3586 => "0001010111100000001000",
			3587 => "0010110010001000000100",
			3588 => "0000000011100010110101",
			3589 => "0000000011100010110101",
			3590 => "0000000011100010110101",
			3591 => "0011010101001000000100",
			3592 => "0000000011100010110101",
			3593 => "0000000011100010110101",
			3594 => "0011000100011000001000",
			3595 => "0001110001101000000100",
			3596 => "1111111011100010110101",
			3597 => "0000000011100010110101",
			3598 => "0000000011100010110101",
			3599 => "0001000001011100000100",
			3600 => "0000000011100010110101",
			3601 => "0001001011110000001100",
			3602 => "0001111000011000001000",
			3603 => "0011001010111000000100",
			3604 => "0000000011100010110101",
			3605 => "0000000011100010110101",
			3606 => "0000000011100010110101",
			3607 => "0000000011100010110101",
			3608 => "0000000010101000100100",
			3609 => "0010100000001000000100",
			3610 => "0000000011100010110101",
			3611 => "0011011010001000001100",
			3612 => "0010011111000000000100",
			3613 => "0000000011100010110101",
			3614 => "0011000100011000000100",
			3615 => "0000000011100010110101",
			3616 => "0000000011100010110101",
			3617 => "0011001001110100001000",
			3618 => "0010010100111100000100",
			3619 => "0000000011100010110101",
			3620 => "0000000011100010110101",
			3621 => "0000100001011100001000",
			3622 => "0010011010100100000100",
			3623 => "0000000011100010110101",
			3624 => "0000000011100010110101",
			3625 => "0000000011100010110101",
			3626 => "0011001000000000000100",
			3627 => "0000000011100010110101",
			3628 => "0000000011100010110101",
			3629 => "0010011001100100001100",
			3630 => "0010101001100100001000",
			3631 => "0001000111010000000100",
			3632 => "0000000011100101100001",
			3633 => "0000000011100101100001",
			3634 => "1111111011100101100001",
			3635 => "0001001100010000010000",
			3636 => "0000111100000000001100",
			3637 => "0000011001011000000100",
			3638 => "0000000011100101100001",
			3639 => "0010011111000000000100",
			3640 => "0000000011100101100001",
			3641 => "0000001011100101100001",
			3642 => "0000000011100101100001",
			3643 => "0011101100111000100100",
			3644 => "0011001001110100011000",
			3645 => "0011011010001000001100",
			3646 => "0000111100111000001000",
			3647 => "0010011010100000000100",
			3648 => "0000000011100101100001",
			3649 => "1111111011100101100001",
			3650 => "0000001011100101100001",
			3651 => "0000111000100000001000",
			3652 => "0000101111010100000100",
			3653 => "0000000011100101100001",
			3654 => "0000000011100101100001",
			3655 => "1111111011100101100001",
			3656 => "0001001011110000001000",
			3657 => "0000010000111100000100",
			3658 => "0000000011100101100001",
			3659 => "0000001011100101100001",
			3660 => "0000000011100101100001",
			3661 => "0011011100010100010000",
			3662 => "0010101001000100001000",
			3663 => "0010111011011100000100",
			3664 => "0000000011100101100001",
			3665 => "0000001011100101100001",
			3666 => "0011010011001000000100",
			3667 => "0000000011100101100001",
			3668 => "0000000011100101100001",
			3669 => "0010111010010100000100",
			3670 => "0000000011100101100001",
			3671 => "1111111011100101100001",
			3672 => "0000000111000101001000",
			3673 => "0001101101011000110000",
			3674 => "0000011011111100100100",
			3675 => "0011111111010100010100",
			3676 => "0010010100111100010000",
			3677 => "0010110010001000001000",
			3678 => "0000111100000000000100",
			3679 => "0000000011100111111101",
			3680 => "0000000011100111111101",
			3681 => "0000101110110100000100",
			3682 => "0000000011100111111101",
			3683 => "0000000011100111111101",
			3684 => "0000000011100111111101",
			3685 => "0010111011110100001100",
			3686 => "0000010001000100001000",
			3687 => "0011000100011000000100",
			3688 => "0000000011100111111101",
			3689 => "0000000011100111111101",
			3690 => "0000000011100111111101",
			3691 => "0000000011100111111101",
			3692 => "0010100010101100001000",
			3693 => "0001111001001000000100",
			3694 => "0000000011100111111101",
			3695 => "0000000011100111111101",
			3696 => "0000000011100111111101",
			3697 => "0010011001111100000100",
			3698 => "0000000011100111111101",
			3699 => "0011000100011000001100",
			3700 => "0001110110100100001000",
			3701 => "0001111001001000000100",
			3702 => "0000000011100111111101",
			3703 => "0000000011100111111101",
			3704 => "0000000011100111111101",
			3705 => "0000110110111100000100",
			3706 => "0000000011100111111101",
			3707 => "0000001011100111111101",
			3708 => "0011100001011100000100",
			3709 => "0000000011100111111101",
			3710 => "0000000011100111111101",
			3711 => "0000000001110101001000",
			3712 => "0000011001011000100000",
			3713 => "0000011001011000010000",
			3714 => "0010101001100100001000",
			3715 => "0001110001111100000100",
			3716 => "1111111011101011011001",
			3717 => "0000111011101011011001",
			3718 => "0001111000011000000100",
			3719 => "1111111011101011011001",
			3720 => "0000000011101011011001",
			3721 => "0011010010011100001000",
			3722 => "0010110101100100000100",
			3723 => "0000000011101011011001",
			3724 => "0000100011101011011001",
			3725 => "0010110110110100000100",
			3726 => "1111111011101011011001",
			3727 => "0000000011101011011001",
			3728 => "0011011110000100001000",
			3729 => "0000100110010000000100",
			3730 => "0000001011101011011001",
			3731 => "1111111011101011011001",
			3732 => "0011010110010000011000",
			3733 => "0010100000001000001100",
			3734 => "0000111100010000000100",
			3735 => "0000001011101011011001",
			3736 => "0011001000000000000100",
			3737 => "1111111011101011011001",
			3738 => "0000000011101011011001",
			3739 => "0011000111001000000100",
			3740 => "0000000011101011011001",
			3741 => "0001010110100000000100",
			3742 => "0000001011101011011001",
			3743 => "0000010011101011011001",
			3744 => "0000000111000100000100",
			3745 => "0000000011101011011001",
			3746 => "1111111011101011011001",
			3747 => "0000001010101100100100",
			3748 => "0010000001010100011000",
			3749 => "0010000001010100010000",
			3750 => "0000000001110100001100",
			3751 => "0001010101110000001000",
			3752 => "0011001010111000000100",
			3753 => "1111111011101011011001",
			3754 => "0000001011101011011001",
			3755 => "1111111011101011011001",
			3756 => "1111111011101011011001",
			3757 => "0011001001110100000100",
			3758 => "0000011011101011011001",
			3759 => "1111111011101011011001",
			3760 => "0001110111010000001000",
			3761 => "0010110100010000000100",
			3762 => "0000001011101011011001",
			3763 => "0000011011101011011001",
			3764 => "1111111011101011011001",
			3765 => "1111111011101011011001",
			3766 => "0000001001101000111000",
			3767 => "0011010101110000010100",
			3768 => "0011001010111000000100",
			3769 => "0000000011101110011101",
			3770 => "0000010111101000001100",
			3771 => "0010110110110100001000",
			3772 => "0001110011100000000100",
			3773 => "0000000011101110011101",
			3774 => "0000000011101110011101",
			3775 => "0000000011101110011101",
			3776 => "0000000011101110011101",
			3777 => "0011001000000000011000",
			3778 => "0010110110110100001100",
			3779 => "0001011100100100000100",
			3780 => "0000000011101110011101",
			3781 => "0011110010000100000100",
			3782 => "0000000011101110011101",
			3783 => "0000000011101110011101",
			3784 => "0000000001110000001000",
			3785 => "0000101110110100000100",
			3786 => "0000000011101110011101",
			3787 => "0000000011101110011101",
			3788 => "0000000011101110011101",
			3789 => "0000101010000100001000",
			3790 => "0000101110110100000100",
			3791 => "0000000011101110011101",
			3792 => "0000000011101110011101",
			3793 => "0000000011101110011101",
			3794 => "0011100111011000000100",
			3795 => "1111111011101110011101",
			3796 => "0011110000010000000100",
			3797 => "0000000011101110011101",
			3798 => "0001110110100100001100",
			3799 => "0000101101101100001000",
			3800 => "0011011110000100000100",
			3801 => "0000000011101110011101",
			3802 => "0000000011101110011101",
			3803 => "0000000011101110011101",
			3804 => "0000101000100000001000",
			3805 => "0011000100011000000100",
			3806 => "0000000011101110011101",
			3807 => "0000000011101110011101",
			3808 => "0000101101101100001000",
			3809 => "0010000101000100000100",
			3810 => "0000000011101110011101",
			3811 => "0000000011101110011101",
			3812 => "0001111000011000000100",
			3813 => "0000000011101110011101",
			3814 => "0000000011101110011101",
			3815 => "0001110110100100010000",
			3816 => "0001001100000000000100",
			3817 => "0000000011110001110001",
			3818 => "0000110111010100001000",
			3819 => "0010110101100100000100",
			3820 => "1111111011110001110001",
			3821 => "0000000011110001110001",
			3822 => "0000000011110001110001",
			3823 => "0010111011011100100100",
			3824 => "0010110101100100010000",
			3825 => "0000011101111100001100",
			3826 => "0000110110111100000100",
			3827 => "0000000011110001110001",
			3828 => "0001000011000000000100",
			3829 => "0000000011110001110001",
			3830 => "0000000011110001110001",
			3831 => "0000000011110001110001",
			3832 => "0001110110100100000100",
			3833 => "0000000011110001110001",
			3834 => "0011111001100000000100",
			3835 => "0000000011110001110001",
			3836 => "0011001010111000000100",
			3837 => "0000000011110001110001",
			3838 => "0001111000011000000100",
			3839 => "0000000011110001110001",
			3840 => "0000000011110001110001",
			3841 => "0001000001011100100000",
			3842 => "0001110110100100001100",
			3843 => "0010011001111100001000",
			3844 => "0000111100000000000100",
			3845 => "0000000011110001110001",
			3846 => "0000000011110001110001",
			3847 => "0000000011110001110001",
			3848 => "0000010000111100010000",
			3849 => "0010101010100000001000",
			3850 => "0000110111010100000100",
			3851 => "0000000011110001110001",
			3852 => "0000000011110001110001",
			3853 => "0001111111011100000100",
			3854 => "0000000011110001110001",
			3855 => "0000000011110001110001",
			3856 => "0000001011110001110001",
			3857 => "0011101100111000001100",
			3858 => "0001010011001000001000",
			3859 => "0000110011000000000100",
			3860 => "0000000011110001110001",
			3861 => "0000000011110001110001",
			3862 => "0000000011110001110001",
			3863 => "0001001000110100001000",
			3864 => "0011011100010100000100",
			3865 => "0000000011110001110001",
			3866 => "0000000011110001110001",
			3867 => "0000000011110001110001",
			3868 => "0000011110010101000000",
			3869 => "0001001000100000111000",
			3870 => "0011010010011100010000",
			3871 => "0000011001011000000100",
			3872 => "0000000011110101001101",
			3873 => "0011010101001000000100",
			3874 => "0000000011110101001101",
			3875 => "0010100111101100000100",
			3876 => "0000000011110101001101",
			3877 => "0000000011110101001101",
			3878 => "0000100010000100010000",
			3879 => "0011010101110000000100",
			3880 => "0000000011110101001101",
			3881 => "0010101010100000001000",
			3882 => "0000100110010000000100",
			3883 => "0000000011110101001101",
			3884 => "0000000011110101001101",
			3885 => "0000000011110101001101",
			3886 => "0001110001101000001100",
			3887 => "0011101100000000001000",
			3888 => "0010110110110100000100",
			3889 => "0000000011110101001101",
			3890 => "0000000011110101001101",
			3891 => "0000000011110101001101",
			3892 => "0000011001011000000100",
			3893 => "0000000011110101001101",
			3894 => "0000101010000100000100",
			3895 => "0000000011110101001101",
			3896 => "0000000011110101001101",
			3897 => "0011000001101000000100",
			3898 => "0000000011110101001101",
			3899 => "0000000011110101001101",
			3900 => "0010101000100100010100",
			3901 => "0001011101000100000100",
			3902 => "0000000011110101001101",
			3903 => "0011001010111000000100",
			3904 => "0000000011110101001101",
			3905 => "0001001011110000001000",
			3906 => "0000011100011000000100",
			3907 => "0000001011110101001101",
			3908 => "0000000011110101001101",
			3909 => "0000000011110101001101",
			3910 => "0011101100111000001000",
			3911 => "0001110110100100000100",
			3912 => "0000000011110101001101",
			3913 => "0000000011110101001101",
			3914 => "0001001000110100010000",
			3915 => "0011000100011000000100",
			3916 => "0000000011110101001101",
			3917 => "0000111101101100000100",
			3918 => "0000000011110101001101",
			3919 => "0001110111010000000100",
			3920 => "0000000011110101001101",
			3921 => "0000000011110101001101",
			3922 => "0000000011110101001101",
			3923 => "0011001010111000010100",
			3924 => "0000000110001000010000",
			3925 => "0000100111011000001000",
			3926 => "0011001010111000000100",
			3927 => "0000000011111000110001",
			3928 => "0000000011111000110001",
			3929 => "0010110000011100000100",
			3930 => "0000000011111000110001",
			3931 => "0000000011111000110001",
			3932 => "1111111011111000110001",
			3933 => "0011001011000001000000",
			3934 => "0011010100101000100100",
			3935 => "0000011101111100011100",
			3936 => "0011011111010000010000",
			3937 => "0001010010110100001000",
			3938 => "0000001011010100000100",
			3939 => "0000000011111000110001",
			3940 => "0000000011111000110001",
			3941 => "0001010110100000000100",
			3942 => "1111111011111000110001",
			3943 => "0000000011111000110001",
			3944 => "0001101101111100000100",
			3945 => "0000000011111000110001",
			3946 => "0010110110110100000100",
			3947 => "0000001011111000110001",
			3948 => "0000000011111000110001",
			3949 => "0010111011011100000100",
			3950 => "0000000011111000110001",
			3951 => "0000000011111000110001",
			3952 => "0011001011000000001100",
			3953 => "0000011110010100001000",
			3954 => "0011100010000100000100",
			3955 => "0000000011111000110001",
			3956 => "1111111011111000110001",
			3957 => "0000000011111000110001",
			3958 => "0011001011000000001100",
			3959 => "0001011111010000001000",
			3960 => "0001010001000000000100",
			3961 => "0000000011111000110001",
			3962 => "0000000011111000110001",
			3963 => "0000000011111000110001",
			3964 => "0000000011111000110001",
			3965 => "0000101110110100001100",
			3966 => "0000010000111100001000",
			3967 => "0001000010000100000100",
			3968 => "0000000011111000110001",
			3969 => "0000000011111000110001",
			3970 => "0000000011111000110001",
			3971 => "0000011100011000010000",
			3972 => "0000011001011000000100",
			3973 => "0000000011111000110001",
			3974 => "0001001000110100001000",
			3975 => "0001011101000100000100",
			3976 => "0000000011111000110001",
			3977 => "0000001011111000110001",
			3978 => "0000000011111000110001",
			3979 => "0000000011111000110001",
			3980 => "0001011101000100011100",
			3981 => "0000000001010100001100",
			3982 => "0011000100011000000100",
			3983 => "0000000011111100110101",
			3984 => "0010110000011100000100",
			3985 => "0000000011111100110101",
			3986 => "0000000011111100110101",
			3987 => "0011100111010100001000",
			3988 => "0001000010000100000100",
			3989 => "0000000011111100110101",
			3990 => "1111111011111100110101",
			3991 => "0001100100111100000100",
			3992 => "0000000011111100110101",
			3993 => "0000000011111100110101",
			3994 => "0000100111011000110000",
			3995 => "0000000001010100100100",
			3996 => "0000011001011000010000",
			3997 => "0001110001101000000100",
			3998 => "0000000011111100110101",
			3999 => "0000110110111100001000",
			4000 => "0011100110010000000100",
			4001 => "0000000011111100110101",
			4002 => "0000001011111100110101",
			4003 => "0000000011111100110101",
			4004 => "0000100010000100010000",
			4005 => "0000100110010000001000",
			4006 => "0010011111000000000100",
			4007 => "0000000011111100110101",
			4008 => "0000000011111100110101",
			4009 => "0001110001101000000100",
			4010 => "0000000011111100110101",
			4011 => "1111111011111100110101",
			4012 => "0000000011111100110101",
			4013 => "0000011001011000000100",
			4014 => "0000000011111100110101",
			4015 => "0000110111010100000100",
			4016 => "0000001011111100110101",
			4017 => "0000000011111100110101",
			4018 => "0010010100101100011100",
			4019 => "0010110100010000001100",
			4020 => "0001011100100100000100",
			4021 => "0000000011111100110101",
			4022 => "0011001001110100000100",
			4023 => "1111111011111100110101",
			4024 => "0000000011111100110101",
			4025 => "0010101010100100000100",
			4026 => "0000000011111100110101",
			4027 => "0010101010100100000100",
			4028 => "0000000011111100110101",
			4029 => "0000100110101100000100",
			4030 => "0000000011111100110101",
			4031 => "0000000011111100110101",
			4032 => "0001000001011100001000",
			4033 => "0001011101000100000100",
			4034 => "0000000011111100110101",
			4035 => "0000001011111100110101",
			4036 => "0000111000100000000100",
			4037 => "1111111011111100110101",
			4038 => "0011001001001000001000",
			4039 => "0000010100110100000100",
			4040 => "0000001011111100110101",
			4041 => "0000000011111100110101",
			4042 => "0001110101110100000100",
			4043 => "0000000011111100110101",
			4044 => "0000000011111100110101",
			4045 => "0000001010101101010000",
			4046 => "0011101100111001000100",
			4047 => "0000001011010100100100",
			4048 => "0010100010101100011000",
			4049 => "0000001001101000010000",
			4050 => "0010001000100100001000",
			4051 => "0001001100010000000100",
			4052 => "0000000011111111011001",
			4053 => "0000000011111111011001",
			4054 => "0011011010001000000100",
			4055 => "0000000011111111011001",
			4056 => "0000000011111111011001",
			4057 => "0001111001001000000100",
			4058 => "0000000011111111011001",
			4059 => "1111111011111111011001",
			4060 => "0001101101011000000100",
			4061 => "0000000011111111011001",
			4062 => "0010110000011100000100",
			4063 => "0000000011111111011001",
			4064 => "0000001011111111011001",
			4065 => "0011101000001100010000",
			4066 => "0001001011101100001000",
			4067 => "0011010101001000000100",
			4068 => "0000000011111111011001",
			4069 => "0000001011111111011001",
			4070 => "0001110001101000000100",
			4071 => "1111111011111111011001",
			4072 => "0000000011111111011001",
			4073 => "0000000111000100001100",
			4074 => "0000000110001000001000",
			4075 => "0010110110110100000100",
			4076 => "0000000011111111011001",
			4077 => "1111111011111111011001",
			4078 => "0000001011111111011001",
			4079 => "1111111011111111011001",
			4080 => "0011011100010100000100",
			4081 => "0000001011111111011001",
			4082 => "0010000001010100000100",
			4083 => "0000000011111111011001",
			4084 => "0000000011111111011001",
			4085 => "1111111011111111011001",
			4086 => "0010111011011101000100",
			4087 => "0011100111011000100100",
			4088 => "0000001100000100011100",
			4089 => "0010001000100100010100",
			4090 => "0001001100010000001100",
			4091 => "0000110111100000000100",
			4092 => "0000000100000011111101",
			4093 => "0000111100010000000100",
			4094 => "0000000100000011111101",
			4095 => "0000000100000011111101",
			4096 => "0010110101100100000100",
			4097 => "1111111100000011111101",
			4098 => "0000000100000011111101",
			4099 => "0000010000111100000100",
			4100 => "0000000100000011111101",
			4101 => "0000000100000011111101",
			4102 => "0001001010000100000100",
			4103 => "0000000100000011111101",
			4104 => "1111111100000011111101",
			4105 => "0010110101100100001000",
			4106 => "0000001111001000000100",
			4107 => "0000001100000011111101",
			4108 => "0000000100000011111101",
			4109 => "0001001111100100000100",
			4110 => "0000000100000011111101",
			4111 => "0010010111101100000100",
			4112 => "1111111100000011111101",
			4113 => "0010011010100000001000",
			4114 => "0010000110011100000100",
			4115 => "0000000100000011111101",
			4116 => "0000000100000011111101",
			4117 => "0011010101110000000100",
			4118 => "0000000100000011111101",
			4119 => "0000000100000011111101",
			4120 => "0001010111100000011000",
			4121 => "0000011101111100010000",
			4122 => "0010110010001000001100",
			4123 => "0001101101111100000100",
			4124 => "0000000100000011111101",
			4125 => "0000000010101000000100",
			4126 => "0000001100000011111101",
			4127 => "0000000100000011111101",
			4128 => "0000000100000011111101",
			4129 => "0001011100100100000100",
			4130 => "0000000100000011111101",
			4131 => "0000000100000011111101",
			4132 => "0011001011000000010000",
			4133 => "0011101100010000000100",
			4134 => "0000000100000011111101",
			4135 => "0000111101101100001000",
			4136 => "0011000100011000000100",
			4137 => "1111111100000011111101",
			4138 => "0000000100000011111101",
			4139 => "0000000100000011111101",
			4140 => "0000000001010100010000",
			4141 => "0000110110111100001000",
			4142 => "0011110010000100000100",
			4143 => "0000000100000011111101",
			4144 => "0000000100000011111101",
			4145 => "0001011111010000000100",
			4146 => "0000000100000011111101",
			4147 => "0000000100000011111101",
			4148 => "0011011100010100010000",
			4149 => "0011000110100100001000",
			4150 => "0000000111000000000100",
			4151 => "0000000100000011111101",
			4152 => "0000000100000011111101",
			4153 => "0001101010011000000100",
			4154 => "0000000100000011111101",
			4155 => "0000000100000011111101",
			4156 => "0010010100101100000100",
			4157 => "0000000100000011111101",
			4158 => "0000000100000011111101",
			4159 => "0011001010111000011000",
			4160 => "0000000110001000010100",
			4161 => "0001111001001000001000",
			4162 => "0000101111010100000100",
			4163 => "0000000100001000000001",
			4164 => "0000000100001000000001",
			4165 => "0010100111101100000100",
			4166 => "0000000100001000000001",
			4167 => "0001110110100100000100",
			4168 => "0000000100001000000001",
			4169 => "0000000100001000000001",
			4170 => "1111111100001000000001",
			4171 => "0001011100100100101100",
			4172 => "0000011101111100100000",
			4173 => "0011011110000100001100",
			4174 => "0000000001010100000100",
			4175 => "0000000100001000000001",
			4176 => "0001110001101000000100",
			4177 => "0000000100001000000001",
			4178 => "0000000100001000000001",
			4179 => "0000001111001000001000",
			4180 => "0001101101111100000100",
			4181 => "0000000100001000000001",
			4182 => "0000001100001000000001",
			4183 => "0010011010100000000100",
			4184 => "0000000100001000000001",
			4185 => "0000111101101100000100",
			4186 => "0000000100001000000001",
			4187 => "0000000100001000000001",
			4188 => "0011000100011000000100",
			4189 => "0000000100001000000001",
			4190 => "0011001000000000000100",
			4191 => "0000000100001000000001",
			4192 => "0000000100001000000001",
			4193 => "0001010111100000010000",
			4194 => "0011010111111100001100",
			4195 => "0000111111100100001000",
			4196 => "0011110110111100000100",
			4197 => "0000000100001000000001",
			4198 => "1111111100001000000001",
			4199 => "0000000100001000000001",
			4200 => "0000000100001000000001",
			4201 => "0000010000111100011000",
			4202 => "0000110110111100001000",
			4203 => "0010001000100100000100",
			4204 => "0000000100001000000001",
			4205 => "0000000100001000000001",
			4206 => "0001111000011000001000",
			4207 => "0001110001101000000100",
			4208 => "0000000100001000000001",
			4209 => "0000000100001000000001",
			4210 => "0000000001010100000100",
			4211 => "1111111100001000000001",
			4212 => "0000000100001000000001",
			4213 => "0011011100010100001100",
			4214 => "0000011010011000001000",
			4215 => "0001000101000000000100",
			4216 => "0000001100001000000001",
			4217 => "0000000100001000000001",
			4218 => "0000000100001000000001",
			4219 => "0001110000011100000100",
			4220 => "0000000100001000000001",
			4221 => "0000101101101100000100",
			4222 => "0000000100001000000001",
			4223 => "0000000100001000000001",
			4224 => "0000001010101101010100",
			4225 => "0011101100111001001000",
			4226 => "0000001011010100100100",
			4227 => "0010001000100100010000",
			4228 => "0001100100110100001100",
			4229 => "0001111111011100001000",
			4230 => "0001101101111100000100",
			4231 => "0000000100001010101101",
			4232 => "0000000100001010101101",
			4233 => "1111111100001010101101",
			4234 => "1111111100001010101101",
			4235 => "0000101100000000001000",
			4236 => "0011010001000000000100",
			4237 => "0000000100001010101101",
			4238 => "0000001100001010101101",
			4239 => "0001101011001100001000",
			4240 => "0000001001101000000100",
			4241 => "0000000100001010101101",
			4242 => "0000000100001010101101",
			4243 => "0000001100001010101101",
			4244 => "0011101000001100010100",
			4245 => "0001010010110100001000",
			4246 => "0010110000011100000100",
			4247 => "0000000100001010101101",
			4248 => "0000000100001010101101",
			4249 => "0001010001000000001000",
			4250 => "0001111001001000000100",
			4251 => "0000000100001010101101",
			4252 => "1111111100001010101101",
			4253 => "0000000100001010101101",
			4254 => "0000000111000100001100",
			4255 => "0000000110001000001000",
			4256 => "0010110110110100000100",
			4257 => "0000000100001010101101",
			4258 => "1111111100001010101101",
			4259 => "0000001100001010101101",
			4260 => "1111111100001010101101",
			4261 => "0011011010001000000100",
			4262 => "0000001100001010101101",
			4263 => "0010000001010100000100",
			4264 => "0000000100001010101101",
			4265 => "0000000100001010101101",
			4266 => "1111111100001010101101",
			4267 => "0011001010111000010000",
			4268 => "0000000110001000001100",
			4269 => "0011101100000000001000",
			4270 => "0001110110100100000100",
			4271 => "0000000100001110110001",
			4272 => "0000000100001110110001",
			4273 => "0000000100001110110001",
			4274 => "1111111100001110110001",
			4275 => "0001011100100100110000",
			4276 => "0000011101111100100100",
			4277 => "0001011101000100011000",
			4278 => "0000111010000100010000",
			4279 => "0000000001010100001000",
			4280 => "0011000100011000000100",
			4281 => "0000000100001110110001",
			4282 => "0000000100001110110001",
			4283 => "0011001010111000000100",
			4284 => "0000000100001110110001",
			4285 => "0000000100001110110001",
			4286 => "0000010001111000000100",
			4287 => "0000001100001110110001",
			4288 => "0000000100001110110001",
			4289 => "0001101101111100000100",
			4290 => "0000000100001110110001",
			4291 => "0000000001110100000100",
			4292 => "0000001100001110110001",
			4293 => "0000000100001110110001",
			4294 => "0011000100011000000100",
			4295 => "0000000100001110110001",
			4296 => "0011001000000000000100",
			4297 => "0000000100001110110001",
			4298 => "0000000100001110110001",
			4299 => "0001010111100000011100",
			4300 => "0011110110111100010000",
			4301 => "0001100100110100001000",
			4302 => "0000111100010000000100",
			4303 => "0000000100001110110001",
			4304 => "0000000100001110110001",
			4305 => "0011100110010000000100",
			4306 => "0000000100001110110001",
			4307 => "0000000100001110110001",
			4308 => "0000111111100100001000",
			4309 => "0010111011011100000100",
			4310 => "1111111100001110110001",
			4311 => "0000000100001110110001",
			4312 => "0000000100001110110001",
			4313 => "0000010000111100011000",
			4314 => "0000110110111100001000",
			4315 => "0010001000100100000100",
			4316 => "0000000100001110110001",
			4317 => "0000001100001110110001",
			4318 => "0001111000011000001000",
			4319 => "0001110001101000000100",
			4320 => "0000000100001110110001",
			4321 => "0000000100001110110001",
			4322 => "0011001001110100000100",
			4323 => "0000000100001110110001",
			4324 => "0000000100001110110001",
			4325 => "0000011010011000001100",
			4326 => "0001000101000000001000",
			4327 => "0001011110010000000100",
			4328 => "0000000100001110110001",
			4329 => "0000000100001110110001",
			4330 => "0000000100001110110001",
			4331 => "0000000100001110110001",
			4332 => "0011000111001000001000",
			4333 => "0001110110100100000100",
			4334 => "1111111100010010001101",
			4335 => "0000000100010010001101",
			4336 => "0000001001101000111000",
			4337 => "0010001000100100011000",
			4338 => "0001001100010000001100",
			4339 => "0000111100010000001000",
			4340 => "0010011111000000000100",
			4341 => "0000000100010010001101",
			4342 => "0000001100010010001101",
			4343 => "0000000100010010001101",
			4344 => "0000101110110100000100",
			4345 => "1111111100010010001101",
			4346 => "0011001000000000000100",
			4347 => "0000000100010010001101",
			4348 => "0000000100010010001101",
			4349 => "0011011010001000010000",
			4350 => "0011010101001000001000",
			4351 => "0000011110010100000100",
			4352 => "0000000100010010001101",
			4353 => "0000000100010010001101",
			4354 => "0000110000010000000100",
			4355 => "0000001100010010001101",
			4356 => "0000000100010010001101",
			4357 => "0001111111011100001000",
			4358 => "0000010000111100000100",
			4359 => "1111111100010010001101",
			4360 => "0000000100010010001101",
			4361 => "0001101100011000000100",
			4362 => "0000001100010010001101",
			4363 => "0000000100010010001101",
			4364 => "0010100010101100000100",
			4365 => "1111111100010010001101",
			4366 => "0000001011010100001100",
			4367 => "0001101101011000000100",
			4368 => "0000000100010010001101",
			4369 => "0000100111011000000100",
			4370 => "0000000100010010001101",
			4371 => "0000001100010010001101",
			4372 => "0011101000001100010000",
			4373 => "0001001011101100001000",
			4374 => "0011010101001000000100",
			4375 => "0000000100010010001101",
			4376 => "0000000100010010001101",
			4377 => "0001110001101000000100",
			4378 => "1111111100010010001101",
			4379 => "0000000100010010001101",
			4380 => "0000000010101000001000",
			4381 => "0000111100111000000100",
			4382 => "0000000100010010001101",
			4383 => "0000001100010010001101",
			4384 => "0000111000101000000100",
			4385 => "1111111100010010001101",
			4386 => "0000000100010010001101",
			4387 => "0010011001100100010100",
			4388 => "0001100000111100010000",
			4389 => "0001100000111100000100",
			4390 => "0000000100010110100001",
			4391 => "0000000011101000000100",
			4392 => "0000000100010110100001",
			4393 => "0000000000110000000100",
			4394 => "0000000100010110100001",
			4395 => "0000000100010110100001",
			4396 => "1111111100010110100001",
			4397 => "0011000100011001000000",
			4398 => "0000000110001000100000",
			4399 => "0001110110100100010000",
			4400 => "0001111001001000001000",
			4401 => "0011010001000000000100",
			4402 => "0000000100010110100001",
			4403 => "0000000100010110100001",
			4404 => "0010110000011100000100",
			4405 => "0000000100010110100001",
			4406 => "1111111100010110100001",
			4407 => "0011010100101000001100",
			4408 => "0010011111000000000100",
			4409 => "0000000100010110100001",
			4410 => "0011000100011000000100",
			4411 => "0000001100010110100001",
			4412 => "0000000100010110100001",
			4413 => "0000000100010110100001",
			4414 => "0010111011011100010000",
			4415 => "0001111000011000001100",
			4416 => "0010011010100000000100",
			4417 => "1111111100010110100001",
			4418 => "0010011010100000000100",
			4419 => "0000000100010110100001",
			4420 => "0000000100010110100001",
			4421 => "0000000100010110100001",
			4422 => "0011000100011000000100",
			4423 => "0000000100010110100001",
			4424 => "0011000100011000001000",
			4425 => "0000101110000000000100",
			4426 => "0000000100010110100001",
			4427 => "0000000100010110100001",
			4428 => "0000000100010110100001",
			4429 => "0011011100010100101000",
			4430 => "0000111011101100011100",
			4431 => "0000001111001000010000",
			4432 => "0001101011001100001000",
			4433 => "0000101000001100000100",
			4434 => "0000000100010110100001",
			4435 => "1111111100010110100001",
			4436 => "0000111111010100000100",
			4437 => "0000000100010110100001",
			4438 => "0000001100010110100001",
			4439 => "0011001000000000001000",
			4440 => "0011000100011000000100",
			4441 => "0000000100010110100001",
			4442 => "1111111100010110100001",
			4443 => "0000000100010110100001",
			4444 => "0000011010011000001000",
			4445 => "0000000111000000000100",
			4446 => "0000001100010110100001",
			4447 => "0000000100010110100001",
			4448 => "0000000100010110100001",
			4449 => "0010010100101100001100",
			4450 => "0000011011111100000100",
			4451 => "0000000100010110100001",
			4452 => "0011011110110100000100",
			4453 => "0000000100010110100001",
			4454 => "0000000100010110100001",
			4455 => "1111111100010110100001",
			4456 => "0011011110000100010100",
			4457 => "0000000101000100001100",
			4458 => "0001111011000000000100",
			4459 => "0000000100011010110101",
			4460 => "0001011101000100000100",
			4461 => "0000000100011010110101",
			4462 => "0000000100011010110101",
			4463 => "0001110110100100000100",
			4464 => "1111111100011010110101",
			4465 => "0000000100011010110101",
			4466 => "0010010111101101010000",
			4467 => "0001000000010000110000",
			4468 => "0011010010011100010100",
			4469 => "0011010101001000001100",
			4470 => "0011000100011000001000",
			4471 => "0001110110100100000100",
			4472 => "0000000100011010110101",
			4473 => "0000000100011010110101",
			4474 => "0000000100011010110101",
			4475 => "0010100000001000000100",
			4476 => "0000000100011010110101",
			4477 => "0000001100011010110101",
			4478 => "0000000001010100001100",
			4479 => "0001011111010000001000",
			4480 => "0000100110010000000100",
			4481 => "0000000100011010110101",
			4482 => "1111111100011010110101",
			4483 => "0000000100011010110101",
			4484 => "0000001100000100001000",
			4485 => "0011000100011000000100",
			4486 => "0000000100011010110101",
			4487 => "0000001100011010110101",
			4488 => "0000011011111100000100",
			4489 => "1111111100011010110101",
			4490 => "0000000100011010110101",
			4491 => "0011001000011000010100",
			4492 => "0001001101101100010000",
			4493 => "0010100010101100001000",
			4494 => "0001111111011100000100",
			4495 => "1111111100011010110101",
			4496 => "0000000100011010110101",
			4497 => "0001011110101000000100",
			4498 => "0000000100011010110101",
			4499 => "0000001100011010110101",
			4500 => "1111111100011010110101",
			4501 => "0000010001000100000100",
			4502 => "0000000100011010110101",
			4503 => "0001101000010000000100",
			4504 => "0000000100011010110101",
			4505 => "0000000100011010110101",
			4506 => "0000000001110100001100",
			4507 => "0010100011101000000100",
			4508 => "0000000100011010110101",
			4509 => "0001010111111100000100",
			4510 => "0000001100011010110101",
			4511 => "0000000100011010110101",
			4512 => "0011101100111000000100",
			4513 => "1111111100011010110101",
			4514 => "0001101000010000001000",
			4515 => "0010101000100100000100",
			4516 => "0000000100011010110101",
			4517 => "0000000100011010110101",
			4518 => "0011111011110000001000",
			4519 => "0000011010011000000100",
			4520 => "0000001100011010110101",
			4521 => "0000000100011010110101",
			4522 => "0011111110000000000100",
			4523 => "0000000100011010110101",
			4524 => "0000000100011010110101",
			4525 => "0000001010101101111000",
			4526 => "0000010000111100111000",
			4527 => "0001111000011000100000",
			4528 => "0001110001101000010100",
			4529 => "0001001100010000001100",
			4530 => "0001101101111100001000",
			4531 => "0001100000111100000100",
			4532 => "0000000100011110101001",
			4533 => "0000000100011110101001",
			4534 => "0000001100011110101001",
			4535 => "0010010100111100000100",
			4536 => "1111111100011110101001",
			4537 => "0000000100011110101001",
			4538 => "0000000101000100001000",
			4539 => "0000111100000000000100",
			4540 => "0000000100011110101001",
			4541 => "0000000100011110101001",
			4542 => "0000001100011110101001",
			4543 => "0000110110111100001000",
			4544 => "0010001000100100000100",
			4545 => "0000000100011110101001",
			4546 => "0000001100011110101001",
			4547 => "0000000001010100000100",
			4548 => "1111111100011110101001",
			4549 => "0001111000011000000100",
			4550 => "1111111100011110101001",
			4551 => "0010001000010100000100",
			4552 => "0000001100011110101001",
			4553 => "0000000100011110101001",
			4554 => "0001110001101000100100",
			4555 => "0001000001011100010100",
			4556 => "0001110001101000010000",
			4557 => "0001010110100000001000",
			4558 => "0000010111101000000100",
			4559 => "0000000100011110101001",
			4560 => "1111111100011110101001",
			4561 => "0011010101110000000100",
			4562 => "0000001100011110101001",
			4563 => "0000000100011110101001",
			4564 => "1111111100011110101001",
			4565 => "0000111111100100000100",
			4566 => "1111111100011110101001",
			4567 => "0000101101101100000100",
			4568 => "0000001100011110101001",
			4569 => "0010000101000100000100",
			4570 => "1111111100011110101001",
			4571 => "0000000100011110101001",
			4572 => "0001010111111100010000",
			4573 => "0000010000111100000100",
			4574 => "0000000100011110101001",
			4575 => "0001011101000100000100",
			4576 => "0000000100011110101001",
			4577 => "0011110110111000000100",
			4578 => "0000001100011110101001",
			4579 => "0000001100011110101001",
			4580 => "0001110101110100001000",
			4581 => "0001011110010000000100",
			4582 => "0000000100011110101001",
			4583 => "1111111100011110101001",
			4584 => "0000000100011110101001",
			4585 => "1111111100011110101001",
			4586 => "0001110110100100010100",
			4587 => "0001000111010100001100",
			4588 => "0000011011111100001000",
			4589 => "0000011101101000000100",
			4590 => "0000000100100011010101",
			4591 => "0000000100100011010101",
			4592 => "0000000100100011010101",
			4593 => "0000111010000100000100",
			4594 => "1111111100100011010101",
			4595 => "0000000100100011010101",
			4596 => "0001110001101000101100",
			4597 => "0001101011001100100000",
			4598 => "0001001011101100011100",
			4599 => "0010101010100000010000",
			4600 => "0001101101111100001000",
			4601 => "0011001011000000000100",
			4602 => "0000000100100011010101",
			4603 => "0000000100100011010101",
			4604 => "0011111001100000000100",
			4605 => "0000000100100011010101",
			4606 => "0000000100100011010101",
			4607 => "0010010100111100000100",
			4608 => "0000000100100011010101",
			4609 => "0000110110111100000100",
			4610 => "0000000100100011010101",
			4611 => "0000000100100011010101",
			4612 => "0000000100100011010101",
			4613 => "0000000001110100001000",
			4614 => "0000111000001100000100",
			4615 => "0000000100100011010101",
			4616 => "0000001100100011010101",
			4617 => "0000000100100011010101",
			4618 => "0001101100011000100100",
			4619 => "0000111010000100011000",
			4620 => "0000101110110100010000",
			4621 => "0001001100000000001000",
			4622 => "0000100010000000000100",
			4623 => "0000000100100011010101",
			4624 => "0000000100100011010101",
			4625 => "0011001011000000000100",
			4626 => "0000000100100011010101",
			4627 => "0000000100100011010101",
			4628 => "0001010001000000000100",
			4629 => "0000000100100011010101",
			4630 => "0000001100100011010101",
			4631 => "0000000001010100000100",
			4632 => "0000000100100011010101",
			4633 => "0011001011000000000100",
			4634 => "0000000100100011010101",
			4635 => "0000000100100011010101",
			4636 => "0001010111100000011100",
			4637 => "0001110001101000001100",
			4638 => "0011011111010000000100",
			4639 => "0000000100100011010101",
			4640 => "0011010100101000000100",
			4641 => "1111111100100011010101",
			4642 => "0000000100100011010101",
			4643 => "0001111000011000001000",
			4644 => "0001100100111100000100",
			4645 => "0000000100100011010101",
			4646 => "0000000100100011010101",
			4647 => "0011010101110000000100",
			4648 => "0000000100100011010101",
			4649 => "0000000100100011010101",
			4650 => "0011011010001000001000",
			4651 => "0000000010101000000100",
			4652 => "0000000100100011010101",
			4653 => "0000000100100011010101",
			4654 => "0011001001110100001000",
			4655 => "0001011001010000000100",
			4656 => "0000000100100011010101",
			4657 => "0000000100100011010101",
			4658 => "0000010000111100000100",
			4659 => "0000000100100011010101",
			4660 => "0000000100100011010101",
			4661 => "0000001010101101110000",
			4662 => "0010010111101101001100",
			4663 => "0000001100000100101100",
			4664 => "0000000001010100011000",
			4665 => "0011010101110000001100",
			4666 => "0001101101111100000100",
			4667 => "0000000100100110111001",
			4668 => "0000111100000000000100",
			4669 => "0000001100100110111001",
			4670 => "0000000100100110111001",
			4671 => "0001011111010000001000",
			4672 => "0011000100011000000100",
			4673 => "0000000100100110111001",
			4674 => "1111111100100110111001",
			4675 => "0000000100100110111001",
			4676 => "0001010110100000000100",
			4677 => "0000000100100110111001",
			4678 => "0000111000001100001000",
			4679 => "0010011111000000000100",
			4680 => "0000000100100110111001",
			4681 => "0000001100100110111001",
			4682 => "0010010100111100000100",
			4683 => "0000000100100110111001",
			4684 => "0000000100100110111001",
			4685 => "0001110111010000011100",
			4686 => "0010100010101100001100",
			4687 => "0001111001001000000100",
			4688 => "0000000100100110111001",
			4689 => "0011011110010000000100",
			4690 => "1111111100100110111001",
			4691 => "0000000100100110111001",
			4692 => "0001001011101100001000",
			4693 => "0001111001001000000100",
			4694 => "0000000100100110111001",
			4695 => "0000000100100110111001",
			4696 => "0001101001100100000100",
			4697 => "1111111100100110111001",
			4698 => "0000000100100110111001",
			4699 => "0000000100100110111001",
			4700 => "0000000001110100010000",
			4701 => "0001101011001100000100",
			4702 => "0000000100100110111001",
			4703 => "0000110111010100000100",
			4704 => "0000000100100110111001",
			4705 => "0001010111111100000100",
			4706 => "0000001100100110111001",
			4707 => "0000000100100110111001",
			4708 => "0011101100111000000100",
			4709 => "1111111100100110111001",
			4710 => "0001101000010000001000",
			4711 => "0001001011110000000100",
			4712 => "0000000100100110111001",
			4713 => "0000000100100110111001",
			4714 => "0001110000011100000100",
			4715 => "0000001100100110111001",
			4716 => "0000000100100110111001",
			4717 => "1111111100100110111001",
			4718 => "0000001010101101100100",
			4719 => "0001100100111101011000",
			4720 => "0000001001101000111000",
			4721 => "0001111000011000011100",
			4722 => "0001010110100000001100",
			4723 => "0000011011111100001000",
			4724 => "0001111011000000000100",
			4725 => "0000000100101010000101",
			4726 => "0000000100101010000101",
			4727 => "1111111100101010000101",
			4728 => "0010100000001000001000",
			4729 => "0011011111010000000100",
			4730 => "0000000100101010000101",
			4731 => "1111111100101010000101",
			4732 => "0011111010000100000100",
			4733 => "0000001100101010000101",
			4734 => "0000000100101010000101",
			4735 => "0001111000011000010000",
			4736 => "0010010100111100001000",
			4737 => "0000110110111100000100",
			4738 => "0000000100101010000101",
			4739 => "1111111100101010000101",
			4740 => "0000111000001100000100",
			4741 => "0000001100101010000101",
			4742 => "1111111100101010000101",
			4743 => "0010110100010000001000",
			4744 => "0010110010001000000100",
			4745 => "0000001100101010000101",
			4746 => "0000000100101010000101",
			4747 => "0000001100101010000101",
			4748 => "0011100111011000001100",
			4749 => "0000001001101000001000",
			4750 => "0000111110110100000100",
			4751 => "0000000100101010000101",
			4752 => "1111110100101010000101",
			4753 => "1111111100101010000101",
			4754 => "0001001000100000000100",
			4755 => "0000001100101010000101",
			4756 => "0011100111010100001000",
			4757 => "0001110110100100000100",
			4758 => "0000000100101010000101",
			4759 => "1111111100101010000101",
			4760 => "0000000111000100000100",
			4761 => "0000000100101010000101",
			4762 => "1111111100101010000101",
			4763 => "0010111010010100001000",
			4764 => "0001011110000100000100",
			4765 => "0000000100101010000101",
			4766 => "0000001100101010000101",
			4767 => "0000000100101010000101",
			4768 => "1111111100101010000101",
			4769 => "0011000111001000000100",
			4770 => "1111111100101110011011",
			4771 => "0001010111100000111100",
			4772 => "0001011100100100101000",
			4773 => "0001011100100100011000",
			4774 => "0000011101111100010000",
			4775 => "0001110110100100001000",
			4776 => "0000001111001000000100",
			4777 => "0000000100101110011011",
			4778 => "0000000100101110011011",
			4779 => "0001010110100000000100",
			4780 => "1111111100101110011011",
			4781 => "0000000100101110011011",
			4782 => "0011010101110000000100",
			4783 => "1111111100101110011011",
			4784 => "0000000100101110011011",
			4785 => "0010110110110100001100",
			4786 => "0000000001110100001000",
			4787 => "0001101101111100000100",
			4788 => "0000000100101110011011",
			4789 => "0000001100101110011011",
			4790 => "0000000100101110011011",
			4791 => "0000000100101110011011",
			4792 => "0011010010011100000100",
			4793 => "0000000100101110011011",
			4794 => "0000010001111000001100",
			4795 => "0010110010001000001000",
			4796 => "0000110111011000000100",
			4797 => "0000000100101110011011",
			4798 => "1111111100101110011011",
			4799 => "0000000100101110011011",
			4800 => "0000000100101110011011",
			4801 => "0001011111010000100000",
			4802 => "0000000101000100001100",
			4803 => "0011010101110000000100",
			4804 => "0000000100101110011011",
			4805 => "0001110001101000000100",
			4806 => "0000000100101110011011",
			4807 => "0000000100101110011011",
			4808 => "0000010100110100001100",
			4809 => "0001000111011000000100",
			4810 => "0000000100101110011011",
			4811 => "0011011010001000000100",
			4812 => "0000001100101110011011",
			4813 => "0000000100101110011011",
			4814 => "0011011010001000000100",
			4815 => "0000000100101110011011",
			4816 => "0000000100101110011011",
			4817 => "0000010000111100010000",
			4818 => "0000101100000000001000",
			4819 => "0001000110111100000100",
			4820 => "0000000100101110011011",
			4821 => "0000000100101110011011",
			4822 => "0001111111011100000100",
			4823 => "1111111100101110011011",
			4824 => "0000000100101110011011",
			4825 => "0011011100010100001100",
			4826 => "0000001010101100001000",
			4827 => "0010110100010000000100",
			4828 => "0000000100101110011011",
			4829 => "0000001100101110011011",
			4830 => "0000000100101110011011",
			4831 => "0011001000011000001000",
			4832 => "0001010011001000000100",
			4833 => "0000000100101110011011",
			4834 => "0000000100101110011011",
			4835 => "0000010111101000000100",
			4836 => "0000000100101110011011",
			4837 => "0000000100101110011011",
			4838 => "0000000100101110011101",
			4839 => "0000000100101110100001",
			4840 => "0011001011000000000100",
			4841 => "0000000100101110110101",
			4842 => "0011000110100100000100",
			4843 => "0000000100101110110101",
			4844 => "0000000100101110110101",
			4845 => "0010110100010000001000",
			4846 => "0010110000011100000100",
			4847 => "0000000100101111001001",
			4848 => "0000000100101111001001",
			4849 => "0000000100101111001001",
			4850 => "0000001100000100001000",
			4851 => "0001000110110100000100",
			4852 => "0000000100101111011101",
			4853 => "0000000100101111011101",
			4854 => "0000000100101111011101",
			4855 => "0000001100000100001000",
			4856 => "0000000011101000000100",
			4857 => "0000000100101111110001",
			4858 => "0000000100101111110001",
			4859 => "0000000100101111110001",
			4860 => "0001011100100100001000",
			4861 => "0001010110110100000100",
			4862 => "0000000100110000001101",
			4863 => "0000000100110000001101",
			4864 => "0001011111010000000100",
			4865 => "0000000100110000001101",
			4866 => "0000000100110000001101",
			4867 => "0010111011011100000100",
			4868 => "0000000100110000101001",
			4869 => "0000101100000000001000",
			4870 => "0000100010000000000100",
			4871 => "0000000100110000101001",
			4872 => "0000000100110000101001",
			4873 => "0000000100110000101001",
			4874 => "0000101100010000001100",
			4875 => "0001000111010100001000",
			4876 => "0000101101000100000100",
			4877 => "0000000100110001001101",
			4878 => "0000000100110001001101",
			4879 => "0000000100110001001101",
			4880 => "0000101010000100000100",
			4881 => "0000000100110001001101",
			4882 => "0000000100110001001101",
			4883 => "0000001001101000001100",
			4884 => "0000101101000100000100",
			4885 => "0000000100110001110001",
			4886 => "0000101010000100000100",
			4887 => "0000000100110001110001",
			4888 => "0000000100110001110001",
			4889 => "0000101000101000000100",
			4890 => "0000000100110001110001",
			4891 => "0000000100110001110001",
			4892 => "0000001100000100001100",
			4893 => "0000101100000000001000",
			4894 => "0000101110110100000100",
			4895 => "0000000100110010011101",
			4896 => "0000000100110010011101",
			4897 => "0000000100110010011101",
			4898 => "0001101000010000001000",
			4899 => "0001100100110100000100",
			4900 => "0000000100110010011101",
			4901 => "0000000100110010011101",
			4902 => "0000000100110010011101",
			4903 => "0000000001110100010000",
			4904 => "0001011100100100001100",
			4905 => "0001110001101000001000",
			4906 => "0001111011000000000100",
			4907 => "0000000100110011000001",
			4908 => "0000000100110011000001",
			4909 => "0000000100110011000001",
			4910 => "0000000100110011000001",
			4911 => "0000000100110011000001",
			4912 => "0011001001110100010000",
			4913 => "0001001100010000000100",
			4914 => "0000000100110011100101",
			4915 => "0001101011001100001000",
			4916 => "0011001010111000000100",
			4917 => "0000000100110011100101",
			4918 => "0000000100110011100101",
			4919 => "0000000100110011100101",
			4920 => "0000000100110011100101",
			4921 => "0010011111000000001000",
			4922 => "0010101001100100000100",
			4923 => "0000000100110100010001",
			4924 => "0000000100110100010001",
			4925 => "0010101001000100001100",
			4926 => "0010100000001000000100",
			4927 => "0000000100110100010001",
			4928 => "0010010010101100000100",
			4929 => "0000000100110100010001",
			4930 => "0000000100110100010001",
			4931 => "0000000100110100010001",
			4932 => "0010111011011100000100",
			4933 => "0000000100110100111101",
			4934 => "0001011111010000001000",
			4935 => "0001011100100100000100",
			4936 => "0000000100110100111101",
			4937 => "0000000100110100111101",
			4938 => "0010111011110100001000",
			4939 => "0010110010001000000100",
			4940 => "0000000100110100111101",
			4941 => "0000000100110100111101",
			4942 => "0000000100110100111101",
			4943 => "0010010111101100001100",
			4944 => "0010011111000000001000",
			4945 => "0010011111000000000100",
			4946 => "0000000100110101110001",
			4947 => "0000000100110101110001",
			4948 => "0000000100110101110001",
			4949 => "0001010111111100001100",
			4950 => "0010010010101100001000",
			4951 => "0001010010110100000100",
			4952 => "0000000100110101110001",
			4953 => "0000000100110101110001",
			4954 => "0000000100110101110001",
			4955 => "0000000100110101110001",
			4956 => "0011000100011000001000",
			4957 => "0010010000001000000100",
			4958 => "0000000100110110100101",
			4959 => "0000000100110110100101",
			4960 => "0010111011011100000100",
			4961 => "0000000100110110100101",
			4962 => "0001001101101100001100",
			4963 => "0011111110110100000100",
			4964 => "0000000100110110100101",
			4965 => "0000011001011000000100",
			4966 => "0000000100110110100101",
			4967 => "0000000100110110100101",
			4968 => "0000000100110110100101",
			4969 => "0000000001110100010100",
			4970 => "0001011100100100010000",
			4971 => "0010011010100000001100",
			4972 => "0001010110110100000100",
			4973 => "0000000100110111010001",
			4974 => "0000001111001000000100",
			4975 => "0000000100110111010001",
			4976 => "0000000100110111010001",
			4977 => "0000000100110111010001",
			4978 => "0000000100110111010001",
			4979 => "0000000100110111010001",
			4980 => "0011001001110100010100",
			4981 => "0001001100010000000100",
			4982 => "0000000100110111111101",
			4983 => "0001101011001100001100",
			4984 => "0011001010111000000100",
			4985 => "0000000100110111111101",
			4986 => "0001111001001000000100",
			4987 => "0000000100110111111101",
			4988 => "0000000100110111111101",
			4989 => "0000000100110111111101",
			4990 => "0000000100110111111101",
			4991 => "0000001001101000010100",
			4992 => "0011110111011000000100",
			4993 => "0000000100111001000001",
			4994 => "0000000001010100000100",
			4995 => "0000000100111001000001",
			4996 => "0011000110100100001000",
			4997 => "0010110101100100000100",
			4998 => "0000000100111001000001",
			4999 => "0000000100111001000001",
			5000 => "0000000100111001000001",
			5001 => "0011100111010100000100",
			5002 => "0000000100111001000001",
			5003 => "0010000101000100001000",
			5004 => "0010000001010000000100",
			5005 => "0000000100111001000001",
			5006 => "0000000100111001000001",
			5007 => "0000000100111001000001",
			5008 => "0011001001110100010000",
			5009 => "0001001100010000000100",
			5010 => "0000000100111010000101",
			5011 => "0011101100111000001000",
			5012 => "0010110101100100000100",
			5013 => "0000000100111010000101",
			5014 => "0000000100111010000101",
			5015 => "0000000100111010000101",
			5016 => "0000100110111000010000",
			5017 => "0000000001010100000100",
			5018 => "0000000100111010000101",
			5019 => "0010110010001000000100",
			5020 => "0000000100111010000101",
			5021 => "0011010010000100000100",
			5022 => "0000000100111010000101",
			5023 => "0000000100111010000101",
			5024 => "0000000100111010000101",
			5025 => "0000000111000100011000",
			5026 => "0010011111000000000100",
			5027 => "0000000100111011000001",
			5028 => "0011011110000100000100",
			5029 => "0000000100111011000001",
			5030 => "0011011010001000001100",
			5031 => "0010100000001000000100",
			5032 => "0000000100111011000001",
			5033 => "0001110110100100000100",
			5034 => "0000000100111011000001",
			5035 => "0000000100111011000001",
			5036 => "0000000100111011000001",
			5037 => "0001101000010000000100",
			5038 => "0000000100111011000001",
			5039 => "0000000100111011000001",
			5040 => "0001000001011100011000",
			5041 => "0010100000001000000100",
			5042 => "0000000100111011111101",
			5043 => "0000011101111100010000",
			5044 => "0000011001011000000100",
			5045 => "0000000100111011111101",
			5046 => "0010110000011100000100",
			5047 => "0000000100111011111101",
			5048 => "0010001100011100000100",
			5049 => "0000000100111011111101",
			5050 => "0000000100111011111101",
			5051 => "0000000100111011111101",
			5052 => "0001100100111100000100",
			5053 => "0000000100111011111101",
			5054 => "0000000100111011111101",
			5055 => "0011101100000000001000",
			5056 => "0011011001010100000100",
			5057 => "0000000100111100111001",
			5058 => "0000000100111100111001",
			5059 => "0011010011001000010100",
			5060 => "0010010100111100000100",
			5061 => "0000000100111100111001",
			5062 => "0011100010010100001100",
			5063 => "0011011110000100000100",
			5064 => "0000000100111100111001",
			5065 => "0010010010101100000100",
			5066 => "0000000100111100111001",
			5067 => "0000000100111100111001",
			5068 => "0000000100111100111001",
			5069 => "0000000100111100111001",
			5070 => "0001101101111100001000",
			5071 => "0011000100011000000100",
			5072 => "0000000100111101110101",
			5073 => "0000000100111101110101",
			5074 => "0001111000011000010100",
			5075 => "0001011100100100000100",
			5076 => "0000000100111101110101",
			5077 => "0011001001110100001100",
			5078 => "0010011010100100001000",
			5079 => "0011010010011100000100",
			5080 => "0000000100111101110101",
			5081 => "0000000100111101110101",
			5082 => "0000000100111101110101",
			5083 => "0000000100111101110101",
			5084 => "0000000100111101110101",
			5085 => "0000000001110100011000",
			5086 => "0001011100100100010100",
			5087 => "0010011010100000010000",
			5088 => "0001010110100000000100",
			5089 => "0000000100111110101001",
			5090 => "0010011111000000000100",
			5091 => "0000000100111110101001",
			5092 => "0000001111001000000100",
			5093 => "0000000100111110101001",
			5094 => "0000000100111110101001",
			5095 => "0000000100111110101001",
			5096 => "0000000100111110101001",
			5097 => "0000000100111110101001",
			5098 => "0001011111010000011000",
			5099 => "0011000100011000000100",
			5100 => "0000000100111111011101",
			5101 => "0000000010101000010000",
			5102 => "0011001001001000001100",
			5103 => "0001110110100100000100",
			5104 => "0000000100111111011101",
			5105 => "0001111111011100000100",
			5106 => "0000000100111111011101",
			5107 => "0000000100111111011101",
			5108 => "0000000100111111011101",
			5109 => "0000000100111111011101",
			5110 => "0000000100111111011101",
			5111 => "0000010000111100010000",
			5112 => "0011101110110100000100",
			5113 => "0000000101000000101001",
			5114 => "0001010101110000001000",
			5115 => "0011010101110000000100",
			5116 => "0000000101000000101001",
			5117 => "0000000101000000101001",
			5118 => "0000000101000000101001",
			5119 => "0011000100011000000100",
			5120 => "0000000101000000101001",
			5121 => "0000000001110100010000",
			5122 => "0011101100000000000100",
			5123 => "0000000101000000101001",
			5124 => "0000010100110100001000",
			5125 => "0001010110100000000100",
			5126 => "0000000101000000101001",
			5127 => "0000000101000000101001",
			5128 => "0000000101000000101001",
			5129 => "0000000101000000101001",
			5130 => "0001000111010100010100",
			5131 => "0010001000100100000100",
			5132 => "0000000101000010001101",
			5133 => "0011111111010100001100",
			5134 => "0011000111001000000100",
			5135 => "0000000101000010001101",
			5136 => "0011110110010000000100",
			5137 => "0000000101000010001101",
			5138 => "0000000101000010001101",
			5139 => "0000000101000010001101",
			5140 => "0001100100111100010000",
			5141 => "0001110000011100001100",
			5142 => "0010001000010100000100",
			5143 => "0000000101000010001101",
			5144 => "0001101111000000000100",
			5145 => "0000000101000010001101",
			5146 => "0000000101000010001101",
			5147 => "0000000101000010001101",
			5148 => "0000001010101100001100",
			5149 => "0000011010011000001000",
			5150 => "0010011010100000000100",
			5151 => "0000000101000010001101",
			5152 => "0000000101000010001101",
			5153 => "0000000101000010001101",
			5154 => "0000000101000010001101",
			5155 => "0000001100000100011000",
			5156 => "0010100000001000010000",
			5157 => "0010000111110100000100",
			5158 => "0000000101000011111001",
			5159 => "0001100100110100001000",
			5160 => "0011111001100000000100",
			5161 => "0000000101000011111001",
			5162 => "0000000101000011111001",
			5163 => "0000000101000011111001",
			5164 => "0011110110010000000100",
			5165 => "0000000101000011111001",
			5166 => "0000000101000011111001",
			5167 => "0010100010101100001100",
			5168 => "0010110101110100001000",
			5169 => "0001101101111100000100",
			5170 => "0000000101000011111001",
			5171 => "0000000101000011111001",
			5172 => "0000000101000011111001",
			5173 => "0010101000100100010000",
			5174 => "0000101101101100001100",
			5175 => "0010000101000100001000",
			5176 => "0000101100000000000100",
			5177 => "0000000101000011111001",
			5178 => "0000000101000011111001",
			5179 => "0000000101000011111001",
			5180 => "0000000101000011111001",
			5181 => "0000000101000011111001",
			5182 => "0001000001011100100000",
			5183 => "0010001000100100001000",
			5184 => "0000011001011000000100",
			5185 => "0000000101000101001101",
			5186 => "0000000101000101001101",
			5187 => "0001110110100100000100",
			5188 => "0000000101000101001101",
			5189 => "0000011001011000000100",
			5190 => "0000000101000101001101",
			5191 => "0001111000011000001100",
			5192 => "0000010111101000001000",
			5193 => "0011010001000000000100",
			5194 => "0000000101000101001101",
			5195 => "0000000101000101001101",
			5196 => "0000000101000101001101",
			5197 => "0000000101000101001101",
			5198 => "0000011100011000001000",
			5199 => "0001110001011000000100",
			5200 => "0000000101000101001101",
			5201 => "0000000101000101001101",
			5202 => "0000000101000101001101",
			5203 => "0010111011011100001100",
			5204 => "0011100111011000001000",
			5205 => "0000111010000100000100",
			5206 => "0000000101000110011001",
			5207 => "0000000101000110011001",
			5208 => "0000000101000110011001",
			5209 => "0001001101101100011000",
			5210 => "0001110110100100000100",
			5211 => "0000000101000110011001",
			5212 => "0000011001011000000100",
			5213 => "0000000101000110011001",
			5214 => "0000000101000100000100",
			5215 => "0000000101000110011001",
			5216 => "0001000111011000000100",
			5217 => "0000000101000110011001",
			5218 => "0000101110110100000100",
			5219 => "0000000101000110011001",
			5220 => "0000000101000110011001",
			5221 => "0000000101000110011001",
			5222 => "0001001101101100011100",
			5223 => "0000011001011000000100",
			5224 => "0000000101000111011101",
			5225 => "0011011110000100000100",
			5226 => "0000000101000111011101",
			5227 => "0000111000100000010000",
			5228 => "0010011111000000000100",
			5229 => "0000000101000111011101",
			5230 => "0011111100000000000100",
			5231 => "0000000101000111011101",
			5232 => "0000011101111100000100",
			5233 => "0000000101000111011101",
			5234 => "0000000101000111011101",
			5235 => "0000000101000111011101",
			5236 => "0010011010100000000100",
			5237 => "0000000101000111011101",
			5238 => "0000000101000111011101",
			5239 => "0011111100000000001100",
			5240 => "0010101010100000001000",
			5241 => "0001110110100100000100",
			5242 => "0000000101001001001001",
			5243 => "0000000101001001001001",
			5244 => "0000000101001001001001",
			5245 => "0011001000000000011000",
			5246 => "0010100010101100001100",
			5247 => "0001111000011000001000",
			5248 => "0011001010111000000100",
			5249 => "0000000101001001001001",
			5250 => "0000000101001001001001",
			5251 => "0000000101001001001001",
			5252 => "0010101000100100001000",
			5253 => "0001111001001000000100",
			5254 => "0000000101001001001001",
			5255 => "0000000101001001001001",
			5256 => "0000000101001001001001",
			5257 => "0011000110100100010000",
			5258 => "0011011100010100001100",
			5259 => "0000010000111100000100",
			5260 => "0000000101001001001001",
			5261 => "0000000111000000000100",
			5262 => "0000000101001001001001",
			5263 => "0000000101001001001001",
			5264 => "0000000101001001001001",
			5265 => "0000000101001001001001",
			5266 => "0001010110100000001000",
			5267 => "0011100111010100000100",
			5268 => "0000000101001010101101",
			5269 => "0000000101001010101101",
			5270 => "0010011001111100011000",
			5271 => "0000101100010000001100",
			5272 => "0011100110010000000100",
			5273 => "0000000101001010101101",
			5274 => "0000100110010000000100",
			5275 => "0000000101001010101101",
			5276 => "0000000101001010101101",
			5277 => "0011101010000100001000",
			5278 => "0000101100000000000100",
			5279 => "0000000101001010101101",
			5280 => "0000000101001010101101",
			5281 => "0000000101001010101101",
			5282 => "0000100110111000010000",
			5283 => "0010010010101100001100",
			5284 => "0011101100010000000100",
			5285 => "0000000101001010101101",
			5286 => "0001111001001000000100",
			5287 => "0000000101001010101101",
			5288 => "0000000101001010101101",
			5289 => "0000000101001010101101",
			5290 => "0000000101001010101101",
			5291 => "0010011111000000001100",
			5292 => "0001101101111100000100",
			5293 => "0000000101001100000001",
			5294 => "0010100000001000000100",
			5295 => "0000000101001100000001",
			5296 => "0000000101001100000001",
			5297 => "0000000001110100011100",
			5298 => "0001110110100100000100",
			5299 => "0000000101001100000001",
			5300 => "0011001001001000010000",
			5301 => "0011011010001000001100",
			5302 => "0001011001010000001000",
			5303 => "0010001000100100000100",
			5304 => "0000000101001100000001",
			5305 => "0000000101001100000001",
			5306 => "0000000101001100000001",
			5307 => "0000000101001100000001",
			5308 => "0011001001110100000100",
			5309 => "0000000101001100000001",
			5310 => "0000000101001100000001",
			5311 => "0000000101001100000001",
			5312 => "0011100111010100011100",
			5313 => "0010110101110100011000",
			5314 => "0001000110010000000100",
			5315 => "0000000101001100111101",
			5316 => "0010100010101100010000",
			5317 => "0001111001001000000100",
			5318 => "0000000101001100111101",
			5319 => "0001011111010000001000",
			5320 => "0001111111011100000100",
			5321 => "0000000101001100111101",
			5322 => "0000000101001100111101",
			5323 => "0000000101001100111101",
			5324 => "0000000101001100111101",
			5325 => "0000000101001100111101",
			5326 => "0000000101001100111101",
			5327 => "0010011111000000000100",
			5328 => "0000000101001101111001",
			5329 => "0001000101000000011000",
			5330 => "0011000100011000000100",
			5331 => "0000000101001101111001",
			5332 => "0001011110010000010000",
			5333 => "0010100000001000000100",
			5334 => "0000000101001101111001",
			5335 => "0010010010101100001000",
			5336 => "0010110100000100000100",
			5337 => "0000000101001101111001",
			5338 => "0000000101001101111001",
			5339 => "0000000101001101111001",
			5340 => "0000000101001101111001",
			5341 => "0000000101001101111001",
			5342 => "0000000010101000011100",
			5343 => "0010011111000000000100",
			5344 => "0000000101001110110101",
			5345 => "0001110110100100000100",
			5346 => "0000000101001110110101",
			5347 => "0000000001010100000100",
			5348 => "0000000101001110110101",
			5349 => "0000011010011000001100",
			5350 => "0011001010111000000100",
			5351 => "0000000101001110110101",
			5352 => "0000010000111100000100",
			5353 => "0000000101001110110101",
			5354 => "0000000101001110110101",
			5355 => "0000000101001110110101",
			5356 => "0000000101001110110101",
			5357 => "0010011111000000000100",
			5358 => "0000000101010000000001",
			5359 => "0001001111100100011000",
			5360 => "0001011111010000010100",
			5361 => "0011011010001000010000",
			5362 => "0011001001001000001100",
			5363 => "0001110110100100000100",
			5364 => "0000000101010000000001",
			5365 => "0010100000001000000100",
			5366 => "0000000101010000000001",
			5367 => "0000000101010000000001",
			5368 => "0000000101010000000001",
			5369 => "0000000101010000000001",
			5370 => "0000000101010000000001",
			5371 => "0010010111101100001000",
			5372 => "0001101101011000000100",
			5373 => "0000000101010000000001",
			5374 => "0000000101010000000001",
			5375 => "0000000101010000000001",
			5376 => "0001001111100100011000",
			5377 => "0011111110110100000100",
			5378 => "0000000101010001110101",
			5379 => "0000110000010000010000",
			5380 => "0001100100110100000100",
			5381 => "0000000101010001110101",
			5382 => "0001110110100100000100",
			5383 => "0000000101010001110101",
			5384 => "0010100011101000000100",
			5385 => "0000000101010001110101",
			5386 => "0000000101010001110101",
			5387 => "0000000101010001110101",
			5388 => "0000111111100100010000",
			5389 => "0011001010111000000100",
			5390 => "0000000101010001110101",
			5391 => "0001010010110100000100",
			5392 => "0000000101010001110101",
			5393 => "0001010111100000000100",
			5394 => "0000000101010001110101",
			5395 => "0000000101010001110101",
			5396 => "0000010001000100000100",
			5397 => "0000000101010001110101",
			5398 => "0011111110000000001100",
			5399 => "0000011010011000001000",
			5400 => "0010101001000100000100",
			5401 => "0000000101010001110101",
			5402 => "0000000101010001110101",
			5403 => "0000000101010001110101",
			5404 => "0000000101010001110101",
			5405 => "0001001011101100110000",
			5406 => "0011010101110000011000",
			5407 => "0001110110100100000100",
			5408 => "0000000101010100000001",
			5409 => "0010011111000000000100",
			5410 => "0000000101010100000001",
			5411 => "0010110110110100001100",
			5412 => "0010100000001000000100",
			5413 => "0000000101010100000001",
			5414 => "0011011110000100000100",
			5415 => "0000000101010100000001",
			5416 => "0000000101010100000001",
			5417 => "0000000101010100000001",
			5418 => "0010110110110100001100",
			5419 => "0000110000010000001000",
			5420 => "0011111001100000000100",
			5421 => "0000000101010100000001",
			5422 => "0000000101010100000001",
			5423 => "0000000101010100000001",
			5424 => "0000110111010100001000",
			5425 => "0011111100000000000100",
			5426 => "0000000101010100000001",
			5427 => "0000000101010100000001",
			5428 => "0000000101010100000001",
			5429 => "0000111111100100001100",
			5430 => "0011101000001100001000",
			5431 => "0000001011010100000100",
			5432 => "0000000101010100000001",
			5433 => "0000000101010100000001",
			5434 => "0000000101010100000001",
			5435 => "0000000111000100001000",
			5436 => "0000001011010100000100",
			5437 => "0000000101010100000001",
			5438 => "0000000101010100000001",
			5439 => "0000000101010100000001",
			5440 => "0000000001110100101000",
			5441 => "0010011111000000001000",
			5442 => "0001111000011000000100",
			5443 => "1111111101010110000101",
			5444 => "0000001101010110000101",
			5445 => "0011010001000000001000",
			5446 => "0000100110010000000100",
			5447 => "0000010101010110000101",
			5448 => "1111111101010110000101",
			5449 => "0011010110010000010100",
			5450 => "0010000101000100001100",
			5451 => "0001101101111100000100",
			5452 => "1111111101010110000101",
			5453 => "0001000001011100000100",
			5454 => "0000010101010110000101",
			5455 => "0000010101010110000101",
			5456 => "0001000110111000000100",
			5457 => "0000010101010110000101",
			5458 => "0000101101010110000101",
			5459 => "1111111101010110000101",
			5460 => "0000001010101100010100",
			5461 => "0010000001010100001100",
			5462 => "0010000001010100000100",
			5463 => "1111111101010110000101",
			5464 => "0001001000000100000100",
			5465 => "0000001101010110000101",
			5466 => "1111111101010110000101",
			5467 => "0001101000010000000100",
			5468 => "1111111101010110000101",
			5469 => "0000100101010110000101",
			5470 => "0000001010101100000100",
			5471 => "1111111101010110000101",
			5472 => "1111111101010110000101",
			5473 => "0010010100111100010100",
			5474 => "0010101010100000001100",
			5475 => "0000110111010100001000",
			5476 => "0000110111100000000100",
			5477 => "0000000101011000010001",
			5478 => "0000000101011000010001",
			5479 => "0000000101011000010001",
			5480 => "0000010000111100000100",
			5481 => "0000000101011000010001",
			5482 => "0000000101011000010001",
			5483 => "0011111111010100010000",
			5484 => "0000001001101000001100",
			5485 => "0011011010001000001000",
			5486 => "0011010111100000000100",
			5487 => "0000000101011000010001",
			5488 => "0000000101011000010001",
			5489 => "0000000101011000010001",
			5490 => "0000000101011000010001",
			5491 => "0000111010000100001100",
			5492 => "0011111010000100001000",
			5493 => "0001011110101000000100",
			5494 => "0000000101011000010001",
			5495 => "0000000101011000010001",
			5496 => "0000000101011000010001",
			5497 => "0000000001110100010000",
			5498 => "0000001001101000000100",
			5499 => "0000000101011000010001",
			5500 => "0001011101000100000100",
			5501 => "0000000101011000010001",
			5502 => "0010010101010000000100",
			5503 => "0000000101011000010001",
			5504 => "0000000101011000010001",
			5505 => "0000111000101000000100",
			5506 => "0000000101011000010001",
			5507 => "0000000101011000010001",
			5508 => "0001001101101100101000",
			5509 => "0011111010000100100100",
			5510 => "0001110001101000010100",
			5511 => "0001001100010000000100",
			5512 => "0000000101011001111101",
			5513 => "0011010111111100001100",
			5514 => "0001111001001000000100",
			5515 => "0000000101011001111101",
			5516 => "0010110000011100000100",
			5517 => "0000000101011001111101",
			5518 => "0000000101011001111101",
			5519 => "0000000101011001111101",
			5520 => "0000000101000100000100",
			5521 => "0000000101011001111101",
			5522 => "0010011111000000000100",
			5523 => "0000000101011001111101",
			5524 => "0001111111011100000100",
			5525 => "0000000101011001111101",
			5526 => "0000000101011001111101",
			5527 => "0000000101011001111101",
			5528 => "0010011010100000001100",
			5529 => "0011001011011100001000",
			5530 => "0010000001010000000100",
			5531 => "0000000101011001111101",
			5532 => "0000000101011001111101",
			5533 => "0000000101011001111101",
			5534 => "0000000101011001111101",
			5535 => "0001001011101100101100",
			5536 => "0010110101100100010100",
			5537 => "0000101111010100010000",
			5538 => "0010010101010000000100",
			5539 => "0000000101011100010001",
			5540 => "0011001101010100000100",
			5541 => "0000000101011100010001",
			5542 => "0011011110000100000100",
			5543 => "0000000101011100010001",
			5544 => "0000000101011100010001",
			5545 => "0000000101011100010001",
			5546 => "0011010101001000000100",
			5547 => "0000000101011100010001",
			5548 => "0000011001011000000100",
			5549 => "0000000101011100010001",
			5550 => "0000101000001100001100",
			5551 => "0011011010001000001000",
			5552 => "0010001000100100000100",
			5553 => "0000000101011100010001",
			5554 => "0000000101011100010001",
			5555 => "0000000101011100010001",
			5556 => "0000000101011100010001",
			5557 => "0001101001100100001100",
			5558 => "0011001001110100001000",
			5559 => "0000001011010100000100",
			5560 => "0000000101011100010001",
			5561 => "0000000101011100010001",
			5562 => "0000000101011100010001",
			5563 => "0000000001110100001100",
			5564 => "0000101101101100001000",
			5565 => "0011110110101100000100",
			5566 => "0000000101011100010001",
			5567 => "0000000101011100010001",
			5568 => "0000000101011100010001",
			5569 => "0010000001110000000100",
			5570 => "0000000101011100010001",
			5571 => "0000000101011100010001",
			5572 => "0001001011101100110000",
			5573 => "0001111000011000011000",
			5574 => "0011001010111000000100",
			5575 => "0000000101011110000101",
			5576 => "0010010111101100010000",
			5577 => "0000011001011000000100",
			5578 => "0000000101011110000101",
			5579 => "0011001001001000001000",
			5580 => "0010110111010000000100",
			5581 => "0000000101011110000101",
			5582 => "0000000101011110000101",
			5583 => "0000000101011110000101",
			5584 => "0000000101011110000101",
			5585 => "0010110100010000010100",
			5586 => "0001011001010000010000",
			5587 => "0001011100100100000100",
			5588 => "0000000101011110000101",
			5589 => "0011000100011000000100",
			5590 => "0000000101011110000101",
			5591 => "0011001001110100000100",
			5592 => "0000000101011110000101",
			5593 => "0000000101011110000101",
			5594 => "0000000101011110000101",
			5595 => "0000000101011110000101",
			5596 => "0011001001110100001000",
			5597 => "0001100100111100000100",
			5598 => "0000000101011110000101",
			5599 => "0000000101011110000101",
			5600 => "0000000101011110000101",
			5601 => "0011010101110000011000",
			5602 => "0000001111001000010000",
			5603 => "0010011111000000000100",
			5604 => "0000000101100000011001",
			5605 => "0010110110110100001000",
			5606 => "0011010001000000000100",
			5607 => "0000000101100000011001",
			5608 => "0000000101100000011001",
			5609 => "0000000101100000011001",
			5610 => "0000111000100000000100",
			5611 => "0000000101100000011001",
			5612 => "0000000101100000011001",
			5613 => "0001010111100000001100",
			5614 => "0010000001010000001000",
			5615 => "0011000100011000000100",
			5616 => "0000000101100000011001",
			5617 => "0000000101100000011001",
			5618 => "0000000101100000011001",
			5619 => "0011011010001000010100",
			5620 => "0011000100011000000100",
			5621 => "0000000101100000011001",
			5622 => "0000101110110100000100",
			5623 => "0000000101100000011001",
			5624 => "0010110101110100001000",
			5625 => "0000001010101100000100",
			5626 => "0000000101100000011001",
			5627 => "0000000101100000011001",
			5628 => "0000000101100000011001",
			5629 => "0000111011111000000100",
			5630 => "0000000101100000011001",
			5631 => "0011001000011000001100",
			5632 => "0001011111010000000100",
			5633 => "0000000101100000011001",
			5634 => "0001010011001000000100",
			5635 => "0000000101100000011001",
			5636 => "0000000101100000011001",
			5637 => "0000000101100000011001",
			5638 => "0001101101111100010000",
			5639 => "0011000100011000000100",
			5640 => "0000000101100010100101",
			5641 => "0011001001110100001000",
			5642 => "0000010000111100000100",
			5643 => "0000000101100010100101",
			5644 => "0000000101100010100101",
			5645 => "0000000101100010100101",
			5646 => "0001111000011000100000",
			5647 => "0010010100101100010100",
			5648 => "0001011100100100000100",
			5649 => "0000000101100010100101",
			5650 => "0011011001011100001100",
			5651 => "0011000100011000000100",
			5652 => "0000000101100010100101",
			5653 => "0011010010011100000100",
			5654 => "0000000101100010100101",
			5655 => "0000000101100010100101",
			5656 => "0000000101100010100101",
			5657 => "0000011101111100001000",
			5658 => "0001111000000000000100",
			5659 => "0000000101100010100101",
			5660 => "0000000101100010100101",
			5661 => "0000000101100010100101",
			5662 => "0011001011000000000100",
			5663 => "0000000101100010100101",
			5664 => "0011010110010000010000",
			5665 => "0011000001101000001100",
			5666 => "0011011100010100001000",
			5667 => "0001100101010000000100",
			5668 => "0000000101100010100101",
			5669 => "0000000101100010100101",
			5670 => "0000000101100010100101",
			5671 => "0000000101100010100101",
			5672 => "0000000101100010100101",
			5673 => "0000000010101000111100",
			5674 => "0000011001011000010000",
			5675 => "0001100000111100001000",
			5676 => "0011111010011100000100",
			5677 => "1111111101100100111001",
			5678 => "0000001101100100111001",
			5679 => "0010011111000000000100",
			5680 => "1111111101100100111001",
			5681 => "0000000101100100111001",
			5682 => "0011010110010000100100",
			5683 => "0011011110000100001100",
			5684 => "0000000001010100000100",
			5685 => "0000001101100100111001",
			5686 => "0001011101000100000100",
			5687 => "1111111101100100111001",
			5688 => "0000000101100100111001",
			5689 => "0010100000001000001100",
			5690 => "0000110010000100001000",
			5691 => "0010000111110100000100",
			5692 => "0000000101100100111001",
			5693 => "0000000101100100111001",
			5694 => "1111111101100100111001",
			5695 => "0001100100111100001000",
			5696 => "0000000110001000000100",
			5697 => "0000001101100100111001",
			5698 => "0000000101100100111001",
			5699 => "0000010101100100111001",
			5700 => "0001110100010000000100",
			5701 => "1111111101100100111001",
			5702 => "0000000101100100111001",
			5703 => "0000001010101100001100",
			5704 => "0010000001010100000100",
			5705 => "1111111101100100111001",
			5706 => "0001101000010000000100",
			5707 => "0000000101100100111001",
			5708 => "0000001101100100111001",
			5709 => "1111111101100100111001",
			5710 => "0011111100000000001100",
			5711 => "0010010100111100001000",
			5712 => "0000010000111100000100",
			5713 => "0000000101100111000101",
			5714 => "0000000101100111000101",
			5715 => "0000000101100111000101",
			5716 => "0011001000000000100100",
			5717 => "0001101011001100010100",
			5718 => "0001111000011000010000",
			5719 => "0001011110101000000100",
			5720 => "0000000101100111000101",
			5721 => "0001101101111100000100",
			5722 => "0000000101100111000101",
			5723 => "0011000100011000000100",
			5724 => "0000000101100111000101",
			5725 => "0000000101100111000101",
			5726 => "0000000101100111000101",
			5727 => "0001110001101000001100",
			5728 => "0000000001110100001000",
			5729 => "0001111001001000000100",
			5730 => "0000000101100111000101",
			5731 => "0000000101100111000101",
			5732 => "0000000101100111000101",
			5733 => "0000000101100111000101",
			5734 => "0011010110010000010100",
			5735 => "0000011001011000000100",
			5736 => "0000000101100111000101",
			5737 => "0011000110100100001100",
			5738 => "0011011100010100001000",
			5739 => "0011101110110100000100",
			5740 => "0000000101100111000101",
			5741 => "0000000101100111000101",
			5742 => "0000000101100111000101",
			5743 => "0000000101100111000101",
			5744 => "0000000101100111000101",
			5745 => "0010011001111100101100",
			5746 => "0000001100000100100100",
			5747 => "0010101010100000011100",
			5748 => "0011010101110000010000",
			5749 => "0001010111100000001100",
			5750 => "0000011101101000000100",
			5751 => "0000000101101001111001",
			5752 => "0000111100000000000100",
			5753 => "0000000101101001111001",
			5754 => "0000000101101001111001",
			5755 => "0000000101101001111001",
			5756 => "0011010111111100001000",
			5757 => "0000100110010000000100",
			5758 => "0000000101101001111001",
			5759 => "0000000101101001111001",
			5760 => "0000000101101001111001",
			5761 => "0000010000111100000100",
			5762 => "0000000101101001111001",
			5763 => "0000000101101001111001",
			5764 => "0011001000011000000100",
			5765 => "0000000101101001111001",
			5766 => "0000000101101001111001",
			5767 => "0000001111001000001100",
			5768 => "0000110110111100000100",
			5769 => "0000000101101001111001",
			5770 => "0001010110100000000100",
			5771 => "0000000101101001111001",
			5772 => "0000001101101001111001",
			5773 => "0011101100111000010000",
			5774 => "0001111000011000001100",
			5775 => "0011001010111000000100",
			5776 => "0000000101101001111001",
			5777 => "0001101000010000000100",
			5778 => "0000000101101001111001",
			5779 => "0000000101101001111001",
			5780 => "0000000101101001111001",
			5781 => "0001001000110100010000",
			5782 => "0011000100011000000100",
			5783 => "0000000101101001111001",
			5784 => "0011010101110000000100",
			5785 => "0000000101101001111001",
			5786 => "0010010010101100000100",
			5787 => "0000000101101001111001",
			5788 => "0000000101101001111001",
			5789 => "0000000101101001111001",
			5790 => "0011010101110000100000",
			5791 => "0000001111001000011000",
			5792 => "0010011111000000000100",
			5793 => "0000000101101100011101",
			5794 => "0001110110100100000100",
			5795 => "0000000101101100011101",
			5796 => "0010110110110100001100",
			5797 => "0011010001000000000100",
			5798 => "0000000101101100011101",
			5799 => "0001010001000000000100",
			5800 => "0000000101101100011101",
			5801 => "0000000101101100011101",
			5802 => "0000000101101100011101",
			5803 => "0000111000100000000100",
			5804 => "0000000101101100011101",
			5805 => "0000000101101100011101",
			5806 => "0001010111100000001100",
			5807 => "0010000001010000001000",
			5808 => "0011000100011000000100",
			5809 => "0000000101101100011101",
			5810 => "0000000101101100011101",
			5811 => "0000000101101100011101",
			5812 => "0011011010001000010100",
			5813 => "0011000100011000000100",
			5814 => "0000000101101100011101",
			5815 => "0000000001010100000100",
			5816 => "0000000101101100011101",
			5817 => "0000001010101100001000",
			5818 => "0011000110100100000100",
			5819 => "0000000101101100011101",
			5820 => "0000000101101100011101",
			5821 => "0000000101101100011101",
			5822 => "0000111000100000000100",
			5823 => "0000000101101100011101",
			5824 => "0011001000011000001100",
			5825 => "0001011111010000000100",
			5826 => "0000000101101100011101",
			5827 => "0001010011001000000100",
			5828 => "0000000101101100011101",
			5829 => "0000000101101100011101",
			5830 => "0000000101101100011101",
			5831 => "0000000010101000111100",
			5832 => "0010011001100100001100",
			5833 => "0001100000111100001000",
			5834 => "0000010111100100000100",
			5835 => "1111111101101110101001",
			5836 => "0000001101101110101001",
			5837 => "1111111101101110101001",
			5838 => "0001010110100000001000",
			5839 => "0000011011111100000100",
			5840 => "0000001101101110101001",
			5841 => "1111111101101110101001",
			5842 => "0001010101110000011000",
			5843 => "0001100100111100010000",
			5844 => "0011001010111000001000",
			5845 => "0000000110001000000100",
			5846 => "0000001101101110101001",
			5847 => "1111111101101110101001",
			5848 => "0010100000001000000100",
			5849 => "0000000101101110101001",
			5850 => "0000001101101110101001",
			5851 => "0001011001010000000100",
			5852 => "0000010101101110101001",
			5853 => "0000001101101110101001",
			5854 => "0001001101101100000100",
			5855 => "0000001101101110101001",
			5856 => "0001110101110100001000",
			5857 => "0001110000011100000100",
			5858 => "1111111101101110101001",
			5859 => "1111111101101110101001",
			5860 => "0000001101101110101001",
			5861 => "0000001010101100001000",
			5862 => "0001101000010000000100",
			5863 => "1111111101101110101001",
			5864 => "0000001101101110101001",
			5865 => "1111111101101110101001",
			5866 => "0001001000001100100100",
			5867 => "0011001010111000000100",
			5868 => "0000000101110001011101",
			5869 => "0001111000011000010000",
			5870 => "0000011011111100001100",
			5871 => "0000011001011000000100",
			5872 => "0000000101110001011101",
			5873 => "0010011111000000000100",
			5874 => "0000000101110001011101",
			5875 => "0000000101110001011101",
			5876 => "0000000101110001011101",
			5877 => "0000000001010100001000",
			5878 => "0000000101000100000100",
			5879 => "0000000101110001011101",
			5880 => "0000000101110001011101",
			5881 => "0000000001010100000100",
			5882 => "0000000101110001011101",
			5883 => "0000000101110001011101",
			5884 => "0000111010000100010000",
			5885 => "0011001011000000001100",
			5886 => "0001110001101000001000",
			5887 => "0011101111010100000100",
			5888 => "1111111101110001011101",
			5889 => "0000000101110001011101",
			5890 => "0000000101110001011101",
			5891 => "0000000101110001011101",
			5892 => "0000101000001100001000",
			5893 => "0000010000111100000100",
			5894 => "0000000101110001011101",
			5895 => "0000000101110001011101",
			5896 => "0011100111010100001100",
			5897 => "0011001011000000001000",
			5898 => "0001110110100100000100",
			5899 => "0000000101110001011101",
			5900 => "0000000101110001011101",
			5901 => "0000000101110001011101",
			5902 => "0000101011111000000100",
			5903 => "0000000101110001011101",
			5904 => "0010110101110100001000",
			5905 => "0001111000011000000100",
			5906 => "0000000101110001011101",
			5907 => "0000000101110001011101",
			5908 => "0011001000011000000100",
			5909 => "0000000101110001011101",
			5910 => "0000000101110001011101",
			5911 => "0010010100101100111000",
			5912 => "0000001100000100101000",
			5913 => "0000111010000100011100",
			5914 => "0010100000001000010100",
			5915 => "0001001100010000001100",
			5916 => "0001011100100100001000",
			5917 => "0011000100011000000100",
			5918 => "0000000101110100101001",
			5919 => "0000000101110100101001",
			5920 => "0000000101110100101001",
			5921 => "0001000111011000000100",
			5922 => "0000000101110100101001",
			5923 => "0000000101110100101001",
			5924 => "0010011111000000000100",
			5925 => "0000000101110100101001",
			5926 => "0000000101110100101001",
			5927 => "0011001001001000001000",
			5928 => "0010001000010100000100",
			5929 => "0000000101110100101001",
			5930 => "0000000101110100101001",
			5931 => "0000000101110100101001",
			5932 => "0011001000011000001100",
			5933 => "0010001000010100000100",
			5934 => "0000000101110100101001",
			5935 => "0010101010100000000100",
			5936 => "0000000101110100101001",
			5937 => "0000000101110100101001",
			5938 => "0000000101110100101001",
			5939 => "0010100010101100001000",
			5940 => "0010010100101100000100",
			5941 => "0000000101110100101001",
			5942 => "0000000101110100101001",
			5943 => "0000000001110100011100",
			5944 => "0001011101000100010000",
			5945 => "0001110110100100001000",
			5946 => "0001111001001000000100",
			5947 => "0000000101110100101001",
			5948 => "0000000101110100101001",
			5949 => "0001001011101100000100",
			5950 => "0000000101110100101001",
			5951 => "0000000101110100101001",
			5952 => "0000110010010100001000",
			5953 => "0010010010101100000100",
			5954 => "0000000101110100101001",
			5955 => "0000000101110100101001",
			5956 => "0000000101110100101001",
			5957 => "0000111000101000001000",
			5958 => "0010000001010100000100",
			5959 => "0000000101110100101001",
			5960 => "0000000101110100101001",
			5961 => "0000000101110100101001",
			5962 => "0000000010101001000100",
			5963 => "0000011001011000010100",
			5964 => "0010101001100100001100",
			5965 => "0000100001101000000100",
			5966 => "0000000101110111011101",
			5967 => "0010011110010100000100",
			5968 => "0000001101110111011101",
			5969 => "0000000101110111011101",
			5970 => "0010011111000000000100",
			5971 => "1111111101110111011101",
			5972 => "0000000101110111011101",
			5973 => "0000001111001000011000",
			5974 => "0010001100011100010000",
			5975 => "0000011101111100001100",
			5976 => "0000111000100000001000",
			5977 => "0011010101110000000100",
			5978 => "0000001101110111011101",
			5979 => "0000000101110111011101",
			5980 => "0000000101110111011101",
			5981 => "1111110101110111011101",
			5982 => "0000111000001100000100",
			5983 => "0000000101110111011101",
			5984 => "0000001101110111011101",
			5985 => "0000111111100100000100",
			5986 => "1111111101110111011101",
			5987 => "0011011010001000001000",
			5988 => "0010111011011100000100",
			5989 => "0000000101110111011101",
			5990 => "0000001101110111011101",
			5991 => "0010101000010100001000",
			5992 => "0001000010010100000100",
			5993 => "0000000101110111011101",
			5994 => "1111111101110111011101",
			5995 => "0000001101110111011101",
			5996 => "0000001010101100010100",
			5997 => "0000001010101100000100",
			5998 => "1111111101110111011101",
			5999 => "0000011010011000001100",
			6000 => "0010010010101100000100",
			6001 => "0000000101110111011101",
			6002 => "0000011100011000000100",
			6003 => "0000000101110111011101",
			6004 => "0000000101110111011101",
			6005 => "0000000101110111011101",
			6006 => "1111111101110111011101",
			6007 => "0000000001110101000000",
			6008 => "0010011111000000010100",
			6009 => "0000011001011000010000",
			6010 => "0001100000111100001000",
			6011 => "0000010111100100000100",
			6012 => "1111111101111010100001",
			6013 => "0000101101111010100001",
			6014 => "0010110010001000000100",
			6015 => "1111111101111010100001",
			6016 => "0000000101111010100001",
			6017 => "0000001101111010100001",
			6018 => "0001010110100000001100",
			6019 => "0000110111010100001000",
			6020 => "0000011011111100000100",
			6021 => "0000001101111010100001",
			6022 => "1111111101111010100001",
			6023 => "0000010101111010100001",
			6024 => "0000110010010100011100",
			6025 => "0000011001011000001100",
			6026 => "0010100000001000001000",
			6027 => "0001011100100100000100",
			6028 => "0000010101111010100001",
			6029 => "1111111101111010100001",
			6030 => "0000001101111010100001",
			6031 => "0000001111001000001000",
			6032 => "0010011111000000000100",
			6033 => "0000011101111010100001",
			6034 => "0000001101111010100001",
			6035 => "0000111111100100000100",
			6036 => "1111111101111010100001",
			6037 => "0000001101111010100001",
			6038 => "1111111101111010100001",
			6039 => "0000000010101000010000",
			6040 => "0010000001010100001100",
			6041 => "0001001011110000001000",
			6042 => "0010000101000100000100",
			6043 => "1111111101111010100001",
			6044 => "0000001101111010100001",
			6045 => "1111111101111010100001",
			6046 => "0000011101111010100001",
			6047 => "0000001010101100010000",
			6048 => "0010000001110000001100",
			6049 => "0001101000010000000100",
			6050 => "1111111101111010100001",
			6051 => "0010000001010100000100",
			6052 => "1111111101111010100001",
			6053 => "0000000101111010100001",
			6054 => "0000010101111010100001",
			6055 => "1111111101111010100001",
			6056 => "0010011001111100110100",
			6057 => "0000001100000100101100",
			6058 => "0010101010100000011100",
			6059 => "0011010101110000010000",
			6060 => "0010110110110100001100",
			6061 => "0000011101101000000100",
			6062 => "0000000101111101100101",
			6063 => "0000111100000000000100",
			6064 => "0000000101111101100101",
			6065 => "0000000101111101100101",
			6066 => "0000000101111101100101",
			6067 => "0011010111111100001000",
			6068 => "0010011111000000000100",
			6069 => "0000000101111101100101",
			6070 => "0000000101111101100101",
			6071 => "0000000101111101100101",
			6072 => "0000111000001100001100",
			6073 => "0001110110100100000100",
			6074 => "0000000101111101100101",
			6075 => "0011111001100000000100",
			6076 => "0000000101111101100101",
			6077 => "0000000101111101100101",
			6078 => "0000000101111101100101",
			6079 => "0011001000011000000100",
			6080 => "0000000101111101100101",
			6081 => "0000000101111101100101",
			6082 => "0000000111000100011000",
			6083 => "0000110110111100000100",
			6084 => "0000000101111101100101",
			6085 => "0011000100011000001100",
			6086 => "0011001010111000001000",
			6087 => "0011000111001000000100",
			6088 => "0000000101111101100101",
			6089 => "0000000101111101100101",
			6090 => "0000000101111101100101",
			6091 => "0011011110000100000100",
			6092 => "0000000101111101100101",
			6093 => "0000001101111101100101",
			6094 => "0000111100111000000100",
			6095 => "0000000101111101100101",
			6096 => "0001001000110100010000",
			6097 => "0001100100111100000100",
			6098 => "0000000101111101100101",
			6099 => "0001001011110000000100",
			6100 => "0000000101111101100101",
			6101 => "0000110110111000000100",
			6102 => "0000000101111101100101",
			6103 => "0000000101111101100101",
			6104 => "0000000101111101100101",
			6105 => "0000000010101001000000",
			6106 => "0000111100111000110000",
			6107 => "0000000111000100101000",
			6108 => "0010010111101100100000",
			6109 => "0011111111010100010000",
			6110 => "0000011001011000001000",
			6111 => "0001100100110100000100",
			6112 => "0000000101111111110001",
			6113 => "0000000101111111110001",
			6114 => "0010110100010000000100",
			6115 => "0000000101111111110001",
			6116 => "0000000101111111110001",
			6117 => "0011001011000000001000",
			6118 => "0010010100101100000100",
			6119 => "1111111101111111110001",
			6120 => "0000000101111111110001",
			6121 => "0000010001000100000100",
			6122 => "0000000101111111110001",
			6123 => "0000000101111111110001",
			6124 => "0000111010000100000100",
			6125 => "0000000101111111110001",
			6126 => "0000001101111111110001",
			6127 => "0011000100011000000100",
			6128 => "0000000101111111110001",
			6129 => "1111111101111111110001",
			6130 => "0000101101101100000100",
			6131 => "0000001101111111110001",
			6132 => "0011011110010000000100",
			6133 => "0000000101111111110001",
			6134 => "0000100011000000000100",
			6135 => "0000000101111111110001",
			6136 => "0000000101111111110001",
			6137 => "0010010010101100000100",
			6138 => "1111111101111111110001",
			6139 => "0000000101111111110001",
			6140 => "0000000001110101000000",
			6141 => "0010011111000000010000",
			6142 => "0010110010001000001100",
			6143 => "0001100000111100001000",
			6144 => "0000010111100100000100",
			6145 => "1111111110000010100101",
			6146 => "0000001110000010100101",
			6147 => "1111111110000010100101",
			6148 => "0000000110000010100101",
			6149 => "0010110100000100001000",
			6150 => "0000101001100000000100",
			6151 => "0000000110000010100101",
			6152 => "1111111110000010100101",
			6153 => "0011011100010100100000",
			6154 => "0000010000111100010000",
			6155 => "0001111000011000001000",
			6156 => "0001010111100000000100",
			6157 => "0000001110000010100101",
			6158 => "1111111110000010100101",
			6159 => "0010110100010000000100",
			6160 => "0000001110000010100101",
			6161 => "0000010110000010100101",
			6162 => "0000001111001000001000",
			6163 => "0011010111100000000100",
			6164 => "0000000110000010100101",
			6165 => "0000001110000010100101",
			6166 => "0000111111100100000100",
			6167 => "1111111110000010100101",
			6168 => "0000001110000010100101",
			6169 => "0000001111001000000100",
			6170 => "0000000110000010100101",
			6171 => "1111111110000010100101",
			6172 => "0000001010101100011000",
			6173 => "0010000001010100010000",
			6174 => "0000000001110100001100",
			6175 => "0000010100110100001000",
			6176 => "0000110110010000000100",
			6177 => "0000000110000010100101",
			6178 => "0000010110000010100101",
			6179 => "1111111110000010100101",
			6180 => "1111111110000010100101",
			6181 => "0001101000010000000100",
			6182 => "0000000110000010100101",
			6183 => "0000001110000010100101",
			6184 => "1111111110000010100101",
			6185 => "0001001111100101000000",
			6186 => "0010101010100000100000",
			6187 => "0011010101110000001000",
			6188 => "0010011111000000000100",
			6189 => "0000000110000110011001",
			6190 => "0000000110000110011001",
			6191 => "0000100010000100001100",
			6192 => "0010001000100100001000",
			6193 => "0011000100011000000100",
			6194 => "0000000110000110011001",
			6195 => "1111111110000110011001",
			6196 => "0000000110000110011001",
			6197 => "0000110111010100001000",
			6198 => "0011001000000000000100",
			6199 => "0000000110000110011001",
			6200 => "0000000110000110011001",
			6201 => "0000000110000110011001",
			6202 => "0000111011111000011000",
			6203 => "0011011110000100001000",
			6204 => "0000001100000100000100",
			6205 => "0000000110000110011001",
			6206 => "0000000110000110011001",
			6207 => "0000010000111100000100",
			6208 => "0000000110000110011001",
			6209 => "0000010111101000001000",
			6210 => "0000111100000000000100",
			6211 => "0000000110000110011001",
			6212 => "0000001110000110011001",
			6213 => "0000000110000110011001",
			6214 => "0010111011110100000100",
			6215 => "0000000110000110011001",
			6216 => "0000000110000110011001",
			6217 => "0000010111101000010100",
			6218 => "0011001001110100001100",
			6219 => "0010000110011000000100",
			6220 => "0000000110000110011001",
			6221 => "0010010100101100000100",
			6222 => "1111111110000110011001",
			6223 => "0000000110000110011001",
			6224 => "0010001100011100000100",
			6225 => "0000000110000110011001",
			6226 => "0000000110000110011001",
			6227 => "0000000110001000001000",
			6228 => "0000111000001100000100",
			6229 => "0000000110000110011001",
			6230 => "0000001110000110011001",
			6231 => "0000111111100100001000",
			6232 => "0010110000011100000100",
			6233 => "0000000110000110011001",
			6234 => "1111111110000110011001",
			6235 => "0000000111000100001000",
			6236 => "0000011100011000000100",
			6237 => "0000000110000110011001",
			6238 => "0000000110000110011001",
			6239 => "0011101100111000001000",
			6240 => "0000000001110100000100",
			6241 => "0000000110000110011001",
			6242 => "1111111110000110011001",
			6243 => "0001101000010000000100",
			6244 => "0000000110000110011001",
			6245 => "0000000110000110011001",
			6246 => "0001001011101101000000",
			6247 => "0010100010101100111000",
			6248 => "0000011110010100110000",
			6249 => "0001110001101000011100",
			6250 => "0001001100010000001100",
			6251 => "0000111100010000001000",
			6252 => "0011001101010100000100",
			6253 => "0000000110001001011101",
			6254 => "0000000110001001011101",
			6255 => "0000000110001001011101",
			6256 => "0001101010011000001000",
			6257 => "0010110101100100000100",
			6258 => "0000000110001001011101",
			6259 => "0000000110001001011101",
			6260 => "0000100010000100000100",
			6261 => "0000000110001001011101",
			6262 => "0000000110001001011101",
			6263 => "0001111000011000001000",
			6264 => "0000011001011000000100",
			6265 => "0000000110001001011101",
			6266 => "0000000110001001011101",
			6267 => "0000010000111100001000",
			6268 => "0000011001011000000100",
			6269 => "0000000110001001011101",
			6270 => "0000000110001001011101",
			6271 => "0000000110001001011101",
			6272 => "0011000100011000000100",
			6273 => "0000000110001001011101",
			6274 => "0000000110001001011101",
			6275 => "0000110110111100000100",
			6276 => "0000000110001001011101",
			6277 => "0000000110001001011101",
			6278 => "0001101111000000001100",
			6279 => "0000001011010100000100",
			6280 => "0000000110001001011101",
			6281 => "0011001000011000000100",
			6282 => "0000000110001001011101",
			6283 => "0000000110001001011101",
			6284 => "0000000001110100010000",
			6285 => "0001110110100100000100",
			6286 => "0000000110001001011101",
			6287 => "0010111011110100001000",
			6288 => "0000111011111000000100",
			6289 => "0000000110001001011101",
			6290 => "0000000110001001011101",
			6291 => "0000000110001001011101",
			6292 => "0001101000010000000100",
			6293 => "0000000110001001011101",
			6294 => "0000000110001001011101",
			6295 => "0001001111100101000100",
			6296 => "0010101010100000100100",
			6297 => "0011010101110000001000",
			6298 => "0010011111000000000100",
			6299 => "0000000110001101000001",
			6300 => "0000000110001101000001",
			6301 => "0000100010000100001100",
			6302 => "0010001000100100001000",
			6303 => "0011000100011000000100",
			6304 => "0000000110001101000001",
			6305 => "1111111110001101000001",
			6306 => "0000000110001101000001",
			6307 => "0000111010000100001000",
			6308 => "0011001000000000000100",
			6309 => "0000000110001101000001",
			6310 => "0000000110001101000001",
			6311 => "0010110100010000000100",
			6312 => "0000000110001101000001",
			6313 => "0000000110001101000001",
			6314 => "0000111011111000011000",
			6315 => "0011011111010000010000",
			6316 => "0011000100011000001000",
			6317 => "0010101010100000000100",
			6318 => "0000000110001101000001",
			6319 => "0000000110001101000001",
			6320 => "0011000100011000000100",
			6321 => "0000000110001101000001",
			6322 => "0000000110001101000001",
			6323 => "0000010000111100000100",
			6324 => "0000000110001101000001",
			6325 => "0000001110001101000001",
			6326 => "0010111011110100000100",
			6327 => "0000000110001101000001",
			6328 => "0000000110001101000001",
			6329 => "0011100111010100001000",
			6330 => "0010110110110100000100",
			6331 => "1111111110001101000001",
			6332 => "0000000110001101000001",
			6333 => "0001001101101100000100",
			6334 => "0000001110001101000001",
			6335 => "0000011110010100001000",
			6336 => "0011001000011000000100",
			6337 => "1111111110001101000001",
			6338 => "0000000110001101000001",
			6339 => "0000111000101000010000",
			6340 => "0000000111000100001000",
			6341 => "0000101111100100000100",
			6342 => "0000000110001101000001",
			6343 => "0000000110001101000001",
			6344 => "0011101100111000000100",
			6345 => "1111111110001101000001",
			6346 => "0000000110001101000001",
			6347 => "0011111110000000001000",
			6348 => "0000001010101100000100",
			6349 => "0000001110001101000001",
			6350 => "0000000110001101000001",
			6351 => "0000000110001101000001",
			6352 => "0010010111101101010000",
			6353 => "0000001001101000111100",
			6354 => "0011010010011100010000",
			6355 => "0011010101001000001000",
			6356 => "0010010101010000000100",
			6357 => "0000000110010000111101",
			6358 => "0000000110010000111101",
			6359 => "0010011111000000000100",
			6360 => "0000000110010000111101",
			6361 => "0000001110010000111101",
			6362 => "0010110110110100010000",
			6363 => "0010110101100100000100",
			6364 => "0000000110010000111101",
			6365 => "0010100010101100001000",
			6366 => "0000100110010000000100",
			6367 => "0000000110010000111101",
			6368 => "1111111110010000111101",
			6369 => "0000000110010000111101",
			6370 => "0001100100110100010000",
			6371 => "0000011001011000001000",
			6372 => "0010110010001000000100",
			6373 => "0000000110010000111101",
			6374 => "0000000110010000111101",
			6375 => "0011001001110100000100",
			6376 => "0000000110010000111101",
			6377 => "0000000110010000111101",
			6378 => "0000111011111000001000",
			6379 => "0010011111000000000100",
			6380 => "0000000110010000111101",
			6381 => "0000000110010000111101",
			6382 => "0000000110010000111101",
			6383 => "0011000001101000001000",
			6384 => "0000010001111000000100",
			6385 => "0000000110010000111101",
			6386 => "0000000110010000111101",
			6387 => "0000010001000100000100",
			6388 => "0000000110010000111101",
			6389 => "0000010111101000000100",
			6390 => "0000000110010000111101",
			6391 => "0000000110010000111101",
			6392 => "0000000111000100010000",
			6393 => "0001101011001100000100",
			6394 => "0000000110010000111101",
			6395 => "0000110111010100000100",
			6396 => "0000000110010000111101",
			6397 => "0010110101110100000100",
			6398 => "0000001110010000111101",
			6399 => "0000000110010000111101",
			6400 => "0011101100111000001100",
			6401 => "0011000100011000000100",
			6402 => "0000000110010000111101",
			6403 => "0000110011000000000100",
			6404 => "0000000110010000111101",
			6405 => "0000000110010000111101",
			6406 => "0011111110000000010000",
			6407 => "0001101000010000000100",
			6408 => "0000000110010000111101",
			6409 => "0011000100011000000100",
			6410 => "0000000110010000111101",
			6411 => "0000111101101100000100",
			6412 => "0000000110010000111101",
			6413 => "0000000110010000111101",
			6414 => "0000000110010000111101",
			6415 => "0001110110100100010100",
			6416 => "0001000111010100001100",
			6417 => "0000011011111100001000",
			6418 => "0000011101101000000100",
			6419 => "0000000110010100100001",
			6420 => "0000000110010100100001",
			6421 => "0000000110010100100001",
			6422 => "0001101011001100000100",
			6423 => "1111111110010100100001",
			6424 => "0000000110010100100001",
			6425 => "0001110001101000101000",
			6426 => "0001101011001100011100",
			6427 => "0001001011101100011000",
			6428 => "0010101010100000001100",
			6429 => "0001101101111100000100",
			6430 => "0000000110010100100001",
			6431 => "0011111001100000000100",
			6432 => "0000000110010100100001",
			6433 => "0000000110010100100001",
			6434 => "0010010100111100000100",
			6435 => "0000000110010100100001",
			6436 => "0000110110111100000100",
			6437 => "0000000110010100100001",
			6438 => "0000000110010100100001",
			6439 => "0000000110010100100001",
			6440 => "0000000001110100001000",
			6441 => "0000111000001100000100",
			6442 => "0000000110010100100001",
			6443 => "0000001110010100100001",
			6444 => "0000000110010100100001",
			6445 => "0010111011011100010000",
			6446 => "0010110101100100000100",
			6447 => "0000000110010100100001",
			6448 => "0000110000010000001000",
			6449 => "0011111001100000000100",
			6450 => "0000000110010100100001",
			6451 => "1111111110010100100001",
			6452 => "0000000110010100100001",
			6453 => "0001001101101100010100",
			6454 => "0000010000111100010000",
			6455 => "0000111010000100001000",
			6456 => "0011001001110100000100",
			6457 => "0000000110010100100001",
			6458 => "0000000110010100100001",
			6459 => "0001111111011100000100",
			6460 => "0000000110010100100001",
			6461 => "0000000110010100100001",
			6462 => "0000001110010100100001",
			6463 => "0000111101101100001000",
			6464 => "0001010111100000000100",
			6465 => "0000000110010100100001",
			6466 => "0000000110010100100001",
			6467 => "0001010111111100001000",
			6468 => "0000000111000000000100",
			6469 => "0000000110010100100001",
			6470 => "0000000110010100100001",
			6471 => "0000000110010100100001",
			6472 => "0000001010101101000000",
			6473 => "0011000111001000001100",
			6474 => "0001110110100100000100",
			6475 => "1111111110010110100101",
			6476 => "0001101101111100000100",
			6477 => "0000000110010110100101",
			6478 => "0000000110010110100101",
			6479 => "0010101000010100110000",
			6480 => "0011010011001000011100",
			6481 => "0000001111001000001100",
			6482 => "0011100111010100001000",
			6483 => "0001001011101100000100",
			6484 => "0000000110010110100101",
			6485 => "1111111110010110100101",
			6486 => "0000001110010110100101",
			6487 => "0011010101110000001000",
			6488 => "0011111011101100000100",
			6489 => "1111111110010110100101",
			6490 => "0000000110010110100101",
			6491 => "0011101100111000000100",
			6492 => "0000000110010110100101",
			6493 => "0000001110010110100101",
			6494 => "0001001101101100001000",
			6495 => "0001111111011100000100",
			6496 => "0000000110010110100101",
			6497 => "0000001110010110100101",
			6498 => "0001110101110100001000",
			6499 => "0010000001010100000100",
			6500 => "1111111110010110100101",
			6501 => "0000000110010110100101",
			6502 => "0000000110010110100101",
			6503 => "0000010110010110100101",
			6504 => "1111111110010110100101",
			6505 => "0011000100011000101100",
			6506 => "0000001011010100011100",
			6507 => "0011110110111100011000",
			6508 => "0011001010111000001000",
			6509 => "0001110110100100000100",
			6510 => "0000000110011010111001",
			6511 => "0000000110011010111001",
			6512 => "0001000111010100001100",
			6513 => "0000110110111100001000",
			6514 => "0001111011000000000100",
			6515 => "0000000110011010111001",
			6516 => "0000000110011010111001",
			6517 => "0000000110011010111001",
			6518 => "0000000110011010111001",
			6519 => "0000000110011010111001",
			6520 => "0001111000011000001100",
			6521 => "0001001011101100000100",
			6522 => "0000000110011010111001",
			6523 => "0010110110110100000100",
			6524 => "1111111110011010111001",
			6525 => "0000000110011010111001",
			6526 => "0000000110011010111001",
			6527 => "0011001011000000111100",
			6528 => "0011010100101000101100",
			6529 => "0001001000101000011100",
			6530 => "0001100100110100010000",
			6531 => "0001001100010000001000",
			6532 => "0001101101111100000100",
			6533 => "0000000110011010111001",
			6534 => "0000000110011010111001",
			6535 => "0011110010000100000100",
			6536 => "0000000110011010111001",
			6537 => "0000000110011010111001",
			6538 => "0000001111001000001000",
			6539 => "0000111100000000000100",
			6540 => "0000000110011010111001",
			6541 => "0000001110011010111001",
			6542 => "0000000110011010111001",
			6543 => "0000111000100000001000",
			6544 => "0010110001011000000100",
			6545 => "0000000110011010111001",
			6546 => "0000000110011010111001",
			6547 => "0000101101101100000100",
			6548 => "0000000110011010111001",
			6549 => "0000000110011010111001",
			6550 => "0000101100010000001000",
			6551 => "0010110010001000000100",
			6552 => "0000000110011010111001",
			6553 => "0000000110011010111001",
			6554 => "0001101011001100000100",
			6555 => "1111111110011010111001",
			6556 => "0000000110011010111001",
			6557 => "0000101110110100001000",
			6558 => "0011010100101000000100",
			6559 => "0000000110011010111001",
			6560 => "0000000110011010111001",
			6561 => "0011000110100100010000",
			6562 => "0000001010101100001100",
			6563 => "0001011101000100000100",
			6564 => "0000000110011010111001",
			6565 => "0011011100010100000100",
			6566 => "0000001110011010111001",
			6567 => "0000000110011010111001",
			6568 => "0000000110011010111001",
			6569 => "0010001100011100001000",
			6570 => "0010110101110100000100",
			6571 => "0000000110011010111001",
			6572 => "0000000110011010111001",
			6573 => "0000000110011010111001",
			6574 => "0010011111000000010000",
			6575 => "0010101001100100001100",
			6576 => "0000100001101000000100",
			6577 => "1111111110011110001101",
			6578 => "0001100101011100000100",
			6579 => "0000001110011110001101",
			6580 => "0000000110011110001101",
			6581 => "1111111110011110001101",
			6582 => "0011011100010101000100",
			6583 => "0001110110100100100100",
			6584 => "0000101100000000001100",
			6585 => "0001010010110100000100",
			6586 => "0000000110011110001101",
			6587 => "0001011100100100000100",
			6588 => "0000001110011110001101",
			6589 => "0000000110011110001101",
			6590 => "0011000100011000001100",
			6591 => "0010100010101100000100",
			6592 => "1111110110011110001101",
			6593 => "0010100011101000000100",
			6594 => "0000000110011110001101",
			6595 => "1111111110011110001101",
			6596 => "0011011111010000000100",
			6597 => "1111111110011110001101",
			6598 => "0001000110111000000100",
			6599 => "0000001110011110001101",
			6600 => "0000000110011110001101",
			6601 => "0010101001000100011100",
			6602 => "0011101100111000010000",
			6603 => "0010001000100100001000",
			6604 => "0001001100010000000100",
			6605 => "0000001110011110001101",
			6606 => "1111111110011110001101",
			6607 => "0000011101111100000100",
			6608 => "0000001110011110001101",
			6609 => "0000000110011110001101",
			6610 => "0011100011000000001000",
			6611 => "0001001000110100000100",
			6612 => "0000001110011110001101",
			6613 => "0000000110011110001101",
			6614 => "0000011110011110001101",
			6615 => "1111111110011110001101",
			6616 => "0010010100101100010100",
			6617 => "0011001001110100000100",
			6618 => "0000000110011110001101",
			6619 => "0001110101100100001000",
			6620 => "0010110001001000000100",
			6621 => "0000001110011110001101",
			6622 => "0000000110011110001101",
			6623 => "0011000100000100000100",
			6624 => "0000000110011110001101",
			6625 => "0000000110011110001101",
			6626 => "1111111110011110001101",
			6627 => "0011001010111000010000",
			6628 => "0000000110001000001100",
			6629 => "0011101100000000001000",
			6630 => "0001110110100100000100",
			6631 => "0000000110100010000001",
			6632 => "0000000110100010000001",
			6633 => "0000000110100010000001",
			6634 => "1111111110100010000001",
			6635 => "0010010100101101000100",
			6636 => "0000101100010000100100",
			6637 => "0011010101001000001000",
			6638 => "0000000001010100000100",
			6639 => "0000000110100010000001",
			6640 => "0000000110100010000001",
			6641 => "0000000101000100010000",
			6642 => "0000111100000000001000",
			6643 => "0010100111101100000100",
			6644 => "0000000110100010000001",
			6645 => "0000000110100010000001",
			6646 => "0000010000111100000100",
			6647 => "0000000110100010000001",
			6648 => "0000000110100010000001",
			6649 => "0010100000001000000100",
			6650 => "0000000110100010000001",
			6651 => "0000111010000100000100",
			6652 => "0000001110100010000001",
			6653 => "0000000110100010000001",
			6654 => "0011001001110100010000",
			6655 => "0011000100011000000100",
			6656 => "0000000110100010000001",
			6657 => "0010110101100100000100",
			6658 => "0000000110100010000001",
			6659 => "0011010010011100000100",
			6660 => "0000000110100010000001",
			6661 => "0000000110100010000001",
			6662 => "0010101010100100000100",
			6663 => "0000001110100010000001",
			6664 => "0000010000111100000100",
			6665 => "0000000110100010000001",
			6666 => "0000101101101100000100",
			6667 => "0000000110100010000001",
			6668 => "0000000110100010000001",
			6669 => "0001000001011100001100",
			6670 => "0000110110111100000100",
			6671 => "0000000110100010000001",
			6672 => "0000011101111100000100",
			6673 => "0000001110100010000001",
			6674 => "0000000110100010000001",
			6675 => "0000101000100000001000",
			6676 => "0010110101100100000100",
			6677 => "0000000110100010000001",
			6678 => "1111111110100010000001",
			6679 => "0000000001110100001000",
			6680 => "0000011100011000000100",
			6681 => "0000001110100010000001",
			6682 => "0000000110100010000001",
			6683 => "0011101100111000000100",
			6684 => "0000000110100010000001",
			6685 => "0011111011110000000100",
			6686 => "0000000110100010000001",
			6687 => "0000000110100010000001",
			6688 => "0010011001100100001100",
			6689 => "0010101001100100001000",
			6690 => "0001000111010000000100",
			6691 => "0000000110100101001101",
			6692 => "0000000110100101001101",
			6693 => "1111111110100101001101",
			6694 => "0001001100010000001100",
			6695 => "0000111100000000001000",
			6696 => "0010011111000000000100",
			6697 => "0000000110100101001101",
			6698 => "0000001110100101001101",
			6699 => "0000000110100101001101",
			6700 => "0001110110100100101000",
			6701 => "0000111010000100011100",
			6702 => "0001000111010100010000",
			6703 => "0000011011111100001000",
			6704 => "0010011000010000000100",
			6705 => "0000000110100101001101",
			6706 => "0000000110100101001101",
			6707 => "0001111001001000000100",
			6708 => "0000000110100101001101",
			6709 => "0000000110100101001101",
			6710 => "0001111001001000001000",
			6711 => "0001111001001000000100",
			6712 => "0000000110100101001101",
			6713 => "0000000110100101001101",
			6714 => "1111111110100101001101",
			6715 => "0001000011000000000100",
			6716 => "0000001110100101001101",
			6717 => "0010111011011100000100",
			6718 => "1111111110100101001101",
			6719 => "0000000110100101001101",
			6720 => "0010001000100100001100",
			6721 => "0011111100000000001000",
			6722 => "0010100000001000000100",
			6723 => "1111111110100101001101",
			6724 => "0000000110100101001101",
			6725 => "0000000110100101001101",
			6726 => "0000101100000000001100",
			6727 => "0010110101110100001000",
			6728 => "0000110010000100000100",
			6729 => "0000000110100101001101",
			6730 => "0000001110100101001101",
			6731 => "0000000110100101001101",
			6732 => "0011101100000000001000",
			6733 => "0010110100010000000100",
			6734 => "1111111110100101001101",
			6735 => "0000000110100101001101",
			6736 => "0000101000001100000100",
			6737 => "0000000110100101001101",
			6738 => "0000000110100101001101",
			6739 => "0011001010111000001000",
			6740 => "0000000110001000000100",
			6741 => "0000000110101000100001",
			6742 => "0000000110101000100001",
			6743 => "0011001000000000110100",
			6744 => "0010110101110100101100",
			6745 => "0001110110100100011000",
			6746 => "0001111001001000001100",
			6747 => "0000001111001000001000",
			6748 => "0001111011000000000100",
			6749 => "0000000110101000100001",
			6750 => "0000000110101000100001",
			6751 => "0000000110101000100001",
			6752 => "0000111000001100001000",
			6753 => "0001001000001100000100",
			6754 => "0000000110101000100001",
			6755 => "0000000110101000100001",
			6756 => "0000000110101000100001",
			6757 => "0000000010101000010000",
			6758 => "0000010000111100001000",
			6759 => "0001111000011000000100",
			6760 => "0000000110101000100001",
			6761 => "0000000110101000100001",
			6762 => "0010110000011100000100",
			6763 => "0000000110101000100001",
			6764 => "0000001110101000100001",
			6765 => "0000000110101000100001",
			6766 => "0010010101010000000100",
			6767 => "0000000110101000100001",
			6768 => "0000000110101000100001",
			6769 => "0010110100010000001100",
			6770 => "0001101000010000001000",
			6771 => "0011001001110100000100",
			6772 => "0000000110101000100001",
			6773 => "0000000110101000100001",
			6774 => "0000000110101000100001",
			6775 => "0011011100010100010000",
			6776 => "0001111000011000000100",
			6777 => "0000000110101000100001",
			6778 => "0011000001101000001000",
			6779 => "0000001000101100000100",
			6780 => "0000000110101000100001",
			6781 => "0000000110101000100001",
			6782 => "0000000110101000100001",
			6783 => "0001110000011100001000",
			6784 => "0010010010101100000100",
			6785 => "0000000110101000100001",
			6786 => "0000000110101000100001",
			6787 => "0000010111101000001000",
			6788 => "0010111110101100000100",
			6789 => "0000000110101000100001",
			6790 => "0000000110101000100001",
			6791 => "0000000110101000100001",
			6792 => "0000000010101001110000",
			6793 => "0011000100011000111100",
			6794 => "0000000110001000101000",
			6795 => "0010010100111100010000",
			6796 => "0011000100011000000100",
			6797 => "1111111110101100101101",
			6798 => "0011000100011000000100",
			6799 => "0000001110101100101101",
			6800 => "0011000100011000000100",
			6801 => "0000000110101100101101",
			6802 => "1111111110101100101101",
			6803 => "0011010101110000010000",
			6804 => "0011011110000100001000",
			6805 => "0000001100000100000100",
			6806 => "0000000110101100101101",
			6807 => "1111111110101100101101",
			6808 => "0000010111101000000100",
			6809 => "0000001110101100101101",
			6810 => "0000000110101100101101",
			6811 => "0001001000001100000100",
			6812 => "0000001110101100101101",
			6813 => "1111111110101100101101",
			6814 => "0001101001100100001100",
			6815 => "0010001100011100001000",
			6816 => "0011111010000100000100",
			6817 => "0000000110101100101101",
			6818 => "1111110110101100101101",
			6819 => "1111111110101100101101",
			6820 => "0000111011111000000100",
			6821 => "1111111110101100101101",
			6822 => "0000001110101100101101",
			6823 => "0001010101110000100100",
			6824 => "0000011001011000001000",
			6825 => "0010011111000000000100",
			6826 => "1111111110101100101101",
			6827 => "0000000110101100101101",
			6828 => "0011001000000000010000",
			6829 => "0000010000111100001000",
			6830 => "0000111010000100000100",
			6831 => "0000001110101100101101",
			6832 => "1111111110101100101101",
			6833 => "0001001000101000000100",
			6834 => "0000001110101100101101",
			6835 => "0000000110101100101101",
			6836 => "0011111110110100000100",
			6837 => "1111111110101100101101",
			6838 => "0001011001010000000100",
			6839 => "0000001110101100101101",
			6840 => "0000000110101100101101",
			6841 => "0001001101101100000100",
			6842 => "0000001110101100101101",
			6843 => "0011001000011000000100",
			6844 => "1111111110101100101101",
			6845 => "0000110010010100000100",
			6846 => "0000001110101100101101",
			6847 => "1111111110101100101101",
			6848 => "0000001010101100010100",
			6849 => "0000001010101100000100",
			6850 => "1111111110101100101101",
			6851 => "0000011010011000001100",
			6852 => "0010010010101100000100",
			6853 => "0000000110101100101101",
			6854 => "0000011100011000000100",
			6855 => "0000000110101100101101",
			6856 => "0000000110101100101101",
			6857 => "0000000110101100101101",
			6858 => "1111111110101100101101",
			6859 => "0000000010101001111100",
			6860 => "0011000100011000110100",
			6861 => "0000000110001000100100",
			6862 => "0010010100111100001100",
			6863 => "0001100000111100001000",
			6864 => "0011000110000100000100",
			6865 => "0000000110110001001001",
			6866 => "0000000110110001001001",
			6867 => "1111111110110001001001",
			6868 => "0011010101110000010000",
			6869 => "0011011110000100001000",
			6870 => "0000100010000000000100",
			6871 => "0000000110110001001001",
			6872 => "1111111110110001001001",
			6873 => "0010001010110000000100",
			6874 => "0000001110110001001001",
			6875 => "0000001110110001001001",
			6876 => "0001110001101000000100",
			6877 => "1111111110110001001001",
			6878 => "0000001110110001001001",
			6879 => "0010001100011100001000",
			6880 => "0011110111010100000100",
			6881 => "0000000110110001001001",
			6882 => "1111101110110001001001",
			6883 => "0010111011011100000100",
			6884 => "1111111110110001001001",
			6885 => "0000000110110001001001",
			6886 => "0001011111010000100100",
			6887 => "0001011111010000011100",
			6888 => "0010011111000000001100",
			6889 => "0000000001010100001000",
			6890 => "0010110010001000000100",
			6891 => "1111111110110001001001",
			6892 => "1111110110110001001001",
			6893 => "0000000110110001001001",
			6894 => "0011001011000000001000",
			6895 => "0000001111001000000100",
			6896 => "0000001110110001001001",
			6897 => "1111111110110001001001",
			6898 => "0001101101111100000100",
			6899 => "0000000110110001001001",
			6900 => "0000001110110001001001",
			6901 => "0000010000111100000100",
			6902 => "0000010110110001001001",
			6903 => "0000001110110001001001",
			6904 => "0001111000011000010000",
			6905 => "0000010000111100001000",
			6906 => "0010001000100100000100",
			6907 => "0000000110110001001001",
			6908 => "1111111110110001001001",
			6909 => "0000111011101100000100",
			6910 => "0000001110110001001001",
			6911 => "0000000110110001001001",
			6912 => "0000100110101100001000",
			6913 => "0010110100010000000100",
			6914 => "0000000110110001001001",
			6915 => "0000001110110001001001",
			6916 => "0000011110010100000100",
			6917 => "1111111110110001001001",
			6918 => "0000010100110100000100",
			6919 => "0000001110110001001001",
			6920 => "1111111110110001001001",
			6921 => "0000001010101100010000",
			6922 => "0000001010101100000100",
			6923 => "0000000110110001001001",
			6924 => "0000011010011000001000",
			6925 => "0000011100011000000100",
			6926 => "0000000110110001001001",
			6927 => "0000000110110001001001",
			6928 => "0000000110110001001001",
			6929 => "1111111110110001001001",
			6930 => "0011000111001000001000",
			6931 => "0001110110100100000100",
			6932 => "1111111110110011110101",
			6933 => "0000000110110011110101",
			6934 => "0001001000110101001100",
			6935 => "0010110110110100101100",
			6936 => "0000011101111100011100",
			6937 => "0011010101110000010000",
			6938 => "0000110111010100001000",
			6939 => "0000010111101000000100",
			6940 => "0000000110110011110101",
			6941 => "1111111110110011110101",
			6942 => "0000001111001000000100",
			6943 => "0000001110110011110101",
			6944 => "0000000110110011110101",
			6945 => "0010000001010000001000",
			6946 => "0011000100011000000100",
			6947 => "0000000110110011110101",
			6948 => "1111111110110011110101",
			6949 => "0000001110110011110101",
			6950 => "0000111111100100000100",
			6951 => "1111111110110011110101",
			6952 => "0000000111000100000100",
			6953 => "0000001110110011110101",
			6954 => "0011000100011000000100",
			6955 => "0000000110110011110101",
			6956 => "1111111110110011110101",
			6957 => "0000101110110100001000",
			6958 => "0011001011000000000100",
			6959 => "0000000110110011110101",
			6960 => "1111111110110011110101",
			6961 => "0000111010000100001000",
			6962 => "0011001011000000000100",
			6963 => "0000000110110011110101",
			6964 => "0000001110110011110101",
			6965 => "0000010101011100001000",
			6966 => "0011001011000000000100",
			6967 => "1111111110110011110101",
			6968 => "0000000110110011110101",
			6969 => "0011011100010100000100",
			6970 => "0000001110110011110101",
			6971 => "0000000110110011110101",
			6972 => "1111111110110011110101",
			6973 => "0000001010101101101100",
			6974 => "0001111000011001001000",
			6975 => "0001111000011000111000",
			6976 => "0001110110100100011000",
			6977 => "0001111001001000001100",
			6978 => "0001111011000000000100",
			6979 => "0000000110110111010001",
			6980 => "0011011001010000000100",
			6981 => "0000000110110111010001",
			6982 => "0000000110110111010001",
			6983 => "0000100110010000000100",
			6984 => "0000000110110111010001",
			6985 => "0010110000011100000100",
			6986 => "0000000110110111010001",
			6987 => "1111111110110111010001",
			6988 => "0001011101000100010000",
			6989 => "0010110000011100001000",
			6990 => "0010110100000100000100",
			6991 => "0000000110110111010001",
			6992 => "0000001110110111010001",
			6993 => "0000011011111100000100",
			6994 => "0000000110110111010001",
			6995 => "1111111110110111010001",
			6996 => "0000011101111100001000",
			6997 => "0010001000010100000100",
			6998 => "0000000110110111010001",
			6999 => "0000000110110111010001",
			7000 => "0010111011011100000100",
			7001 => "1111111110110111010001",
			7002 => "0000000110110111010001",
			7003 => "0001100100110100000100",
			7004 => "0000000110110111010001",
			7005 => "0011010101110000000100",
			7006 => "0000000110110111010001",
			7007 => "0001101011001100000100",
			7008 => "1111111110110111010001",
			7009 => "0000000110110111010001",
			7010 => "0011011010001000001000",
			7011 => "0010001000100100000100",
			7012 => "0000000110110111010001",
			7013 => "0000001110110111010001",
			7014 => "0010110101110100001000",
			7015 => "0001011001010000000100",
			7016 => "0000000110110111010001",
			7017 => "1111111110110111010001",
			7018 => "0011011100010100001000",
			7019 => "0011011110010000000100",
			7020 => "0000000110110111010001",
			7021 => "0000001110110111010001",
			7022 => "0001110101110100001000",
			7023 => "0001101000010000000100",
			7024 => "0000000110110111010001",
			7025 => "0000000110110111010001",
			7026 => "0000000110110111010001",
			7027 => "1111111110110111010001",
			7028 => "0011000111001000001000",
			7029 => "0001110110100100000100",
			7030 => "1111111110111011010101",
			7031 => "0000000110111011010101",
			7032 => "0000101000001101001000",
			7033 => "0010101010100000100000",
			7034 => "0001011110101000001000",
			7035 => "0011001010111000000100",
			7036 => "0000000110111011010101",
			7037 => "0000000110111011010101",
			7038 => "0000100010000100001100",
			7039 => "0010001000100100001000",
			7040 => "0000100110010000000100",
			7041 => "0000000110111011010101",
			7042 => "1111111110111011010101",
			7043 => "0000000110111011010101",
			7044 => "0000101100000000001000",
			7045 => "0000011001011000000100",
			7046 => "0000000110111011010101",
			7047 => "0000000110111011010101",
			7048 => "0000000110111011010101",
			7049 => "0001011101000100011000",
			7050 => "0001010010110100001100",
			7051 => "0001110110100100000100",
			7052 => "0000000110111011010101",
			7053 => "0000000110001000000100",
			7054 => "0000000110111011010101",
			7055 => "0000000110111011010101",
			7056 => "0010010100101100001000",
			7057 => "0010110101100100000100",
			7058 => "0000000110111011010101",
			7059 => "0000000110111011010101",
			7060 => "0000000110111011010101",
			7061 => "0000111011111000001000",
			7062 => "0000010000111100000100",
			7063 => "0000000110111011010101",
			7064 => "0000001110111011010101",
			7065 => "0000101010000100000100",
			7066 => "0000000110111011010101",
			7067 => "0000000110111011010101",
			7068 => "0011100111010100010000",
			7069 => "0001101101011000000100",
			7070 => "0000000110111011010101",
			7071 => "0001111001001000000100",
			7072 => "0000000110111011010101",
			7073 => "0011111000001100000100",
			7074 => "0000000110111011010101",
			7075 => "1111111110111011010101",
			7076 => "0000101011111000000100",
			7077 => "0000000110111011010101",
			7078 => "0011101100111000010000",
			7079 => "0010111010010100001000",
			7080 => "0001110001101000000100",
			7081 => "0000000110111011010101",
			7082 => "0000000110111011010101",
			7083 => "0000100001011100000100",
			7084 => "0000000110111011010101",
			7085 => "0000000110111011010101",
			7086 => "0001101000010000001000",
			7087 => "0000000001110100000100",
			7088 => "0000000110111011010101",
			7089 => "0000000110111011010101",
			7090 => "0000001010101100000100",
			7091 => "0000001110111011010101",
			7092 => "0000000110111011010101",
			7093 => "0000001010101101111100",
			7094 => "0010110110110101000000",
			7095 => "0001001100010000010100",
			7096 => "0010011111000000001100",
			7097 => "0010000100101100001000",
			7098 => "0010111110110000000100",
			7099 => "0000000110111111010001",
			7100 => "0000001110111111010001",
			7101 => "1111111110111111010001",
			7102 => "0001011100100100000100",
			7103 => "0000001110111111010001",
			7104 => "0000000110111111010001",
			7105 => "0011100111010100011100",
			7106 => "0000101000001100010000",
			7107 => "0011100111011000001000",
			7108 => "0000001001101000000100",
			7109 => "0000000110111111010001",
			7110 => "1111111110111111010001",
			7111 => "0011000100011000000100",
			7112 => "0000000110111111010001",
			7113 => "0000001110111111010001",
			7114 => "0001110001101000001000",
			7115 => "0011001010111000000100",
			7116 => "0000000110111111010001",
			7117 => "1111111110111111010001",
			7118 => "1111110110111111010001",
			7119 => "0000000111000100001000",
			7120 => "0010010111101100000100",
			7121 => "0000000110111111010001",
			7122 => "0000001110111111010001",
			7123 => "0000101000101000000100",
			7124 => "1111111110111111010001",
			7125 => "0000000110111111010001",
			7126 => "0001011111010000011100",
			7127 => "0010001000100100000100",
			7128 => "1111111110111111010001",
			7129 => "0010110101110100010000",
			7130 => "0011001011000000001000",
			7131 => "0011000100011000000100",
			7132 => "0000000110111111010001",
			7133 => "0000000110111111010001",
			7134 => "0011001001110100000100",
			7135 => "0000001110111111010001",
			7136 => "0000000110111111010001",
			7137 => "0011110110111100000100",
			7138 => "0000000110111111010001",
			7139 => "0000000110111111010001",
			7140 => "0010000001010100011000",
			7141 => "0011001001110100001100",
			7142 => "0001010010011100001000",
			7143 => "0010010100111100000100",
			7144 => "0000000110111111010001",
			7145 => "0000001110111111010001",
			7146 => "1111111110111111010001",
			7147 => "0000000111000100001000",
			7148 => "0011110110111100000100",
			7149 => "0000000110111111010001",
			7150 => "0000001110111111010001",
			7151 => "1111111110111111010001",
			7152 => "0010111010010100000100",
			7153 => "0000001110111111010001",
			7154 => "0000000110111111010001",
			7155 => "1111111110111111010001",
			7156 => "0000001010101101111000",
			7157 => "0001110110100100100100",
			7158 => "0001001010000100001100",
			7159 => "0000010000111100001000",
			7160 => "0001100000111100000100",
			7161 => "0000000111000011000101",
			7162 => "0000000111000011000101",
			7163 => "0000000111000011000101",
			7164 => "0001101011001100001000",
			7165 => "0010101010100000000100",
			7166 => "0000000111000011000101",
			7167 => "1111111111000011000101",
			7168 => "0010101000100100001100",
			7169 => "0010110000011100000100",
			7170 => "0000000111000011000101",
			7171 => "0011100111011000000100",
			7172 => "0000000111000011000101",
			7173 => "0000000111000011000101",
			7174 => "1111111111000011000101",
			7175 => "0001110001101000011100",
			7176 => "0011100111010100010100",
			7177 => "0011110000010000010000",
			7178 => "0010000111110100001000",
			7179 => "0001010010110100000100",
			7180 => "0000000111000011000101",
			7181 => "0000000111000011000101",
			7182 => "0010110000011100000100",
			7183 => "0000000111000011000101",
			7184 => "0000001111000011000101",
			7185 => "0000000111000011000101",
			7186 => "0010101000100100000100",
			7187 => "0000001111000011000101",
			7188 => "0000000111000011000101",
			7189 => "0011111111010100100000",
			7190 => "0001111000011000010000",
			7191 => "0001101101111100001000",
			7192 => "0001011110101000000100",
			7193 => "0000000111000011000101",
			7194 => "0000000111000011000101",
			7195 => "0011010101001000000100",
			7196 => "0000000111000011000101",
			7197 => "0000001111000011000101",
			7198 => "0000000001010100001000",
			7199 => "0000110110111100000100",
			7200 => "0000001111000011000101",
			7201 => "1111111111000011000101",
			7202 => "0011100010000100000100",
			7203 => "0000000111000011000101",
			7204 => "0000001111000011000101",
			7205 => "0011101011111000001100",
			7206 => "0000000110001000001000",
			7207 => "0001101101011000000100",
			7208 => "1111111111000011000101",
			7209 => "0000001111000011000101",
			7210 => "1111111111000011000101",
			7211 => "0010000001010100001000",
			7212 => "0000010100110100000100",
			7213 => "0000000111000011000101",
			7214 => "1111111111000011000101",
			7215 => "0000001111000011000101",
			7216 => "1111111111000011000101",
			7217 => "0000001010101110000000",
			7218 => "0000010000111100111100",
			7219 => "0000111010000100101100",
			7220 => "0000101110110100011100",
			7221 => "0001001100010000001100",
			7222 => "0001101101111100001000",
			7223 => "0001100000111100000100",
			7224 => "0000000111000111001011",
			7225 => "0000000111000111001011",
			7226 => "0000001111000111001011",
			7227 => "0001100100110100001000",
			7228 => "0010001000100100000100",
			7229 => "1111111111000111001011",
			7230 => "0000000111000111001011",
			7231 => "0000111100010000000100",
			7232 => "0000000111000111001011",
			7233 => "0000000111000111001011",
			7234 => "0010110010001000001100",
			7235 => "0001100100110100000100",
			7236 => "1111111111000111001011",
			7237 => "0000011001011000000100",
			7238 => "0000000111000111001011",
			7239 => "0000001111000111001011",
			7240 => "0000001111000111001011",
			7241 => "0010011111000000000100",
			7242 => "1111111111000111001011",
			7243 => "0000110111010100000100",
			7244 => "0000000111000111001011",
			7245 => "0010110100010000000100",
			7246 => "1111111111000111001011",
			7247 => "0000000111000111001011",
			7248 => "0001110001101000100000",
			7249 => "0000010101011100000100",
			7250 => "0000001111000111001011",
			7251 => "0010011001111100001100",
			7252 => "0000100111011000001000",
			7253 => "0010101010100000000100",
			7254 => "1111111111000111001011",
			7255 => "0000001111000111001011",
			7256 => "1111111111000111001011",
			7257 => "0011101100010000001000",
			7258 => "0001000111010100000100",
			7259 => "0000000111000111001011",
			7260 => "1111111111000111001011",
			7261 => "0001000001011100000100",
			7262 => "0000001111000111001011",
			7263 => "0000000111000111001011",
			7264 => "0001010111111100011000",
			7265 => "0010010100111100001000",
			7266 => "0001000111010100000100",
			7267 => "0000000111000111001011",
			7268 => "0000000111000111001011",
			7269 => "0010111011011100001000",
			7270 => "0001000001011100000100",
			7271 => "0000000111000111001011",
			7272 => "0000000111000111001011",
			7273 => "0001110111010000000100",
			7274 => "0000001111000111001011",
			7275 => "0000000111000111001011",
			7276 => "0001110101110100001000",
			7277 => "0001011110010000000100",
			7278 => "0000000111000111001011",
			7279 => "1111111111000111001011",
			7280 => "0000000111000111001011",
			7281 => "1111111111000111001011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2358, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4838, initial_addr_3'length));
	end generate gen_rom_2;

	gen_rom_3: if SELECT_ROM = 3 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000010101100000100",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0011001100110000000100",
			26 => "0000000000000001110001",
			27 => "0000000000000001110001",
			28 => "0000101000000000000100",
			29 => "0000000000000001111101",
			30 => "0000000000000001111101",
			31 => "0001000111001000000100",
			32 => "0000000000000010001001",
			33 => "0000000000000010001001",
			34 => "0011111011000000000100",
			35 => "0000000000000010010101",
			36 => "0000000000000010010101",
			37 => "0001000110110100000100",
			38 => "0000000000000010100001",
			39 => "0000000000000010100001",
			40 => "0000101000000000000100",
			41 => "0000000000000010101101",
			42 => "0000000000000010101101",
			43 => "0001000111010000000100",
			44 => "0000000000000011000001",
			45 => "0010011110010100000100",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0010010000111100000100",
			49 => "0000000000000011010101",
			50 => "0010011001100100000100",
			51 => "0000000000000011010101",
			52 => "0000000000000011010101",
			53 => "0000000010101100000100",
			54 => "0000000000000011101001",
			55 => "0011111100010100000100",
			56 => "0000000000000011101001",
			57 => "0000000000000011101001",
			58 => "0011111001001000001000",
			59 => "0000000101000100000100",
			60 => "0000000000000011111101",
			61 => "0000000000000011111101",
			62 => "0000000000000011111101",
			63 => "0000000110011000001000",
			64 => "0011100010001000000100",
			65 => "0000001000000100010001",
			66 => "1101011000000100010001",
			67 => "1100010000000100010001",
			68 => "0010101101011000001000",
			69 => "0011000110000100000100",
			70 => "0000001000000100101101",
			71 => "0000000000000100101101",
			72 => "0010010101011100000100",
			73 => "0000000000000100101101",
			74 => "0000000000000100101101",
			75 => "0000101000000000001000",
			76 => "0001101101011100000100",
			77 => "0000000000000101001001",
			78 => "0000000000000101001001",
			79 => "0000010111100100000100",
			80 => "0000000000000101001001",
			81 => "0000000000000101001001",
			82 => "0000101000000000001000",
			83 => "0011000100000000000100",
			84 => "0000000000000101100101",
			85 => "0000000000000101100101",
			86 => "0001110111010000000100",
			87 => "0000000000000101100101",
			88 => "0000000000000101100101",
			89 => "0010010101011100001100",
			90 => "0000100100001000000100",
			91 => "0000000000000110000001",
			92 => "0000010110101000000100",
			93 => "0000000000000110000001",
			94 => "0000000000000110000001",
			95 => "0000000000000110000001",
			96 => "0000010110101000000100",
			97 => "0000000000000110011101",
			98 => "0011100111110000001000",
			99 => "0010000111110100000100",
			100 => "0000000000000110011101",
			101 => "0000000000000110011101",
			102 => "0000000000000110011101",
			103 => "0010010000111100001100",
			104 => "0011100100001000000100",
			105 => "0000000000000110111001",
			106 => "0000010110101000000100",
			107 => "0000000000000110111001",
			108 => "0000000000000110111001",
			109 => "0000000000000110111001",
			110 => "0001000111010000000100",
			111 => "0000000000000111010101",
			112 => "0000000010101100000100",
			113 => "0000000000000111010101",
			114 => "0011111010011100000100",
			115 => "0000000000000111010101",
			116 => "0000000000000111010101",
			117 => "0000000010101100001000",
			118 => "0011000110000100000100",
			119 => "0000000000000111111001",
			120 => "0000000000000111111001",
			121 => "0000010111100100001000",
			122 => "0011001110001100000100",
			123 => "0000000000000111111001",
			124 => "0000000000000111111001",
			125 => "0000000000000111111001",
			126 => "0000100000110100010000",
			127 => "0010010000111100001000",
			128 => "0011100100001000000100",
			129 => "0000000000001000011101",
			130 => "0000000000001000011101",
			131 => "0011111011011100000100",
			132 => "0000000000001000011101",
			133 => "0000000000001000011101",
			134 => "0000000000001000011101",
			135 => "0011000100000000001100",
			136 => "0001000111001000000100",
			137 => "0000000000001001001001",
			138 => "0001111101100000000100",
			139 => "0000000000001001001001",
			140 => "0000000000001001001001",
			141 => "0010110100001000001000",
			142 => "0000000101000100000100",
			143 => "0000000000001001001001",
			144 => "0000000000001001001001",
			145 => "0000000000001001001001",
			146 => "0010010000111100000100",
			147 => "0000000000001001101101",
			148 => "0010011001100100001100",
			149 => "0001110101101100000100",
			150 => "0000000000001001101101",
			151 => "0000111001100000000100",
			152 => "0000000000001001101101",
			153 => "0000000000001001101101",
			154 => "0000000000001001101101",
			155 => "0010010000111100000100",
			156 => "0000000000001010010001",
			157 => "0010011001100100001100",
			158 => "0011010010011100001000",
			159 => "0011010110100100000100",
			160 => "0000000000001010010001",
			161 => "0000000000001010010001",
			162 => "0000000000001010010001",
			163 => "0000000000001010010001",
			164 => "0001000110110100010000",
			165 => "0010010101011100001100",
			166 => "0000111010111100000100",
			167 => "0000000000001010111101",
			168 => "0001111101100000000100",
			169 => "0000000000001010111101",
			170 => "0000000000001010111101",
			171 => "0000000000001010111101",
			172 => "0010010111101000000100",
			173 => "0000000000001010111101",
			174 => "0000000000001010111101",
			175 => "0000010110101000010000",
			176 => "0011110001111100000100",
			177 => "0000000000001011101001",
			178 => "0010110000001100001000",
			179 => "0001110110000100000100",
			180 => "0000000000001011101001",
			181 => "0000000000001011101001",
			182 => "0000000000001011101001",
			183 => "0011111011011100000100",
			184 => "0000001000001011101001",
			185 => "0000000000001011101001",
			186 => "0000101000000000001000",
			187 => "0000010110101000000100",
			188 => "0000000000001100010101",
			189 => "0000000000001100010101",
			190 => "0010010111101000001100",
			191 => "0000011101101000001000",
			192 => "0001000001101000000100",
			193 => "0000000000001100010101",
			194 => "0000000000001100010101",
			195 => "0000000000001100010101",
			196 => "0000000000001100010101",
			197 => "0011001100110000001000",
			198 => "0010010101011100000100",
			199 => "0000000000001101000001",
			200 => "0000000000001101000001",
			201 => "0010011001100100001100",
			202 => "0011001000000000001000",
			203 => "0010011101011100000100",
			204 => "0000000000001101000001",
			205 => "0000000000001101000001",
			206 => "0000000000001101000001",
			207 => "0000000000001101000001",
			208 => "0000100000110100010100",
			209 => "0010010000111100001100",
			210 => "0011100100001000000100",
			211 => "0000000000001101101101",
			212 => "0001111101100000000100",
			213 => "0000000000001101101101",
			214 => "0000000000001101101101",
			215 => "0011111011011100000100",
			216 => "0000000000001101101101",
			217 => "0000000000001101101101",
			218 => "0000000000001101101101",
			219 => "0010010101011100001100",
			220 => "0011100100001000000100",
			221 => "0000000000001110100001",
			222 => "0000010111100100000100",
			223 => "0000000000001110100001",
			224 => "0000000000001110100001",
			225 => "0000011001011000001100",
			226 => "0011101010001000001000",
			227 => "0001111101100000000100",
			228 => "0000000000001110100001",
			229 => "0000000000001110100001",
			230 => "0000000000001110100001",
			231 => "0000000000001110100001",
			232 => "0001000110110100010100",
			233 => "0000010110101000001100",
			234 => "0000111010111100000100",
			235 => "0000000000001111011101",
			236 => "0001111101100000000100",
			237 => "0000000000001111011101",
			238 => "0000000000001111011101",
			239 => "0001101001011000000100",
			240 => "0000000000001111011101",
			241 => "0000000000001111011101",
			242 => "0001111100101000001000",
			243 => "0011001110001100000100",
			244 => "0000000000001111011101",
			245 => "0000000000001111011101",
			246 => "0000000000001111011101",
			247 => "0010010000111100010000",
			248 => "0001000111001000000100",
			249 => "0000000000010000011001",
			250 => "0000010110101000001000",
			251 => "0001111110001100000100",
			252 => "0000000000010000011001",
			253 => "0000000000010000011001",
			254 => "0000000000010000011001",
			255 => "0010100111101100001100",
			256 => "0011101010001000001000",
			257 => "0000010111100100000100",
			258 => "0000000000010000011001",
			259 => "0000000000010000011001",
			260 => "0000000000010000011001",
			261 => "0000000000010000011001",
			262 => "0010000111110100011000",
			263 => "0010010000111100001100",
			264 => "0011111011000000001000",
			265 => "0001111001110000000100",
			266 => "0000000000010001001101",
			267 => "0000000000010001001101",
			268 => "0000000000010001001101",
			269 => "0001110110000100000100",
			270 => "0000000000010001001101",
			271 => "0000111001100000000100",
			272 => "0000000000010001001101",
			273 => "0000000000010001001101",
			274 => "0000000000010001001101",
			275 => "0010110101101100001000",
			276 => "0001000111001000000100",
			277 => "0000000000010010000001",
			278 => "0000000000010010000001",
			279 => "0001001001100000010000",
			280 => "0010010000111100000100",
			281 => "0000000000010010000001",
			282 => "0011101010001000001000",
			283 => "0000011001011000000100",
			284 => "0000000000010010000001",
			285 => "0000000000010010000001",
			286 => "0000000000010010000001",
			287 => "0000000000010010000001",
			288 => "0010010000111100001000",
			289 => "0011000110000100000100",
			290 => "0000000000010010110101",
			291 => "0000000000010010110101",
			292 => "0010011001100100010000",
			293 => "0001011110101000001100",
			294 => "0001111101100000000100",
			295 => "0000000000010010110101",
			296 => "0011001000000000000100",
			297 => "0000000000010010110101",
			298 => "0000000000010010110101",
			299 => "0000000000010010110101",
			300 => "0000000000010010110101",
			301 => "0000000010101100000100",
			302 => "0000000000010011100001",
			303 => "0000010111100100000100",
			304 => "0000000000010011100001",
			305 => "0000101110010000001100",
			306 => "0001101101111100001000",
			307 => "0001011101000100000100",
			308 => "0000000000010011100001",
			309 => "0000000000010011100001",
			310 => "0000000000010011100001",
			311 => "0000000000010011100001",
			312 => "0000000110011000010100",
			313 => "0011000100000000000100",
			314 => "0000000000010100011101",
			315 => "0011110001001000001100",
			316 => "0000010111100100001000",
			317 => "0000110110100100000100",
			318 => "0000001000010100011101",
			319 => "1111111000010100011101",
			320 => "0000001000010100011101",
			321 => "0000000000010100011101",
			322 => "0001001100010100001000",
			323 => "0010100100101100000100",
			324 => "1111111000010100011101",
			325 => "0000010000010100011101",
			326 => "1111111000010100011101",
			327 => "0011001100110000001100",
			328 => "0010100100110100000100",
			329 => "0000000000010101011001",
			330 => "0000010111100100000100",
			331 => "0000000000010101011001",
			332 => "0000000000010101011001",
			333 => "0000010110101000000100",
			334 => "0000000000010101011001",
			335 => "0000101110010000001100",
			336 => "0000011001011000001000",
			337 => "0000111001100000000100",
			338 => "0000000000010101011001",
			339 => "0000000000010101011001",
			340 => "0000000000010101011001",
			341 => "0000000000010101011001",
			342 => "0000000110011000011000",
			343 => "0011111011000000001000",
			344 => "0010110101101100000100",
			345 => "0000000000010110001101",
			346 => "0000001000010110001101",
			347 => "0010010101011100000100",
			348 => "1111111000010110001101",
			349 => "0011110010001000000100",
			350 => "0000001000010110001101",
			351 => "0010011101111100000100",
			352 => "1111111000010110001101",
			353 => "0000001000010110001101",
			354 => "1111111000010110001101",
			355 => "0010101001111100011000",
			356 => "0000110001001000010100",
			357 => "0011000100000000001000",
			358 => "0001000111001000000100",
			359 => "0000001000010111010001",
			360 => "0000000000010111010001",
			361 => "0011110010001000001000",
			362 => "0000100001101000000100",
			363 => "0000001000010111010001",
			364 => "0000001000010111010001",
			365 => "0000000000010111010001",
			366 => "0000011000010111010001",
			367 => "0001001100010100001000",
			368 => "0001001110010000000100",
			369 => "1111111000010111010001",
			370 => "0000000000010111010001",
			371 => "1111111000010111010001",
			372 => "0011001100110000010000",
			373 => "0000100100001000000100",
			374 => "0000000000011000010101",
			375 => "0010010101011100001000",
			376 => "0011011111011100000100",
			377 => "0000000000011000010101",
			378 => "0000000000011000010101",
			379 => "0000000000011000010101",
			380 => "0010010000111100000100",
			381 => "0000000000011000010101",
			382 => "0000101110010000001100",
			383 => "0010011001100100001000",
			384 => "0001011110101000000100",
			385 => "0000000000011000010101",
			386 => "0000000000011000010101",
			387 => "0000000000011000010101",
			388 => "0000000000011000010101",
			389 => "0000000110011000011000",
			390 => "0000011001111000000100",
			391 => "0000000000011001100001",
			392 => "0011110010001000001100",
			393 => "0011001000111000001000",
			394 => "0000110011100000000100",
			395 => "0000001000011001100001",
			396 => "0000000000011001100001",
			397 => "0000001000011001100001",
			398 => "0001110100001000000100",
			399 => "1111111000011001100001",
			400 => "0000001000011001100001",
			401 => "0001001001100000001100",
			402 => "0010100111101100000100",
			403 => "1111111000011001100001",
			404 => "0010000111110100000100",
			405 => "0000010000011001100001",
			406 => "0000000000011001100001",
			407 => "1111111000011001100001",
			408 => "0000010111100100011000",
			409 => "0011111011000000001100",
			410 => "0011000100000000000100",
			411 => "0000000000011010110101",
			412 => "0001100111101000000100",
			413 => "0000000000011010110101",
			414 => "0000000000011010110101",
			415 => "0011001110001100001000",
			416 => "0001101001011000000100",
			417 => "0000000000011010110101",
			418 => "0000000000011010110101",
			419 => "0000000000011010110101",
			420 => "0000101110010000010000",
			421 => "0001100000111100000100",
			422 => "0000000000011010110101",
			423 => "0000011001011000001000",
			424 => "0001011110101000000100",
			425 => "0000000000011010110101",
			426 => "0000000000011010110101",
			427 => "0000000000011010110101",
			428 => "0000000000011010110101",
			429 => "0001001100010100100000",
			430 => "0000010111100100010000",
			431 => "0001001001001000001000",
			432 => "0001101111001100000100",
			433 => "0000000000011011111001",
			434 => "0000001000011011111001",
			435 => "0000010110101000000100",
			436 => "1111111000011011111001",
			437 => "0000000000011011111001",
			438 => "0011110010001000000100",
			439 => "0000001000011011111001",
			440 => "0011010101110100000100",
			441 => "0000000000011011111001",
			442 => "0011111010001000000100",
			443 => "0000000000011011111001",
			444 => "0000000000011011111001",
			445 => "1111111000011011111001",
			446 => "0010110101101100001000",
			447 => "0001000111001000000100",
			448 => "0000000000011100111101",
			449 => "0000000000011100111101",
			450 => "0001000111010000000100",
			451 => "0000000000011100111101",
			452 => "0011001000000000001100",
			453 => "0011001000111100000100",
			454 => "0000000000011100111101",
			455 => "0011000110000100000100",
			456 => "0000000000011100111101",
			457 => "0000000000011100111101",
			458 => "0011001000000000001000",
			459 => "0010110101100100000100",
			460 => "0000000000011100111101",
			461 => "0000000000011100111101",
			462 => "0000000000011100111101",
			463 => "0010110101101100001000",
			464 => "0001000111001000000100",
			465 => "0000000000011110001001",
			466 => "0000000000011110001001",
			467 => "0011111010011100001000",
			468 => "0000001100000100000100",
			469 => "0000000000011110001001",
			470 => "0000000000011110001001",
			471 => "0000010111100100001000",
			472 => "0011001110001100000100",
			473 => "0000000000011110001001",
			474 => "0000000000011110001001",
			475 => "0010000111110100001100",
			476 => "0011101010001000001000",
			477 => "0010000100101100000100",
			478 => "0000000000011110001001",
			479 => "0000000000011110001001",
			480 => "0000000000011110001001",
			481 => "0000000000011110001001",
			482 => "0010000111110100100100",
			483 => "0000010111100100010100",
			484 => "0010000101010000001100",
			485 => "0011100100001000000100",
			486 => "0000000000011111010101",
			487 => "0001111101100000000100",
			488 => "0000000000011111010101",
			489 => "0000000000011111010101",
			490 => "0011000011011100000100",
			491 => "0000000000011111010101",
			492 => "0000000000011111010101",
			493 => "0011101010001000001100",
			494 => "0001011110101000001000",
			495 => "0000101110010000000100",
			496 => "0000000000011111010101",
			497 => "0000000000011111010101",
			498 => "0000000000011111010101",
			499 => "0000000000011111010101",
			500 => "1111111000011111010101",
			501 => "0001001100010100011100",
			502 => "0000010010001100000100",
			503 => "1111111000100000010001",
			504 => "0011111011000000000100",
			505 => "0000001000100000010001",
			506 => "0001110110000100001100",
			507 => "0000010111100100000100",
			508 => "1111111000100000010001",
			509 => "0011000011011100000100",
			510 => "0000000000100000010001",
			511 => "0000000000100000010001",
			512 => "0011111010001000000100",
			513 => "0000001000100000010001",
			514 => "0000000000100000010001",
			515 => "1111111000100000010001",
			516 => "0010000111110100100100",
			517 => "0000010111100100010000",
			518 => "0000000010101100001100",
			519 => "0000011001111000000100",
			520 => "0000000000100001011101",
			521 => "0000010110101000000100",
			522 => "0000000000100001011101",
			523 => "0000000000100001011101",
			524 => "0000000000100001011101",
			525 => "0011110010001000000100",
			526 => "0000000000100001011101",
			527 => "0011001000000000000100",
			528 => "0000000000100001011101",
			529 => "0000001100011100000100",
			530 => "0000000000100001011101",
			531 => "0000101100010100000100",
			532 => "0000000000100001011101",
			533 => "0000000000100001011101",
			534 => "1111111000100001011101",
			535 => "0010000111110100101000",
			536 => "0000010111100100010100",
			537 => "0011100100001000001000",
			538 => "0001101001011000000100",
			539 => "0000000000100010110001",
			540 => "0000000000100010110001",
			541 => "0000010110101000000100",
			542 => "0000000000100010110001",
			543 => "0001100000111100000100",
			544 => "0000000000100010110001",
			545 => "0000000000100010110001",
			546 => "0011101010001000010000",
			547 => "0001100000111100000100",
			548 => "0000000000100010110001",
			549 => "0011001100110000000100",
			550 => "0000000000100010110001",
			551 => "0001011101000100000100",
			552 => "0000000000100010110001",
			553 => "0000000000100010110001",
			554 => "0000000000100010110001",
			555 => "0000000000100010110001",
			556 => "0000000110011100011100",
			557 => "0011000100000000000100",
			558 => "0000000000100011101101",
			559 => "0001000111010000000100",
			560 => "0000001000100011101101",
			561 => "0011001100110000000100",
			562 => "0000000000100011101101",
			563 => "0011101010001000001100",
			564 => "0010010111101000000100",
			565 => "0000000000100011101101",
			566 => "0000111001100000000100",
			567 => "0000000000100011101101",
			568 => "0000000000100011101101",
			569 => "0000000000100011101101",
			570 => "1111111000100011101101",
			571 => "0000000110011100100100",
			572 => "0001110001101000011100",
			573 => "0000100000110100011000",
			574 => "0010010000111100001100",
			575 => "0001001001001000001000",
			576 => "0011000100000000000100",
			577 => "0000000000100100111001",
			578 => "0000001000100100111001",
			579 => "1111111000100100111001",
			580 => "0011110010001000000100",
			581 => "0000001000100100111001",
			582 => "0001011011011100000100",
			583 => "0000000000100100111001",
			584 => "0000001000100100111001",
			585 => "1111111000100100111001",
			586 => "0000101110010000000100",
			587 => "0000010000100100111001",
			588 => "0000000000100100111001",
			589 => "1111111000100100111001",
			590 => "0001001100010100100000",
			591 => "0000010010001100000100",
			592 => "1111111000100101111101",
			593 => "0000100001001000010100",
			594 => "0000010110101000010000",
			595 => "0011110111001000001100",
			596 => "0011100100001000000100",
			597 => "0000001000100101111101",
			598 => "0011100001111100000100",
			599 => "0000000000100101111101",
			600 => "0000001000100101111101",
			601 => "1111111000100101111101",
			602 => "0000001000100101111101",
			603 => "0010011101011000000100",
			604 => "1111111000100101111101",
			605 => "0000010000100101111101",
			606 => "1111111000100101111101",
			607 => "0000000110011100101000",
			608 => "0011001000000000011100",
			609 => "0000100000110100011000",
			610 => "0010010000111100001100",
			611 => "0001001001001000001000",
			612 => "0011000100000000000100",
			613 => "0000000000100111010001",
			614 => "0000001000100111010001",
			615 => "1111111000100111010001",
			616 => "0011100101100100000100",
			617 => "0000001000100111010001",
			618 => "0001110001111100000100",
			619 => "1111111000100111010001",
			620 => "0000001000100111010001",
			621 => "1111111000100111010001",
			622 => "0010110101100100000100",
			623 => "0000000000100111010001",
			624 => "0001011110101000000100",
			625 => "0000001000100111010001",
			626 => "0000000000100111010001",
			627 => "1111111000100111010001",
			628 => "0000000110011100100100",
			629 => "0001110001101000011100",
			630 => "0011110000110100011000",
			631 => "0011000100000000001000",
			632 => "0001000111001000000100",
			633 => "0000000000101000011101",
			634 => "1111111000101000011101",
			635 => "0011000011011100000100",
			636 => "0000001000101000011101",
			637 => "0000010111100100001000",
			638 => "0000110110100100000100",
			639 => "0000000000101000011101",
			640 => "0000000000101000011101",
			641 => "0000001000101000011101",
			642 => "0000000000101000011101",
			643 => "0000111001100000000100",
			644 => "0000001000101000011101",
			645 => "0000000000101000011101",
			646 => "1111111000101000011101",
			647 => "0010000111110100100100",
			648 => "0000011001111000001000",
			649 => "0011110000001100000100",
			650 => "0000000000101001101001",
			651 => "0000000000101001101001",
			652 => "0010110100001000000100",
			653 => "0000001000101001101001",
			654 => "0011001100110000001000",
			655 => "0011111010011100000100",
			656 => "0000000000101001101001",
			657 => "1111111000101001101001",
			658 => "0011101010001000001100",
			659 => "0000010111100100000100",
			660 => "0000000000101001101001",
			661 => "0001100000111100000100",
			662 => "0000000000101001101001",
			663 => "0000000000101001101001",
			664 => "0000000000101001101001",
			665 => "1111111000101001101001",
			666 => "0000000110011100101100",
			667 => "0000010111100100010100",
			668 => "0000000010101100001100",
			669 => "0011000100000000000100",
			670 => "0000000000101011000101",
			671 => "0011000110000100000100",
			672 => "0000001000101011000101",
			673 => "0000000000101011000101",
			674 => "0000010111100100000100",
			675 => "1111111000101011000101",
			676 => "0000000000101011000101",
			677 => "0001100000111100000100",
			678 => "0000000000101011000101",
			679 => "0000101110010000010000",
			680 => "0011001100110000000100",
			681 => "0000000000101011000101",
			682 => "0000011001011000001000",
			683 => "0001011101000100000100",
			684 => "0000001000101011000101",
			685 => "0000000000101011000101",
			686 => "0000000000101011000101",
			687 => "0000000000101011000101",
			688 => "1111111000101011000101",
			689 => "0000000110011100101000",
			690 => "0011000100000000000100",
			691 => "0000000000101100011011",
			692 => "0011111010011100001100",
			693 => "0010010000111100001000",
			694 => "0010010000111100000100",
			695 => "0000000000101100011011",
			696 => "0000000000101100011011",
			697 => "0000001000101100011011",
			698 => "0010101001100100001000",
			699 => "0000011101101000000100",
			700 => "0000000000101100011011",
			701 => "0000000000101100011011",
			702 => "0011101010001000001100",
			703 => "0011001100110000000100",
			704 => "0000000000101100011011",
			705 => "0000111001100000000100",
			706 => "0000000000101100011011",
			707 => "0000000000101100011011",
			708 => "0000000000101100011011",
			709 => "1111111000101100011011",
			710 => "0000000000101100011101",
			711 => "0000000000101100100001",
			712 => "0000000000101100100101",
			713 => "0000000000101100101001",
			714 => "0000000000101100101101",
			715 => "0000000000101100110001",
			716 => "0000000000101100110101",
			717 => "0000000000101100111001",
			718 => "0000000000101100111101",
			719 => "0000000000101101000001",
			720 => "0000000000101101000101",
			721 => "0000000000101101001001",
			722 => "0000000000101101001101",
			723 => "0000000000101101010001",
			724 => "0000000000101101010101",
			725 => "0000000000101101011001",
			726 => "0000000000101101011101",
			727 => "0000000000101101100001",
			728 => "0000000000101101100101",
			729 => "0000000000101101101001",
			730 => "0000000000101101101101",
			731 => "0000000000101101110001",
			732 => "0000000010101100000100",
			733 => "0000000000101101111101",
			734 => "0000000000101101111101",
			735 => "0011001100110000000100",
			736 => "0000000000101110001001",
			737 => "0000000000101110001001",
			738 => "0000101000000000000100",
			739 => "0000000000101110010101",
			740 => "0000000000101110010101",
			741 => "0001000111001000000100",
			742 => "0000000000101110100001",
			743 => "0000000000101110100001",
			744 => "0011111011000000000100",
			745 => "0000000000101110101101",
			746 => "0000000000101110101101",
			747 => "0001000110110100000100",
			748 => "0000000000101110111001",
			749 => "0000000000101110111001",
			750 => "0000101000000000000100",
			751 => "0000000000101111000101",
			752 => "0000000000101111000101",
			753 => "0000100001101000000100",
			754 => "0000000000101111011001",
			755 => "0010011110010100000100",
			756 => "0000000000101111011001",
			757 => "0000000000101111011001",
			758 => "0010010000111100000100",
			759 => "0000000000101111101101",
			760 => "0010011001100100000100",
			761 => "0000000000101111101101",
			762 => "0000000000101111101101",
			763 => "0000000010101100000100",
			764 => "0000000000110000000001",
			765 => "0011111100010100000100",
			766 => "0000000000110000000001",
			767 => "0000000000110000000001",
			768 => "0011001000000000001000",
			769 => "0000111100101100000100",
			770 => "0000000000110000010101",
			771 => "0000000000110000010101",
			772 => "0000000000110000010101",
			773 => "0010101101011000001000",
			774 => "0011000110000100000100",
			775 => "0000001000110000110001",
			776 => "0000000000110000110001",
			777 => "0010010101011100000100",
			778 => "0000000000110000110001",
			779 => "0000000000110000110001",
			780 => "0010010000111100001000",
			781 => "0001000111001000000100",
			782 => "0000000000110001001101",
			783 => "0000000000110001001101",
			784 => "0011110111010000000100",
			785 => "0000000000110001001101",
			786 => "0000000000110001001101",
			787 => "0000101000000000001000",
			788 => "0011000100000000000100",
			789 => "0000000000110001101001",
			790 => "0000000000110001101001",
			791 => "0011001100110000000100",
			792 => "0000000000110001101001",
			793 => "0000000000110001101001",
			794 => "0000101000000000001000",
			795 => "0011000100000000000100",
			796 => "0000000000110010000101",
			797 => "0000000000110010000101",
			798 => "0010010111101000000100",
			799 => "0000000000110010000101",
			800 => "0000000000110010000101",
			801 => "0010010101011100001100",
			802 => "0000100100001000000100",
			803 => "0000000000110010100001",
			804 => "0000010110101000000100",
			805 => "0000000000110010100001",
			806 => "0000000000110010100001",
			807 => "0000000000110010100001",
			808 => "0000010110101000000100",
			809 => "0000000000110010111101",
			810 => "0011100111110000001000",
			811 => "0001111101100000000100",
			812 => "0000000000110010111101",
			813 => "0000000000110010111101",
			814 => "0000000000110010111101",
			815 => "0001000111010000000100",
			816 => "0000000000110011011001",
			817 => "0000000010101100000100",
			818 => "0000000000110011011001",
			819 => "0011111010011100000100",
			820 => "0000000000110011011001",
			821 => "0000000000110011011001",
			822 => "0000000010101100001000",
			823 => "0011000110000100000100",
			824 => "0000000000110011111101",
			825 => "0000000000110011111101",
			826 => "0000010111100100001000",
			827 => "0011001110001100000100",
			828 => "0000000000110011111101",
			829 => "0000000000110011111101",
			830 => "0000000000110011111101",
			831 => "0000000010101100001000",
			832 => "0011000110000100000100",
			833 => "0000000000110100100001",
			834 => "0000000000110100100001",
			835 => "0000010111100100001000",
			836 => "0011001110001100000100",
			837 => "0000000000110100100001",
			838 => "0000000000110100100001",
			839 => "0000000000110100100001",
			840 => "0000100000110100010000",
			841 => "0000010111100100001000",
			842 => "0010001001111100000100",
			843 => "0000000000110101000101",
			844 => "0000000000110101000101",
			845 => "0011101101010100000100",
			846 => "0000000000110101000101",
			847 => "0000000000110101000101",
			848 => "0000000000110101000101",
			849 => "0011111001001000001100",
			850 => "0011000100000000000100",
			851 => "0000000000110101110001",
			852 => "0000001010000000000100",
			853 => "0000000000110101110001",
			854 => "0000000000110101110001",
			855 => "0010010111101000001000",
			856 => "0000011101101000000100",
			857 => "0000000000110101110001",
			858 => "0000000000110101110001",
			859 => "0000000000110101110001",
			860 => "0010010000111100000100",
			861 => "0000000000110110010101",
			862 => "0010011001100100001100",
			863 => "0011010010011100001000",
			864 => "0011011001110100000100",
			865 => "0000000000110110010101",
			866 => "0000000000110110010101",
			867 => "0000000000110110010101",
			868 => "0000000000110110010101",
			869 => "0010010000111100000100",
			870 => "0000000000110110111001",
			871 => "0010011001100100001100",
			872 => "0011010010011100001000",
			873 => "0011010110100100000100",
			874 => "0000000000110110111001",
			875 => "0000000000110110111001",
			876 => "0000000000110110111001",
			877 => "0000000000110110111001",
			878 => "0010110101101100001000",
			879 => "0010100100110100000100",
			880 => "0000000000110111100101",
			881 => "0000000000110111100101",
			882 => "0000000110011100001100",
			883 => "0010010000111100000100",
			884 => "0000000000110111100101",
			885 => "0011101010001000000100",
			886 => "0000000000110111100101",
			887 => "0000000000110111100101",
			888 => "0000000000110111100101",
			889 => "0000010110101000010000",
			890 => "0000100100001000000100",
			891 => "0000000000111000010001",
			892 => "0010110000001100001000",
			893 => "0001110110000100000100",
			894 => "0000000000111000010001",
			895 => "0000000000111000010001",
			896 => "0000000000111000010001",
			897 => "0001000110110100000100",
			898 => "0000001000111000010001",
			899 => "0000000000111000010001",
			900 => "0011001100110000001000",
			901 => "0000010111100100000100",
			902 => "0000000000111000111101",
			903 => "0000000000111000111101",
			904 => "0000011001011000001100",
			905 => "0011001000000000001000",
			906 => "0010011101011100000100",
			907 => "0000000000111000111101",
			908 => "0000000000111000111101",
			909 => "0000000000111000111101",
			910 => "0000000000111000111101",
			911 => "0000010110101000001000",
			912 => "0010110000001100000100",
			913 => "0000000000111001101001",
			914 => "0000000000111001101001",
			915 => "0000011001011000001100",
			916 => "0001011101000100001000",
			917 => "0001010011100000000100",
			918 => "0000000000111001101001",
			919 => "0000000000111001101001",
			920 => "0000000000111001101001",
			921 => "0000000000111001101001",
			922 => "0000000110011000010100",
			923 => "0010010000111100001100",
			924 => "0011100100001000000100",
			925 => "0000000000111010010101",
			926 => "0001111101100000000100",
			927 => "0000000000111010010101",
			928 => "0000000000111010010101",
			929 => "0011111011011100000100",
			930 => "0000000000111010010101",
			931 => "0000000000111010010101",
			932 => "0000000000111010010101",
			933 => "0000010110101000001100",
			934 => "0000110100001000000100",
			935 => "0000000000111011001001",
			936 => "0001110110000100000100",
			937 => "0000000000111011001001",
			938 => "0000000000111011001001",
			939 => "0000011001011000001100",
			940 => "0000111001100000001000",
			941 => "0001111001110000000100",
			942 => "0000000000111011001001",
			943 => "0000000000111011001001",
			944 => "0000000000111011001001",
			945 => "0000000000111011001001",
			946 => "0000000110011000010100",
			947 => "0011100100010000010000",
			948 => "0011000100000000001000",
			949 => "0011111101111000000100",
			950 => "0000001000111011110101",
			951 => "0000000000111011110101",
			952 => "0011111011011100000100",
			953 => "0000001000111011110101",
			954 => "0000001000111011110101",
			955 => "0000011000111011110101",
			956 => "1111111000111011110101",
			957 => "0000100001001000010100",
			958 => "0001001001001000000100",
			959 => "0000000000111100101001",
			960 => "0000010111100100001100",
			961 => "0001111110001100001000",
			962 => "0001101001011000000100",
			963 => "0000000000111100101001",
			964 => "0000000000111100101001",
			965 => "0000000000111100101001",
			966 => "0000000000111100101001",
			967 => "0001110111010000000100",
			968 => "1111111000111100101001",
			969 => "0000000000111100101001",
			970 => "0001000110110100010100",
			971 => "0010010101011100010000",
			972 => "0000111010111100000100",
			973 => "0000000000111101011101",
			974 => "0000010110101000001000",
			975 => "0001111101100000000100",
			976 => "0000000000111101011101",
			977 => "0000000000111101011101",
			978 => "0000000000111101011101",
			979 => "0000000000111101011101",
			980 => "0010010111101000000100",
			981 => "0000000000111101011101",
			982 => "0000000000111101011101",
			983 => "0000010110101000001000",
			984 => "0010110000001100000100",
			985 => "0000000000111110010001",
			986 => "0000000000111110010001",
			987 => "0000011001011000010000",
			988 => "0001011110101000001100",
			989 => "0011001000000000001000",
			990 => "0001010011100000000100",
			991 => "0000000000111110010001",
			992 => "0000000000111110010001",
			993 => "0000000000111110010001",
			994 => "0000000000111110010001",
			995 => "0000000000111110010001",
			996 => "0001001100010100010100",
			997 => "0001001001001000000100",
			998 => "0000000000111110111101",
			999 => "0010010000111100000100",
			1000 => "0000000000111110111101",
			1001 => "0011111010011100000100",
			1002 => "0000000000111110111101",
			1003 => "0000010111100100000100",
			1004 => "0000000000111110111101",
			1005 => "0000000000111110111101",
			1006 => "1111111000111110111101",
			1007 => "0000000110011000011000",
			1008 => "0001000110110100001100",
			1009 => "0011101011000000000100",
			1010 => "0000001001000000000001",
			1011 => "0011011111011100000100",
			1012 => "0000000001000000000001",
			1013 => "0000001001000000000001",
			1014 => "0011000110000100000100",
			1015 => "1111110001000000000001",
			1016 => "0000011011101000000100",
			1017 => "0000000001000000000001",
			1018 => "0000001001000000000001",
			1019 => "0001001100010100001000",
			1020 => "0000001100011100000100",
			1021 => "1111111001000000000001",
			1022 => "0000011001000000000001",
			1023 => "1111111001000000000001",
			1024 => "0000010110101000001100",
			1025 => "0010110000001100001000",
			1026 => "0001110110000100000100",
			1027 => "0000000001000000111101",
			1028 => "0000000001000000111101",
			1029 => "0000000001000000111101",
			1030 => "0000011001011000010000",
			1031 => "0001011110101000001100",
			1032 => "0011001000000000001000",
			1033 => "0001111001110000000100",
			1034 => "0000000001000000111101",
			1035 => "0000000001000000111101",
			1036 => "0000000001000000111101",
			1037 => "0000000001000000111101",
			1038 => "0000000001000000111101",
			1039 => "0000010110101000001100",
			1040 => "0011100100001000000100",
			1041 => "0000000001000001111001",
			1042 => "0010110000001100000100",
			1043 => "0000000001000001111001",
			1044 => "0000000001000001111001",
			1045 => "0000011001011000010000",
			1046 => "0011101010001000001100",
			1047 => "0001011101000100001000",
			1048 => "0001010011100000000100",
			1049 => "0000000001000001111001",
			1050 => "0000000001000001111001",
			1051 => "0000000001000001111001",
			1052 => "0000000001000001111001",
			1053 => "0000000001000001111001",
			1054 => "0000000110011000011000",
			1055 => "0011111011000000001000",
			1056 => "0000011001111000000100",
			1057 => "0000000001000010101101",
			1058 => "0000001001000010101101",
			1059 => "0010010101011100000100",
			1060 => "1111111001000010101101",
			1061 => "0011110010001000000100",
			1062 => "0000001001000010101101",
			1063 => "0000011011101000000100",
			1064 => "1111111001000010101101",
			1065 => "0000001001000010101101",
			1066 => "1111111001000010101101",
			1067 => "0000000110011000010100",
			1068 => "0011000100000000000100",
			1069 => "0000000001000011110001",
			1070 => "0000100000110100001100",
			1071 => "0000111001010100001000",
			1072 => "0011111011011100000100",
			1073 => "0000001001000011110001",
			1074 => "0000001001000011110001",
			1075 => "0000010001000011110001",
			1076 => "1111111001000011110001",
			1077 => "0001001001100000001100",
			1078 => "0010100111101100000100",
			1079 => "1111111001000011110001",
			1080 => "0010000111110100000100",
			1081 => "0000011001000011110001",
			1082 => "0000000001000011110001",
			1083 => "1111111001000011110001",
			1084 => "0010101001111100011100",
			1085 => "0000010111100100010100",
			1086 => "0000110110100100001000",
			1087 => "0011000100000000000100",
			1088 => "0000000001000100101101",
			1089 => "0000001001000100101101",
			1090 => "0001111110001100001000",
			1091 => "0001101001011000000100",
			1092 => "1111111001000100101101",
			1093 => "0000000001000100101101",
			1094 => "0000000001000100101101",
			1095 => "0000100001001000000100",
			1096 => "0000001001000100101101",
			1097 => "0000000001000100101101",
			1098 => "1111111001000100101101",
			1099 => "0000100001101000000100",
			1100 => "0000000001000101100001",
			1101 => "0000010111100100000100",
			1102 => "1111111001000101100001",
			1103 => "0001001001100000010000",
			1104 => "0001110001101000001000",
			1105 => "0011110000110100000100",
			1106 => "0000000001000101100001",
			1107 => "0000000001000101100001",
			1108 => "0010100111101100000100",
			1109 => "0000000001000101100001",
			1110 => "0000000001000101100001",
			1111 => "0000000001000101100001",
			1112 => "0010101001111100011000",
			1113 => "0011110000110100010100",
			1114 => "0011000100000000000100",
			1115 => "0000000001000110100101",
			1116 => "0011110101110100001100",
			1117 => "0011110110110100001000",
			1118 => "0011111011011100000100",
			1119 => "0000001001000110100101",
			1120 => "0000000001000110100101",
			1121 => "0000000001000110100101",
			1122 => "0000010001000110100101",
			1123 => "1111111001000110100101",
			1124 => "0001001100010100001000",
			1125 => "0001001110010000000100",
			1126 => "1111111001000110100101",
			1127 => "0000000001000110100101",
			1128 => "1111111001000110100101",
			1129 => "0000000110011100100000",
			1130 => "0000010111100100010000",
			1131 => "0011111001001000001000",
			1132 => "0011000110000100000100",
			1133 => "0000001001000111101001",
			1134 => "0000000001000111101001",
			1135 => "0000010111100100000100",
			1136 => "1111111001000111101001",
			1137 => "0000000001000111101001",
			1138 => "0011101010001000001100",
			1139 => "0010011011001100001000",
			1140 => "0011110000110100000100",
			1141 => "0000001001000111101001",
			1142 => "0000000001000111101001",
			1143 => "0000001001000111101001",
			1144 => "0000000001000111101001",
			1145 => "1111111001000111101001",
			1146 => "0010110101101100001000",
			1147 => "0001000111001000000100",
			1148 => "0000000001001000101101",
			1149 => "0000000001001000101101",
			1150 => "0000100001101000000100",
			1151 => "0000000001001000101101",
			1152 => "0011001000000000001100",
			1153 => "0011001000111100000100",
			1154 => "0000000001001000101101",
			1155 => "0011000110000100000100",
			1156 => "0000000001001000101101",
			1157 => "0000000001001000101101",
			1158 => "0011001000000000001000",
			1159 => "0010110101100100000100",
			1160 => "0000000001001000101101",
			1161 => "0000000001001000101101",
			1162 => "0000000001001000101101",
			1163 => "0000000110011100100000",
			1164 => "0000000010101100001100",
			1165 => "0011000110000100000100",
			1166 => "0000001001001001110001",
			1167 => "0011000110000100000100",
			1168 => "1111111001001001110001",
			1169 => "0000000001001001110001",
			1170 => "0010011011111100000100",
			1171 => "1111111001001001110001",
			1172 => "0011111010001000001100",
			1173 => "0011001100110000000100",
			1174 => "0000000001001001110001",
			1175 => "0001111101111000000100",
			1176 => "0000000001001001110001",
			1177 => "0000001001001001110001",
			1178 => "0000000001001001110001",
			1179 => "1111111001001001110001",
			1180 => "0010101001111100100100",
			1181 => "0001000110110100010100",
			1182 => "0001111001110000000100",
			1183 => "0000000001001011010101",
			1184 => "0011011000011000000100",
			1185 => "0000001001001011010101",
			1186 => "0011011010011100000100",
			1187 => "0000000001001011010101",
			1188 => "0011011010011100000100",
			1189 => "0000000001001011010101",
			1190 => "0000001001001011010101",
			1191 => "0010010111101000001000",
			1192 => "0001011111011100000100",
			1193 => "1111111001001011010101",
			1194 => "0000000001001011010101",
			1195 => "0011100111110000000100",
			1196 => "0000001001001011010101",
			1197 => "0000000001001011010101",
			1198 => "0001001001100000001100",
			1199 => "0010100111101100000100",
			1200 => "1111111001001011010101",
			1201 => "0001000110010000000100",
			1202 => "0000000001001011010101",
			1203 => "0000111001001011010101",
			1204 => "1111111001001011010101",
			1205 => "0000000110011000100000",
			1206 => "0000100111010000010100",
			1207 => "0001111001110000000100",
			1208 => "0000000001001100111001",
			1209 => "0000110110100100000100",
			1210 => "0000001001001100111001",
			1211 => "0011011010011100000100",
			1212 => "1111111001001100111001",
			1213 => "0011011010011100000100",
			1214 => "0000000001001100111001",
			1215 => "0000001001001100111001",
			1216 => "0000010111100100000100",
			1217 => "1111111001001100111001",
			1218 => "0011100101110100000100",
			1219 => "0000001001001100111001",
			1220 => "0000000001001100111001",
			1221 => "0010000111110100010000",
			1222 => "0010100111101100000100",
			1223 => "1111111001001100111001",
			1224 => "0000000110011100000100",
			1225 => "0000000001001100111001",
			1226 => "0010100111101100000100",
			1227 => "0000011001001100111001",
			1228 => "0000000001001100111001",
			1229 => "1111111001001100111001",
			1230 => "0010000111110100101000",
			1231 => "0000010111100100011000",
			1232 => "0011100100001000001000",
			1233 => "0000010010001100000100",
			1234 => "0000000001001110001101",
			1235 => "0000000001001110001101",
			1236 => "0000010110101000000100",
			1237 => "0000000001001110001101",
			1238 => "0000010110101000000100",
			1239 => "0000000001001110001101",
			1240 => "0001110110000100000100",
			1241 => "0000000001001110001101",
			1242 => "0000000001001110001101",
			1243 => "0011101010001000001100",
			1244 => "0001011110101000001000",
			1245 => "0000101110010000000100",
			1246 => "0000000001001110001101",
			1247 => "0000000001001110001101",
			1248 => "0000000001001110001101",
			1249 => "0000000001001110001101",
			1250 => "1111111001001110001101",
			1251 => "0000000110011100100000",
			1252 => "0010110101100100011000",
			1253 => "0011111011000000000100",
			1254 => "0000001001001111010001",
			1255 => "0010010101011100000100",
			1256 => "1111111001001111010001",
			1257 => "0011110010001000000100",
			1258 => "0000001001001111010001",
			1259 => "0001101011111100000100",
			1260 => "0000000001001111010001",
			1261 => "0001101110010100000100",
			1262 => "0000000001001111010001",
			1263 => "0000000001001111010001",
			1264 => "0011101010001000000100",
			1265 => "0000001001001111010001",
			1266 => "0000000001001111010001",
			1267 => "1111111001001111010001",
			1268 => "0001001001100000100100",
			1269 => "0011001000000000011100",
			1270 => "0000100000110100011000",
			1271 => "0000010111100100010000",
			1272 => "0001001001001000001000",
			1273 => "0011000100000000000100",
			1274 => "0000000001010000011101",
			1275 => "0000001001010000011101",
			1276 => "0010010000111100000100",
			1277 => "1111111001010000011101",
			1278 => "0000000001010000011101",
			1279 => "0011110010001000000100",
			1280 => "0000001001010000011101",
			1281 => "0000000001010000011101",
			1282 => "1111111001010000011101",
			1283 => "0010110101100100000100",
			1284 => "0000000001010000011101",
			1285 => "0000011001010000011101",
			1286 => "1111111001010000011101",
			1287 => "0001001001100000100100",
			1288 => "0001000111010000001000",
			1289 => "0011000100000000000100",
			1290 => "0000000001010001101001",
			1291 => "0000001001010001101001",
			1292 => "0000011101101000001000",
			1293 => "0011001000111100000100",
			1294 => "0000000001010001101001",
			1295 => "0000000001010001101001",
			1296 => "0011101010001000010000",
			1297 => "0011000110000100000100",
			1298 => "0000000001010001101001",
			1299 => "0000011001011000001000",
			1300 => "0000111001100000000100",
			1301 => "0000000001010001101001",
			1302 => "0000000001010001101001",
			1303 => "0000000001010001101001",
			1304 => "0000000001010001101001",
			1305 => "1111111001010001101001",
			1306 => "0001001100010100100000",
			1307 => "0000010010001100000100",
			1308 => "1111111001010010101101",
			1309 => "0000100001001000010100",
			1310 => "0000010110101000010000",
			1311 => "0011110111001000001100",
			1312 => "0011100100001000000100",
			1313 => "0000001001010010101101",
			1314 => "0011100001111100000100",
			1315 => "0000000001010010101101",
			1316 => "0000001001010010101101",
			1317 => "1111111001010010101101",
			1318 => "0000001001010010101101",
			1319 => "0001110110100100000100",
			1320 => "1111111001010010101101",
			1321 => "0000010001010010101101",
			1322 => "1111111001010010101101",
			1323 => "0010100111101100101000",
			1324 => "0000010111100100010000",
			1325 => "0011100100001000001000",
			1326 => "0000010010001100000100",
			1327 => "0000000001010100000001",
			1328 => "0000000001010100000001",
			1329 => "0000010110101000000100",
			1330 => "0000000001010100000001",
			1331 => "0000000001010100000001",
			1332 => "0000111001100000010100",
			1333 => "0010011011111100000100",
			1334 => "0000000001010100000001",
			1335 => "0011001100110000000100",
			1336 => "0000000001010100000001",
			1337 => "0001011101000100001000",
			1338 => "0000011001011000000100",
			1339 => "0000000001010100000001",
			1340 => "0000000001010100000001",
			1341 => "0000000001010100000001",
			1342 => "0000000001010100000001",
			1343 => "0000000001010100000001",
			1344 => "0001001001100000100100",
			1345 => "0000011001111000001000",
			1346 => "0000100100001000000100",
			1347 => "0000000001010101001101",
			1348 => "1111111001010101001101",
			1349 => "0010110100001000000100",
			1350 => "0000001001010101001101",
			1351 => "0011001100110000001000",
			1352 => "0000010111100100000100",
			1353 => "1111111001010101001101",
			1354 => "0000000001010101001101",
			1355 => "0000101110010000001100",
			1356 => "0000010111100100000100",
			1357 => "0000000001010101001101",
			1358 => "0001100000111100000100",
			1359 => "0000000001010101001101",
			1360 => "0000001001010101001101",
			1361 => "0000000001010101001101",
			1362 => "1111111001010101001101",
			1363 => "0010000111110100101000",
			1364 => "0000010111100100010000",
			1365 => "0000000010101100001100",
			1366 => "0011000100000000000100",
			1367 => "0000000001010110100001",
			1368 => "0011000110000100000100",
			1369 => "0000001001010110100001",
			1370 => "0000000001010110100001",
			1371 => "1111111001010110100001",
			1372 => "0011101010001000010100",
			1373 => "0001100000111100000100",
			1374 => "0000000001010110100001",
			1375 => "0000010111100100000100",
			1376 => "0000000001010110100001",
			1377 => "0011001100110000000100",
			1378 => "0000000001010110100001",
			1379 => "0001011101000100000100",
			1380 => "0000001001010110100001",
			1381 => "0000000001010110100001",
			1382 => "0000000001010110100001",
			1383 => "1111111001010110100001",
			1384 => "0000000110011100100100",
			1385 => "0011000100000000000100",
			1386 => "0000000001010111101101",
			1387 => "0011111010011100001100",
			1388 => "0010010000111100001000",
			1389 => "0010010000111100000100",
			1390 => "0000000001010111101101",
			1391 => "0000000001010111101101",
			1392 => "0000001001010111101101",
			1393 => "0011001100110000000100",
			1394 => "0000000001010111101101",
			1395 => "0011101010001000001100",
			1396 => "0010011110010100000100",
			1397 => "0000000001010111101101",
			1398 => "0000111001100000000100",
			1399 => "0000000001010111101101",
			1400 => "0000000001010111101101",
			1401 => "0000000001010111101101",
			1402 => "1111111001010111101101",
			1403 => "0000000110011100110000",
			1404 => "0000010111100100011000",
			1405 => "0000000010101100010000",
			1406 => "0011000100000000000100",
			1407 => "0000000001011001010011",
			1408 => "0011000110000100000100",
			1409 => "0000001001011001010011",
			1410 => "0011011010011100000100",
			1411 => "0000000001011001010011",
			1412 => "0000000001011001010011",
			1413 => "0000010111100100000100",
			1414 => "1111111001011001010011",
			1415 => "0000000001011001010011",
			1416 => "0011101010001000010100",
			1417 => "0001100000111100000100",
			1418 => "0000000001011001010011",
			1419 => "0011001100110000000100",
			1420 => "0000000001011001010011",
			1421 => "0001011101000100001000",
			1422 => "0000111001100000000100",
			1423 => "0000001001011001010011",
			1424 => "0000000001011001010011",
			1425 => "0000000001011001010011",
			1426 => "0000000001011001010011",
			1427 => "1111111001011001010011",
			1428 => "0000000001011001010101",
			1429 => "0000000001011001011001",
			1430 => "0000000001011001011101",
			1431 => "0000000001011001100001",
			1432 => "0000000001011001100101",
			1433 => "0000000001011001101001",
			1434 => "0000000001011001101101",
			1435 => "0000000001011001110001",
			1436 => "0000000001011001110101",
			1437 => "0000000001011001111001",
			1438 => "0000000001011001111101",
			1439 => "0000000001011010000001",
			1440 => "0000000001011010000101",
			1441 => "0000000001011010001001",
			1442 => "0000000001011010001101",
			1443 => "0000000001011010010001",
			1444 => "0000000001011010010101",
			1445 => "0000000001011010011001",
			1446 => "0000000001011010011101",
			1447 => "0000000001011010100001",
			1448 => "0000000001011010100101",
			1449 => "0000000010101100000100",
			1450 => "0000000001011010110001",
			1451 => "0000000001011010110001",
			1452 => "0000000010101100000100",
			1453 => "0000000001011010111101",
			1454 => "0000000001011010111101",
			1455 => "0011001100110000000100",
			1456 => "0000000001011011001001",
			1457 => "0000000001011011001001",
			1458 => "0001000111001000000100",
			1459 => "0000000001011011010101",
			1460 => "0000000001011011010101",
			1461 => "0011111011000000000100",
			1462 => "0000000001011011100001",
			1463 => "0000000001011011100001",
			1464 => "0001000110110100000100",
			1465 => "0000000001011011101101",
			1466 => "0000000001011011101101",
			1467 => "0000101000000000000100",
			1468 => "0000000001011011111001",
			1469 => "0000000001011011111001",
			1470 => "0001000111010000000100",
			1471 => "0000000001011100001101",
			1472 => "0001111100101000000100",
			1473 => "0000000001011100001101",
			1474 => "0000000001011100001101",
			1475 => "0001000111010000000100",
			1476 => "0000000001011100100001",
			1477 => "0010011110010100000100",
			1478 => "0000000001011100100001",
			1479 => "0000000001011100100001",
			1480 => "0011011010011100000100",
			1481 => "0000000001011100110101",
			1482 => "0011010010011100000100",
			1483 => "0000000001011100110101",
			1484 => "0000000001011100110101",
			1485 => "0000101000000000001000",
			1486 => "0011111010111100000100",
			1487 => "0000000001011101001001",
			1488 => "0000000001011101001001",
			1489 => "0000000001011101001001",
			1490 => "0010010000111100000100",
			1491 => "0000000001011101011101",
			1492 => "0010011001100100000100",
			1493 => "0000000001011101011101",
			1494 => "0000000001011101011101",
			1495 => "0000101000000000001000",
			1496 => "0000010110101000000100",
			1497 => "0000000001011101111001",
			1498 => "0000001001011101111001",
			1499 => "0010010101011100000100",
			1500 => "0000000001011101111001",
			1501 => "0000000001011101111001",
			1502 => "0010010000111100001000",
			1503 => "0001000111001000000100",
			1504 => "0000000001011110010101",
			1505 => "0000000001011110010101",
			1506 => "0011110111010000000100",
			1507 => "0000000001011110010101",
			1508 => "0000000001011110010101",
			1509 => "0000101000000000001000",
			1510 => "0011000100000000000100",
			1511 => "0000000001011110110001",
			1512 => "0000000001011110110001",
			1513 => "0001110111010000000100",
			1514 => "0000000001011110110001",
			1515 => "0000000001011110110001",
			1516 => "0001000111010000000100",
			1517 => "0000000001011111001101",
			1518 => "0000010111100100001000",
			1519 => "0001011111011100000100",
			1520 => "0000000001011111001101",
			1521 => "0000000001011111001101",
			1522 => "0000000001011111001101",
			1523 => "0010010101011100001100",
			1524 => "0000100100001000000100",
			1525 => "0000000001011111101001",
			1526 => "0000010110101000000100",
			1527 => "0000000001011111101001",
			1528 => "0000000001011111101001",
			1529 => "0000000001011111101001",
			1530 => "0010010000111100001100",
			1531 => "0001000111001000000100",
			1532 => "0000000001100000000101",
			1533 => "0000010110101000000100",
			1534 => "0000000001100000000101",
			1535 => "0000000001100000000101",
			1536 => "0000000001100000000101",
			1537 => "0001000111010000000100",
			1538 => "0000000001100000100001",
			1539 => "0000000010101100000100",
			1540 => "0000000001100000100001",
			1541 => "0011111010011100000100",
			1542 => "0000000001100000100001",
			1543 => "0000000001100000100001",
			1544 => "0000000010101100001000",
			1545 => "0011000110000100000100",
			1546 => "0000000001100001000101",
			1547 => "0000000001100001000101",
			1548 => "0000010111100100001000",
			1549 => "0011001110001100000100",
			1550 => "0000000001100001000101",
			1551 => "0000000001100001000101",
			1552 => "0000000001100001000101",
			1553 => "0000010110101000001100",
			1554 => "0011100100001000000100",
			1555 => "0000000001100001101001",
			1556 => "0010110000001100000100",
			1557 => "0000000001100001101001",
			1558 => "0000000001100001101001",
			1559 => "0011100110100100000100",
			1560 => "0000000001100001101001",
			1561 => "0000000001100001101001",
			1562 => "0000100000110100010000",
			1563 => "0000010111100100001000",
			1564 => "0010001001111100000100",
			1565 => "0000000001100010001101",
			1566 => "0000000001100010001101",
			1567 => "0011101101010100000100",
			1568 => "0000000001100010001101",
			1569 => "0000000001100010001101",
			1570 => "0000000001100010001101",
			1571 => "0010000111110100010000",
			1572 => "0010011101101000000100",
			1573 => "0000000001100010110001",
			1574 => "0000111001100000001000",
			1575 => "0010010000111100000100",
			1576 => "0000000001100010110001",
			1577 => "0000000001100010110001",
			1578 => "0000000001100010110001",
			1579 => "0000000001100010110001",
			1580 => "0010010000111100000100",
			1581 => "0000000001100011010101",
			1582 => "0010011001100100001100",
			1583 => "0011010010011100001000",
			1584 => "0011011001110100000100",
			1585 => "0000000001100011010101",
			1586 => "0000000001100011010101",
			1587 => "0000000001100011010101",
			1588 => "0000000001100011010101",
			1589 => "0010010000111100000100",
			1590 => "0000000001100011111001",
			1591 => "0010011001100100001100",
			1592 => "0011010010011100001000",
			1593 => "0011010110100100000100",
			1594 => "0000000001100011111001",
			1595 => "0000000001100011111001",
			1596 => "0000000001100011111001",
			1597 => "0000000001100011111001",
			1598 => "0010010101011100001000",
			1599 => "0000010111100100000100",
			1600 => "0000000001100100100101",
			1601 => "0000000001100100100101",
			1602 => "0000011001011000001100",
			1603 => "0001011110101000001000",
			1604 => "0001111101100000000100",
			1605 => "0000000001100100100101",
			1606 => "0000000001100100100101",
			1607 => "0000000001100100100101",
			1608 => "0000000001100100100101",
			1609 => "0000010110101000010000",
			1610 => "0011110001111100000100",
			1611 => "0000000001100101010001",
			1612 => "0010110000001100001000",
			1613 => "0001110110000100000100",
			1614 => "0000000001100101010001",
			1615 => "0000000001100101010001",
			1616 => "0000000001100101010001",
			1617 => "0011111011011100000100",
			1618 => "0000001001100101010001",
			1619 => "0000000001100101010001",
			1620 => "0011001100110000001000",
			1621 => "0000010111100100000100",
			1622 => "0000000001100101111101",
			1623 => "0000000001100101111101",
			1624 => "0000011001011000001100",
			1625 => "0011001000000000001000",
			1626 => "0010011101011100000100",
			1627 => "0000000001100101111101",
			1628 => "0000000001100101111101",
			1629 => "0000000001100101111101",
			1630 => "0000000001100101111101",
			1631 => "0010010000111100001100",
			1632 => "0000100100001000001000",
			1633 => "0010001000010000000100",
			1634 => "0000000001100110110001",
			1635 => "0000000001100110110001",
			1636 => "1111111001100110110001",
			1637 => "0000100001001000001000",
			1638 => "0010010101011100000100",
			1639 => "0000000001100110110001",
			1640 => "0000000001100110110001",
			1641 => "0001110111010000000100",
			1642 => "0000000001100110110001",
			1643 => "0000000001100110110001",
			1644 => "0010010101011100001100",
			1645 => "0011100100001000000100",
			1646 => "0000000001100111100101",
			1647 => "0000010111100100000100",
			1648 => "0000000001100111100101",
			1649 => "0000000001100111100101",
			1650 => "0000011001011000001100",
			1651 => "0011101010001000001000",
			1652 => "0001111101100000000100",
			1653 => "0000000001100111100101",
			1654 => "0000000001100111100101",
			1655 => "0000000001100111100101",
			1656 => "0000000001100111100101",
			1657 => "0011001100110000001100",
			1658 => "0011110001111100000100",
			1659 => "0000000001101000011001",
			1660 => "0000010111100100000100",
			1661 => "0000000001101000011001",
			1662 => "0000000001101000011001",
			1663 => "0000010110101000000100",
			1664 => "0000000001101000011001",
			1665 => "0000101110010000001000",
			1666 => "0000011001011000000100",
			1667 => "0000000001101000011001",
			1668 => "0000000001101000011001",
			1669 => "0000000001101000011001",
			1670 => "0000000110011000010000",
			1671 => "0011000100000000000100",
			1672 => "0000000001101001010101",
			1673 => "0011110000110100001000",
			1674 => "0000100101110100000100",
			1675 => "0000001001101001010101",
			1676 => "0000011001101001010101",
			1677 => "1111111001101001010101",
			1678 => "0001001001100000001100",
			1679 => "0010000111110100000100",
			1680 => "1111111001101001010101",
			1681 => "0010000111110100000100",
			1682 => "0000110001101001010101",
			1683 => "0000000001101001010101",
			1684 => "1111111001101001010101",
			1685 => "0001001001100000011000",
			1686 => "0010010000111100001100",
			1687 => "0011111011000000001000",
			1688 => "0001111001110000000100",
			1689 => "0000000001101010001001",
			1690 => "0000000001101010001001",
			1691 => "0000000001101010001001",
			1692 => "0001110110000100000100",
			1693 => "0000000001101010001001",
			1694 => "0011101010001000000100",
			1695 => "0000000001101010001001",
			1696 => "0000000001101010001001",
			1697 => "0000000001101010001001",
			1698 => "0000010111100100001000",
			1699 => "0010001001111100000100",
			1700 => "0000000001101010111101",
			1701 => "0000000001101010111101",
			1702 => "0000101110010000010000",
			1703 => "0001100000111100000100",
			1704 => "0000000001101010111101",
			1705 => "0000011001011000001000",
			1706 => "0001011110101000000100",
			1707 => "0000000001101010111101",
			1708 => "0000000001101010111101",
			1709 => "0000000001101010111101",
			1710 => "0000000001101010111101",
			1711 => "0010010000111100001000",
			1712 => "0001111110001100000100",
			1713 => "0000000001101011110001",
			1714 => "0000000001101011110001",
			1715 => "0010011001100100010000",
			1716 => "0001011110101000001100",
			1717 => "0001111101100000000100",
			1718 => "0000000001101011110001",
			1719 => "0011001000000000000100",
			1720 => "0000000001101011110001",
			1721 => "0000000001101011110001",
			1722 => "0000000001101011110001",
			1723 => "0000000001101011110001",
			1724 => "0000000010101100000100",
			1725 => "0000000001101100011101",
			1726 => "0000010111100100000100",
			1727 => "0000000001101100011101",
			1728 => "0000101110010000001100",
			1729 => "0001101101111100001000",
			1730 => "0001011101000100000100",
			1731 => "0000000001101100011101",
			1732 => "0000000001101100011101",
			1733 => "0000000001101100011101",
			1734 => "0000000001101100011101",
			1735 => "0000000110011000010100",
			1736 => "0001000110110100001100",
			1737 => "0001001001001000000100",
			1738 => "0000001001101101100001",
			1739 => "0010010101011100000100",
			1740 => "1111111001101101100001",
			1741 => "0000001001101101100001",
			1742 => "0010010111101000000100",
			1743 => "1111111001101101100001",
			1744 => "0000001001101101100001",
			1745 => "0001001001100000001100",
			1746 => "0010100111101100000100",
			1747 => "1111111001101101100001",
			1748 => "0001000110010000000100",
			1749 => "0000000001101101100001",
			1750 => "0000100001101101100001",
			1751 => "1111111001101101100001",
			1752 => "0010010000111100001100",
			1753 => "0000010110101000001000",
			1754 => "0001111110001100000100",
			1755 => "0000000001101110011101",
			1756 => "0000000001101110011101",
			1757 => "0000000001101110011101",
			1758 => "0000011001011000010000",
			1759 => "0001011110101000001100",
			1760 => "0001111101100000000100",
			1761 => "0000000001101110011101",
			1762 => "0011001000000000000100",
			1763 => "0000000001101110011101",
			1764 => "0000000001101110011101",
			1765 => "0000000001101110011101",
			1766 => "0000000001101110011101",
			1767 => "0010010000111100010100",
			1768 => "0001001001001000001100",
			1769 => "0001000111001000000100",
			1770 => "0000000001101111101001",
			1771 => "0001101101011100000100",
			1772 => "0000000001101111101001",
			1773 => "0000000001101111101001",
			1774 => "0000010110101000000100",
			1775 => "1111111001101111101001",
			1776 => "0000000001101111101001",
			1777 => "0011100111110000001100",
			1778 => "0010010101011100000100",
			1779 => "0000000001101111101001",
			1780 => "0000000110011100000100",
			1781 => "0000000001101111101001",
			1782 => "0000000001101111101001",
			1783 => "0001110111010000000100",
			1784 => "0000000001101111101001",
			1785 => "0000000001101111101001",
			1786 => "0000100001001000011000",
			1787 => "0001001001001000000100",
			1788 => "0000000001110000100101",
			1789 => "0010010000111100001000",
			1790 => "0001101001011000000100",
			1791 => "0000000001110000100101",
			1792 => "0000000001110000100101",
			1793 => "0011111010011100000100",
			1794 => "0000000001110000100101",
			1795 => "0011000110000100000100",
			1796 => "0000000001110000100101",
			1797 => "0000000001110000100101",
			1798 => "0001110111010000000100",
			1799 => "1111111001110000100101",
			1800 => "0000000001110000100101",
			1801 => "0000100001001000011100",
			1802 => "0010010101011100010100",
			1803 => "0011110001111100001000",
			1804 => "0000010010001100000100",
			1805 => "0000000001110001101001",
			1806 => "0000000001110001101001",
			1807 => "0010010000111100001000",
			1808 => "0001111101100000000100",
			1809 => "0000000001110001101001",
			1810 => "0000000001110001101001",
			1811 => "0000000001110001101001",
			1812 => "0011110010001000000100",
			1813 => "0000000001110001101001",
			1814 => "0000000001110001101001",
			1815 => "0001110111010000000100",
			1816 => "1111111001110001101001",
			1817 => "0000000001110001101001",
			1818 => "0001001100010100011100",
			1819 => "0000010111100100001100",
			1820 => "0001001001001000001000",
			1821 => "0001101111001100000100",
			1822 => "0000000001110010100101",
			1823 => "0000001001110010100101",
			1824 => "1111111001110010100101",
			1825 => "0011110010001000000100",
			1826 => "0000001001110010100101",
			1827 => "0000110001001000000100",
			1828 => "0000000001110010100101",
			1829 => "0011111010001000000100",
			1830 => "0000000001110010100101",
			1831 => "0000000001110010100101",
			1832 => "1111111001110010100101",
			1833 => "0000010111100100011000",
			1834 => "0011111011000000001100",
			1835 => "0011000100000000000100",
			1836 => "0000000001110011111001",
			1837 => "0001100111101000000100",
			1838 => "0000000001110011111001",
			1839 => "0000000001110011111001",
			1840 => "0011001110001100001000",
			1841 => "0001101001011000000100",
			1842 => "0000000001110011111001",
			1843 => "0000000001110011111001",
			1844 => "0000000001110011111001",
			1845 => "0000101110010000010000",
			1846 => "0001100000111100000100",
			1847 => "0000000001110011111001",
			1848 => "0000011001011000001000",
			1849 => "0011101010001000000100",
			1850 => "0000000001110011111001",
			1851 => "0000000001110011111001",
			1852 => "0000000001110011111001",
			1853 => "0000000001110011111001",
			1854 => "0001001100010100100000",
			1855 => "0000010111100100010000",
			1856 => "0001001001001000001000",
			1857 => "0001101111001100000100",
			1858 => "0000000001110100111101",
			1859 => "0000001001110100111101",
			1860 => "0000010110101000000100",
			1861 => "1111111001110100111101",
			1862 => "0000000001110100111101",
			1863 => "0011110010001000000100",
			1864 => "0000001001110100111101",
			1865 => "0011010101110100000100",
			1866 => "0000000001110100111101",
			1867 => "0011111010001000000100",
			1868 => "0000000001110100111101",
			1869 => "0000000001110100111101",
			1870 => "1111111001110100111101",
			1871 => "0000000110011100100000",
			1872 => "0000010111100100010000",
			1873 => "0011111001001000001000",
			1874 => "0011000110000100000100",
			1875 => "0000001001110110000001",
			1876 => "0000000001110110000001",
			1877 => "0000010111100100000100",
			1878 => "1111111001110110000001",
			1879 => "0000000001110110000001",
			1880 => "0000111001100000001100",
			1881 => "0001100000111100000100",
			1882 => "0000000001110110000001",
			1883 => "0000101110010000000100",
			1884 => "0000001001110110000001",
			1885 => "0000000001110110000001",
			1886 => "0000000001110110000001",
			1887 => "1111111001110110000001",
			1888 => "0000000010101100000100",
			1889 => "0000000001110110110101",
			1890 => "0000010111100100000100",
			1891 => "0000000001110110110101",
			1892 => "0001101101111100010000",
			1893 => "0011101010001000001100",
			1894 => "0001011101000100001000",
			1895 => "0011001100110000000100",
			1896 => "0000000001110110110101",
			1897 => "0000000001110110110101",
			1898 => "0000000001110110110101",
			1899 => "0000000001110110110101",
			1900 => "0000000001110110110101",
			1901 => "0000000110011000011100",
			1902 => "0011110000110100011000",
			1903 => "0011110101110100010100",
			1904 => "0001000110110100001100",
			1905 => "0011110111010000000100",
			1906 => "0000001001111000000001",
			1907 => "0011101010001100000100",
			1908 => "0000000001111000000001",
			1909 => "0000001001111000000001",
			1910 => "0001100101011100000100",
			1911 => "1111111001111000000001",
			1912 => "0000001001111000000001",
			1913 => "0000010001111000000001",
			1914 => "1111111001111000000001",
			1915 => "0001001100010100001000",
			1916 => "0001001110010000000100",
			1917 => "1111111001111000000001",
			1918 => "0000000001111000000001",
			1919 => "1111111001111000000001",
			1920 => "0000000110011000011000",
			1921 => "0010010100110100010100",
			1922 => "0011110001001000010000",
			1923 => "0011000100000000000100",
			1924 => "0000000001111001010101",
			1925 => "0011110110110100001000",
			1926 => "0011111011011100000100",
			1927 => "0000001001111001010101",
			1928 => "0000001001111001010101",
			1929 => "0000010001111001010101",
			1930 => "1111111001111001010101",
			1931 => "0000011001111001010101",
			1932 => "0000000110011100010000",
			1933 => "0010000111110100000100",
			1934 => "1111111001111001010101",
			1935 => "0010000111110100001000",
			1936 => "0010100111101100000100",
			1937 => "0000000001111001010101",
			1938 => "0000010001111001010101",
			1939 => "0000000001111001010101",
			1940 => "1111111001111001010101",
			1941 => "0000000110011000100000",
			1942 => "0000011001111000000100",
			1943 => "0000000001111010110001",
			1944 => "0011110010001000010100",
			1945 => "0000011001111000001000",
			1946 => "0011101100110000000100",
			1947 => "0000001001111010110001",
			1948 => "0000000001111010110001",
			1949 => "0011101011000000000100",
			1950 => "0000001001111010110001",
			1951 => "0011001100110000000100",
			1952 => "0000000001111010110001",
			1953 => "0000001001111010110001",
			1954 => "0001110100001000000100",
			1955 => "1111111001111010110001",
			1956 => "0000001001111010110001",
			1957 => "0000000110011100001100",
			1958 => "0010000111110100000100",
			1959 => "1111111001111010110001",
			1960 => "0010000111110100000100",
			1961 => "0000001001111010110001",
			1962 => "0000000001111010110001",
			1963 => "1111111001111010110001",
			1964 => "0010000111110100101000",
			1965 => "0000010111100100010100",
			1966 => "0010000101010000001100",
			1967 => "0011100100001000000100",
			1968 => "0000000001111100000101",
			1969 => "0011111101010100000100",
			1970 => "0000000001111100000101",
			1971 => "0000000001111100000101",
			1972 => "0010010000111100000100",
			1973 => "0000000001111100000101",
			1974 => "0000000001111100000101",
			1975 => "0011101010001000010000",
			1976 => "0001011110101000001100",
			1977 => "0000111001100000001000",
			1978 => "0000101110010000000100",
			1979 => "0000000001111100000101",
			1980 => "0000000001111100000101",
			1981 => "0000000001111100000101",
			1982 => "0000000001111100000101",
			1983 => "0000000001111100000101",
			1984 => "1111111001111100000101",
			1985 => "0010000111110100100000",
			1986 => "0000011001111000001000",
			1987 => "0000100100001000000100",
			1988 => "0000000001111101001001",
			1989 => "0000000001111101001001",
			1990 => "0011111010011100000100",
			1991 => "0000000001111101001001",
			1992 => "0000010111100100000100",
			1993 => "0000000001111101001001",
			1994 => "0011101010001000001100",
			1995 => "0001100101011100000100",
			1996 => "0000000001111101001001",
			1997 => "0001011110101000000100",
			1998 => "0000000001111101001001",
			1999 => "0000000001111101001001",
			2000 => "0000000001111101001001",
			2001 => "1111111001111101001001",
			2002 => "0001001001100000100100",
			2003 => "0011001000000000011100",
			2004 => "0000100000110100011000",
			2005 => "0000010111100100010000",
			2006 => "0001001001001000001000",
			2007 => "0011000100000000000100",
			2008 => "0000000001111110010101",
			2009 => "0000001001111110010101",
			2010 => "0010010000111100000100",
			2011 => "1111111001111110010101",
			2012 => "0000000001111110010101",
			2013 => "0011110010001000000100",
			2014 => "0000001001111110010101",
			2015 => "0000000001111110010101",
			2016 => "1111111001111110010101",
			2017 => "0010110101100100000100",
			2018 => "0000000001111110010101",
			2019 => "0000010001111110010101",
			2020 => "1111111001111110010101",
			2021 => "0010101001111100011100",
			2022 => "0000011001111000000100",
			2023 => "1111111001111111110001",
			2024 => "0000100000110100010100",
			2025 => "0011111011000000000100",
			2026 => "0000001001111111110001",
			2027 => "0000010111100100000100",
			2028 => "1111111001111111110001",
			2029 => "0001110110000100001000",
			2030 => "0001100000111100000100",
			2031 => "0000001001111111110001",
			2032 => "0000000001111111110001",
			2033 => "0000001001111111110001",
			2034 => "1111111001111111110001",
			2035 => "0001001001100000010000",
			2036 => "0010100111101100000100",
			2037 => "1111111001111111110001",
			2038 => "0010100111101100001000",
			2039 => "0010000111110100000100",
			2040 => "0000000001111111110001",
			2041 => "0000100001111111110001",
			2042 => "0000000001111111110001",
			2043 => "1111111001111111110001",
			2044 => "0010000111110100100000",
			2045 => "0000100001101000000100",
			2046 => "0000000010000000110101",
			2047 => "0000011101101000001000",
			2048 => "0011001000111100000100",
			2049 => "0000000010000000110101",
			2050 => "0000000010000000110101",
			2051 => "0011101010001000010000",
			2052 => "0011000110000100000100",
			2053 => "0000000010000000110101",
			2054 => "0001011110101000001000",
			2055 => "0000101110010000000100",
			2056 => "0000000010000000110101",
			2057 => "0000000010000000110101",
			2058 => "0000000010000000110101",
			2059 => "0000000010000000110101",
			2060 => "1111111010000000110101",
			2061 => "0000010110101000010000",
			2062 => "0000100100001000000100",
			2063 => "0000000010000010011001",
			2064 => "0001110110000100001000",
			2065 => "0010110000001100000100",
			2066 => "1111111010000010011001",
			2067 => "0000000010000010011001",
			2068 => "0000000010000010011001",
			2069 => "0000000010101100000100",
			2070 => "0000000010000010011001",
			2071 => "0000010111100100001100",
			2072 => "0011100110100100000100",
			2073 => "0000000010000010011001",
			2074 => "0001110101101100000100",
			2075 => "0000000010000010011001",
			2076 => "0000000010000010011001",
			2077 => "0000101110010000010000",
			2078 => "0011001100110000000100",
			2079 => "0000000010000010011001",
			2080 => "0010011110010100000100",
			2081 => "0000000010000010011001",
			2082 => "0000011001011000000100",
			2083 => "0000000010000010011001",
			2084 => "0000000010000010011001",
			2085 => "0000000010000010011001",
			2086 => "0001001001100000100100",
			2087 => "0000011001111000001000",
			2088 => "0000100100001000000100",
			2089 => "0000000010000011100101",
			2090 => "1111111010000011100101",
			2091 => "0010110100001000000100",
			2092 => "0000001010000011100101",
			2093 => "0011001100110000001000",
			2094 => "0000010111100100000100",
			2095 => "0000000010000011100101",
			2096 => "0000000010000011100101",
			2097 => "0011101010001000001100",
			2098 => "0000010111100100000100",
			2099 => "0000000010000011100101",
			2100 => "0001100000111100000100",
			2101 => "0000000010000011100101",
			2102 => "0000001010000011100101",
			2103 => "0000000010000011100101",
			2104 => "1111111010000011100101",
			2105 => "0010000111110100101000",
			2106 => "0000011001111000001000",
			2107 => "0011110001111100000100",
			2108 => "0000000010000100111001",
			2109 => "0000000010000100111001",
			2110 => "0011111010011100001100",
			2111 => "0010110100001000000100",
			2112 => "0000001010000100111001",
			2113 => "0010110001111100000100",
			2114 => "0000000010000100111001",
			2115 => "0000000010000100111001",
			2116 => "0000010111100100000100",
			2117 => "0000000010000100111001",
			2118 => "0011101010001000001100",
			2119 => "0001100101011100000100",
			2120 => "0000000010000100111001",
			2121 => "0001011110101000000100",
			2122 => "0000000010000100111001",
			2123 => "0000000010000100111001",
			2124 => "0000000010000100111001",
			2125 => "1111111010000100111001",
			2126 => "0010000111110100101000",
			2127 => "0011001000000000100000",
			2128 => "0000100000110100011100",
			2129 => "0000010111100100010000",
			2130 => "0010000101010000001000",
			2131 => "0011000100000000000100",
			2132 => "0000000010000110001101",
			2133 => "0000001010000110001101",
			2134 => "0000001010100000000100",
			2135 => "0000000010000110001101",
			2136 => "1111111010000110001101",
			2137 => "0001110110000100001000",
			2138 => "0011110110100100000100",
			2139 => "0000001010000110001101",
			2140 => "0000000010000110001101",
			2141 => "0000001010000110001101",
			2142 => "1111111010000110001101",
			2143 => "0000111001100000000100",
			2144 => "0000110010000110001101",
			2145 => "0000000010000110001101",
			2146 => "1111111010000110001101",
			2147 => "0001001100010100100100",
			2148 => "0010011101101000000100",
			2149 => "0000000010000111011011",
			2150 => "0011111011000000000100",
			2151 => "0000001010000111011011",
			2152 => "0001110110000100001100",
			2153 => "0010010101011100000100",
			2154 => "1111111010000111011011",
			2155 => "0011001100110000000100",
			2156 => "0000000010000111011011",
			2157 => "0000000010000111011011",
			2158 => "0011110000110100000100",
			2159 => "0000001010000111011011",
			2160 => "0000100111111100000100",
			2161 => "0000000010000111011011",
			2162 => "0000101001011100000100",
			2163 => "0000001010000111011011",
			2164 => "0000000010000111011011",
			2165 => "1111111010000111011011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(710, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1428, initial_addr_3'length));
	end generate gen_rom_3;

	gen_rom_4: if SELECT_ROM = 4 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0010110100010000001000",
			10 => "0010111011011100000100",
			11 => "0000000000000001000001",
			12 => "0000000000000001000001",
			13 => "0010110111111100000100",
			14 => "0000000000000001000001",
			15 => "0000000000000001000001",
			16 => "0010100000001000001000",
			17 => "0010101011001100000100",
			18 => "0000000000000001011101",
			19 => "0000000000000001011101",
			20 => "0010100110011000000100",
			21 => "0000000000000001011101",
			22 => "0000000000000001011101",
			23 => "0000010110101000000100",
			24 => "0000000000000001111001",
			25 => "0011011010001000001000",
			26 => "0001111111011100000100",
			27 => "0000000000000001111001",
			28 => "0000000000000001111001",
			29 => "0000000000000001111001",
			30 => "0001011111010000001100",
			31 => "0001110001101000000100",
			32 => "0000000000000010011101",
			33 => "0001011101000100000100",
			34 => "0000000000000010011101",
			35 => "0000000000000010011101",
			36 => "0001110001001000000100",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0010010101011100001100",
			40 => "0011100100001000000100",
			41 => "0000000000000011000001",
			42 => "0000001100011100000100",
			43 => "0000000000000011000001",
			44 => "0000000000000011000001",
			45 => "0001101101111100000100",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0001111000011000001000",
			49 => "0001110001101000000100",
			50 => "0000000000000011100101",
			51 => "0000000000000011100101",
			52 => "0000111010000100000100",
			53 => "0000000000000011100101",
			54 => "0000110010100100000100",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0010110101100100001100",
			58 => "0011001100110000000100",
			59 => "0000000000000100010001",
			60 => "0011001000000000000100",
			61 => "0000000000000100010001",
			62 => "0000000000000100010001",
			63 => "0000010000111100001000",
			64 => "0001110111010000000100",
			65 => "0000000000000100010001",
			66 => "0000000000000100010001",
			67 => "0000000000000100010001",
			68 => "0010100000001000001100",
			69 => "0000000010101100000100",
			70 => "0000000000000100111101",
			71 => "0000000001110000000100",
			72 => "0000000000000100111101",
			73 => "0000000000000100111101",
			74 => "0010100110011000001000",
			75 => "0000000001010100000100",
			76 => "0000000000000100111101",
			77 => "0000000000000100111101",
			78 => "0000000000000100111101",
			79 => "0010110100010000010000",
			80 => "0010111000011000000100",
			81 => "0000000000000101100001",
			82 => "0000010000111100001000",
			83 => "0000011111001100000100",
			84 => "0000000000000101100001",
			85 => "0000000000000101100001",
			86 => "0000000000000101100001",
			87 => "0000000000000101100001",
			88 => "0001001111100100010000",
			89 => "0000101100010000000100",
			90 => "0000000000000110000101",
			91 => "0000101010000100001000",
			92 => "0010001001000100000100",
			93 => "0000000000000110000101",
			94 => "0000000000000110000101",
			95 => "0000000000000110000101",
			96 => "0000000000000110000101",
			97 => "0011001100110000000100",
			98 => "0000000000000110101001",
			99 => "0001011111010000001100",
			100 => "0011011010001000001000",
			101 => "0001111111011100000100",
			102 => "0000000000000110101001",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0001011110010000010000",
			107 => "0000001100011100001000",
			108 => "0010100100111100000100",
			109 => "0000000000000111011101",
			110 => "0000000000000111011101",
			111 => "0010100111101100000100",
			112 => "0000000000000111011101",
			113 => "0000000000000111011101",
			114 => "0001101000010000001000",
			115 => "0000011101111100000100",
			116 => "0000000000000111011101",
			117 => "0000000000000111011101",
			118 => "0000000000000111011101",
			119 => "0001111000011000010000",
			120 => "0011111011000000000100",
			121 => "0000000000001000010001",
			122 => "0011111010000100001000",
			123 => "0010110100010000000100",
			124 => "0000000000001000010001",
			125 => "0000000000001000010001",
			126 => "0000000000001000010001",
			127 => "0011110110111100001000",
			128 => "0011110010000100000100",
			129 => "0000000000001000010001",
			130 => "0000000000001000010001",
			131 => "0000000000001000010001",
			132 => "0010100000001000010000",
			133 => "0010100100110100000100",
			134 => "0000000000001001000101",
			135 => "0000000001010100001000",
			136 => "0010100111101100000100",
			137 => "0000000000001001000101",
			138 => "0000000000001001000101",
			139 => "0000000000001001000101",
			140 => "0000000101000100000100",
			141 => "0000000000001001000101",
			142 => "0010100110011000000100",
			143 => "0000000000001001000101",
			144 => "0000000000001001000101",
			145 => "0000111110110100001100",
			146 => "0010010000111100000100",
			147 => "0000000000001001111001",
			148 => "0000010110101000000100",
			149 => "0000000000001001111001",
			150 => "0000000000001001111001",
			151 => "0000100111010100001100",
			152 => "0010110101110100001000",
			153 => "0000010000111100000100",
			154 => "0000000000001001111001",
			155 => "0000000000001001111001",
			156 => "0000000000001001111001",
			157 => "0000000000001001111001",
			158 => "0010100000001000001100",
			159 => "0011100100001000000100",
			160 => "0000000000001010110101",
			161 => "0001111101100000000100",
			162 => "0000000000001010110101",
			163 => "0000000000001010110101",
			164 => "0000111010000100001000",
			165 => "0001011111010000000100",
			166 => "0000000000001010110101",
			167 => "0000000000001010110101",
			168 => "0001011110000100000100",
			169 => "0000000000001010110101",
			170 => "0001011000100000000100",
			171 => "0000000000001010110101",
			172 => "0000000000001010110101",
			173 => "0001001111100100010100",
			174 => "0000101100010000000100",
			175 => "0000000000001011101001",
			176 => "0010110101110100001100",
			177 => "0010011000010000001000",
			178 => "0000010000111100000100",
			179 => "0000000000001011101001",
			180 => "0000000000001011101001",
			181 => "0000000000001011101001",
			182 => "0000000000001011101001",
			183 => "0010110111111100000100",
			184 => "0000000000001011101001",
			185 => "0000000000001011101001",
			186 => "0011001100110000000100",
			187 => "0000000000001100010101",
			188 => "0001011111010000010000",
			189 => "0011011010001000001100",
			190 => "0011001001110100001000",
			191 => "0000100110101100000100",
			192 => "0000000000001100010101",
			193 => "0000000000001100010101",
			194 => "0000000000001100010101",
			195 => "0000000000001100010101",
			196 => "0000000000001100010101",
			197 => "0010001001101000010100",
			198 => "0011100100001000000100",
			199 => "0000000000001101000001",
			200 => "0000011001011000001100",
			201 => "0010101010100100001000",
			202 => "0001111101100000000100",
			203 => "0000000000001101000001",
			204 => "0000000000001101000001",
			205 => "0000000000001101000001",
			206 => "0000000000001101000001",
			207 => "0000000000001101000001",
			208 => "0011100110100100000100",
			209 => "0000000000001101110101",
			210 => "0001010101001000001000",
			211 => "0011001011000000000100",
			212 => "0000000000001101110101",
			213 => "0000000000001101110101",
			214 => "0011001011011100001100",
			215 => "0001011111010000000100",
			216 => "0000000000001101110101",
			217 => "0011001011000000000100",
			218 => "0000000000001101110101",
			219 => "0000000000001101110101",
			220 => "0000000000001101110101",
			221 => "0001110110000100010000",
			222 => "0011000100000000000100",
			223 => "0000000000001110111001",
			224 => "0011000110000100001000",
			225 => "0000011101101000000100",
			226 => "0000000000001110111001",
			227 => "0000000000001110111001",
			228 => "0000000000001110111001",
			229 => "0000010000111100010000",
			230 => "0001111111011100001100",
			231 => "0011000011011100000100",
			232 => "0000000000001110111001",
			233 => "0000010110101000000100",
			234 => "0000000000001110111001",
			235 => "0000000000001110111001",
			236 => "0000000000001110111001",
			237 => "0000000000001110111001",
			238 => "0000111100010000010000",
			239 => "0011111011000000000100",
			240 => "0000000000010000000101",
			241 => "0011010010011100001000",
			242 => "0011001000000000000100",
			243 => "0000000000010000000101",
			244 => "0000000000010000000101",
			245 => "0000000000010000000101",
			246 => "0011111100000000001000",
			247 => "0001100100110100000100",
			248 => "0000000000010000000101",
			249 => "0000000000010000000101",
			250 => "0011101110111000001100",
			251 => "0000000001010100000100",
			252 => "0000000000010000000101",
			253 => "0011100010000100000100",
			254 => "0000000000010000000101",
			255 => "0000000000010000000101",
			256 => "0000000000010000000101",
			257 => "0000000001010100100000",
			258 => "0011110000011100001100",
			259 => "0000010110101000001000",
			260 => "0011100100001000000100",
			261 => "0000000000010001010001",
			262 => "0000000000010001010001",
			263 => "1111111000010001010001",
			264 => "0001110001101000001100",
			265 => "0010011111000000001000",
			266 => "0010100100111100000100",
			267 => "0000000000010001010001",
			268 => "0000000000010001010001",
			269 => "0000000000010001010001",
			270 => "0001111000011000000100",
			271 => "0000000000010001010001",
			272 => "0000000000010001010001",
			273 => "0001101101111100000100",
			274 => "0000000000010001010001",
			275 => "0000000000010001010001",
			276 => "0000111100010000011100",
			277 => "0010010000111100001100",
			278 => "0011100100001000000100",
			279 => "0000000000010010100101",
			280 => "0000000101000100000100",
			281 => "0000000000010010100101",
			282 => "0000000000010010100101",
			283 => "0000010110101000000100",
			284 => "0000000000010010100101",
			285 => "0011010010011100001000",
			286 => "0011001000000000000100",
			287 => "0000000000010010100101",
			288 => "0000000000010010100101",
			289 => "0000000000010010100101",
			290 => "0010100001010000001100",
			291 => "0001011110101000000100",
			292 => "0000000000010010100101",
			293 => "0000011101111100000100",
			294 => "0000000000010010100101",
			295 => "0000000000010010100101",
			296 => "0000000000010010100101",
			297 => "0011011110101100001100",
			298 => "0010001001111100000100",
			299 => "0000000000010011101001",
			300 => "0011101110101000000100",
			301 => "0000000000010011101001",
			302 => "0000000000010011101001",
			303 => "0000010101011100010100",
			304 => "0011001000011000010000",
			305 => "0001101011001100001100",
			306 => "0011001110001100000100",
			307 => "0000000000010011101001",
			308 => "0011011110101000000100",
			309 => "0000000000010011101001",
			310 => "0000000000010011101001",
			311 => "0000000000010011101001",
			312 => "0000000000010011101001",
			313 => "0000000000010011101001",
			314 => "0010011100011000011000",
			315 => "0011001100110000010000",
			316 => "0001111101100000000100",
			317 => "0000000000010100111101",
			318 => "0011100100001000000100",
			319 => "0000000000010100111101",
			320 => "0000000101000100000100",
			321 => "0000000000010100111101",
			322 => "0000000000010100111101",
			323 => "0010011100011000000100",
			324 => "0000000000010100111101",
			325 => "0000000000010100111101",
			326 => "0000010000111100010000",
			327 => "0001111111011100001100",
			328 => "0001110001111100000100",
			329 => "0000000000010100111101",
			330 => "0001101011001100000100",
			331 => "0000000000010100111101",
			332 => "0000000000010100111101",
			333 => "0000000000010100111101",
			334 => "0000000000010100111101",
			335 => "0001010101001000000100",
			336 => "0000000000010101110001",
			337 => "0001111000011000000100",
			338 => "0000000000010101110001",
			339 => "0001111111011100010000",
			340 => "0000101010000100001100",
			341 => "0010110010001000000100",
			342 => "0000000000010101110001",
			343 => "0010011000010000000100",
			344 => "0000000000010101110001",
			345 => "0000000000010101110001",
			346 => "0000000000010101110001",
			347 => "0000000000010101110001",
			348 => "0001111000011000011100",
			349 => "0011111011000000000100",
			350 => "0000000000010110101101",
			351 => "0000111100010000001100",
			352 => "0001110001101000001000",
			353 => "0011010010011100000100",
			354 => "0000000000010110101101",
			355 => "0000000000010110101101",
			356 => "0000000000010110101101",
			357 => "0011111100000000000100",
			358 => "0000000000010110101101",
			359 => "0011111010000100000100",
			360 => "0000000000010110101101",
			361 => "0000000000010110101101",
			362 => "0000000000010110101101",
			363 => "0001010110100100001100",
			364 => "0011111000000000000100",
			365 => "0000000000011000000001",
			366 => "0011101000011000000100",
			367 => "0000000000011000000001",
			368 => "0000000000011000000001",
			369 => "0010011001100100010100",
			370 => "0011101011000000000100",
			371 => "0000000000011000000001",
			372 => "0011010111111100001100",
			373 => "0010100111110100001000",
			374 => "0010110100001000000100",
			375 => "0000000000011000000001",
			376 => "0000000000011000000001",
			377 => "0000000000011000000001",
			378 => "0000000000011000000001",
			379 => "0011011001011100001000",
			380 => "0000111010000100000100",
			381 => "0000000000011000000001",
			382 => "0000000000011000000001",
			383 => "0000000000011000000001",
			384 => "0000000001010100100100",
			385 => "0001011100100100011000",
			386 => "0001111100101000001100",
			387 => "0000100100001000000100",
			388 => "0000000000011001011101",
			389 => "0011001110001100000100",
			390 => "0000000000011001011101",
			391 => "0000000000011001011101",
			392 => "0011001000000000001000",
			393 => "0000100110010000000100",
			394 => "0000000000011001011101",
			395 => "0000000000011001011101",
			396 => "0000000000011001011101",
			397 => "0001100100110100001000",
			398 => "0011001011000000000100",
			399 => "0000000000011001011101",
			400 => "0000000000011001011101",
			401 => "0000000000011001011101",
			402 => "0011110110001100001000",
			403 => "0010100000001000000100",
			404 => "0000000000011001011101",
			405 => "0000000000011001011101",
			406 => "0000000000011001011101",
			407 => "0001010110100100001100",
			408 => "0011000110000100001000",
			409 => "0001101101011100000100",
			410 => "0000000000011011000001",
			411 => "1111111000011011000001",
			412 => "0000000000011011000001",
			413 => "0000011001011000010000",
			414 => "0011010010110100000100",
			415 => "0000000000011011000001",
			416 => "0001010010011100001000",
			417 => "0000011111001100000100",
			418 => "0000000000011011000001",
			419 => "0000000000011011000001",
			420 => "0000000000011011000001",
			421 => "0011011010001000001100",
			422 => "0001011111010000001000",
			423 => "0010011011001100000100",
			424 => "0000000000011011000001",
			425 => "0000000000011011000001",
			426 => "0000000000011011000001",
			427 => "0000011101111100001000",
			428 => "0010011111000000000100",
			429 => "0000000000011011000001",
			430 => "0000000000011011000001",
			431 => "0000000000011011000001",
			432 => "0010100000001000011000",
			433 => "0010010101011100010000",
			434 => "0000010110101000001100",
			435 => "0000100100001000000100",
			436 => "0000000000011100101101",
			437 => "0000000011101000000100",
			438 => "0000000000011100101101",
			439 => "0000000000011100101101",
			440 => "0000000000011100101101",
			441 => "0000101101000100000100",
			442 => "0000000000011100101101",
			443 => "0000000000011100101101",
			444 => "0000111010000100001100",
			445 => "0011111111010100001000",
			446 => "0000010000111100000100",
			447 => "0000000000011100101101",
			448 => "0000000000011100101101",
			449 => "0000000000011100101101",
			450 => "0011001011000000000100",
			451 => "0000000000011100101101",
			452 => "0001010010011100001100",
			453 => "0000010000111100001000",
			454 => "0001111111011100000100",
			455 => "0000000000011100101101",
			456 => "0000000000011100101101",
			457 => "0000000000011100101101",
			458 => "0000000000011100101101",
			459 => "0000111100010000011100",
			460 => "0010010000111100010000",
			461 => "0000000011101000001100",
			462 => "0000100100001000000100",
			463 => "0000000000011110010001",
			464 => "0001000111001000000100",
			465 => "0000000000011110010001",
			466 => "0000000000011110010001",
			467 => "0000000000011110010001",
			468 => "0011001100110000000100",
			469 => "0000000000011110010001",
			470 => "0000111001100000000100",
			471 => "0000000000011110010001",
			472 => "0000000000011110010001",
			473 => "0010011100011000000100",
			474 => "0000000000011110010001",
			475 => "0000011101111100010000",
			476 => "0011011111010000000100",
			477 => "0000000000011110010001",
			478 => "0010100001010000001000",
			479 => "0011000111001000000100",
			480 => "0000000000011110010001",
			481 => "0000000000011110010001",
			482 => "0000000000011110010001",
			483 => "0000000000011110010001",
			484 => "0011010111111100011100",
			485 => "0000111001001000000100",
			486 => "0000000000011111011101",
			487 => "0010101010100000010100",
			488 => "0010010100111100010000",
			489 => "0011000011011100000100",
			490 => "0000000000011111011101",
			491 => "0011111011000000000100",
			492 => "0000000000011111011101",
			493 => "0011001011000000000100",
			494 => "0000000000011111011101",
			495 => "0000000000011111011101",
			496 => "0000000000011111011101",
			497 => "0000000000011111011101",
			498 => "0010101010100000001000",
			499 => "0000101100000000000100",
			500 => "0000000000011111011101",
			501 => "0000000000011111011101",
			502 => "0000000000011111011101",
			503 => "0001111000000000010100",
			504 => "0000100000110100001100",
			505 => "0000010110101000001000",
			506 => "0011100100001000000100",
			507 => "0000000000100001010001",
			508 => "0000000000100001010001",
			509 => "0000000000100001010001",
			510 => "0011000100011000000100",
			511 => "0000000000100001010001",
			512 => "0000000000100001010001",
			513 => "0011001011000000010000",
			514 => "0010011111000000001100",
			515 => "0001111000011000001000",
			516 => "0001001000001000000100",
			517 => "0000000000100001010001",
			518 => "0000000000100001010001",
			519 => "0000000000100001010001",
			520 => "0000000000100001010001",
			521 => "0000110110111100001000",
			522 => "0001011101000100000100",
			523 => "0000000000100001010001",
			524 => "0000000000100001010001",
			525 => "0001010111100000000100",
			526 => "0000000000100001010001",
			527 => "0000110010100100001000",
			528 => "0000111111010100000100",
			529 => "0000000000100001010001",
			530 => "0000000000100001010001",
			531 => "0000000000100001010001",
			532 => "0001101001011000001100",
			533 => "0000010110101000001000",
			534 => "0011100100001000000100",
			535 => "0000000000100010110101",
			536 => "0000000000100010110101",
			537 => "0000000000100010110101",
			538 => "0001010101001000011000",
			539 => "0010100111101100000100",
			540 => "0000000000100010110101",
			541 => "0000111100010000001000",
			542 => "0010000111110100000100",
			543 => "0000000000100010110101",
			544 => "0000000000100010110101",
			545 => "0010001000100100000100",
			546 => "0000000000100010110101",
			547 => "0010000001010000000100",
			548 => "0000000000100010110101",
			549 => "0000000000100010110101",
			550 => "0011001001110100001100",
			551 => "0000010101011100001000",
			552 => "0000111010000100000100",
			553 => "0000000000100010110101",
			554 => "0000000000100010110101",
			555 => "0000000000100010110101",
			556 => "0000000000100010110101",
			557 => "0010100010101100100000",
			558 => "0011111001001000001000",
			559 => "0011000110000100000100",
			560 => "0000000000100011111001",
			561 => "0000000000100011111001",
			562 => "0000010000111100010100",
			563 => "0001111000011000010000",
			564 => "0011001001110100001100",
			565 => "0011000011011100000100",
			566 => "0000000000100011111001",
			567 => "0010010100111100000100",
			568 => "0000000000100011111001",
			569 => "0000000000100011111001",
			570 => "0000000000100011111001",
			571 => "0000000000100011111001",
			572 => "0000000000100011111001",
			573 => "0000000000100011111001",
			574 => "0010100000001000100100",
			575 => "0000110000110100010100",
			576 => "0010010101011100010000",
			577 => "0011001100110000001100",
			578 => "0011110001111100000100",
			579 => "0000000000100101111101",
			580 => "0011000100000000000100",
			581 => "0000000000100101111101",
			582 => "0000000000100101111101",
			583 => "0000000000100101111101",
			584 => "0000000000100101111101",
			585 => "0001100100110100001100",
			586 => "0011001000000000001000",
			587 => "0010010100111100000100",
			588 => "0000000000100101111101",
			589 => "0000000000100101111101",
			590 => "0000000000100101111101",
			591 => "0000000000100101111101",
			592 => "0000111010000100001000",
			593 => "0011110110111100000100",
			594 => "0000000000100101111101",
			595 => "0000000000100101111101",
			596 => "0010011111000000001100",
			597 => "0010011100011000000100",
			598 => "0000000000100101111101",
			599 => "0001101011001100000100",
			600 => "0000000000100101111101",
			601 => "0000000000100101111101",
			602 => "0001110001001000001000",
			603 => "0000000001010100000100",
			604 => "0000000000100101111101",
			605 => "0000000000100101111101",
			606 => "0000000000100101111101",
			607 => "0001010110100100001100",
			608 => "0011000110000100001000",
			609 => "0001101101011100000100",
			610 => "0000000000100111110001",
			611 => "1111111000100111110001",
			612 => "0000000000100111110001",
			613 => "0000111111010100011100",
			614 => "0000011001011000010000",
			615 => "0000110000110100000100",
			616 => "0000000000100111110001",
			617 => "0011001000000000001000",
			618 => "0011000011011100000100",
			619 => "0000000000100111110001",
			620 => "0000000000100111110001",
			621 => "0000000000100111110001",
			622 => "0011000100011000000100",
			623 => "0000000000100111110001",
			624 => "0011001001110100000100",
			625 => "0000000000100111110001",
			626 => "0000000000100111110001",
			627 => "0011001000000000000100",
			628 => "0000000000100111110001",
			629 => "0000011101111100001100",
			630 => "0011001011011100001000",
			631 => "0000011111001100000100",
			632 => "0000000000100111110001",
			633 => "0000000000100111110001",
			634 => "0000000000100111110001",
			635 => "0000000000100111110001",
			636 => "0011101010001000011100",
			637 => "0000001100011100011000",
			638 => "0010100100111100010000",
			639 => "0001010001101000001100",
			640 => "0000110110100100000100",
			641 => "0000000000101001110101",
			642 => "0001100000111100000100",
			643 => "0000000000101001110101",
			644 => "0000000000101001110101",
			645 => "0000000000101001110101",
			646 => "0011110010001000000100",
			647 => "0000000000101001110101",
			648 => "0000000000101001110101",
			649 => "1111111000101001110101",
			650 => "0000010000111100011100",
			651 => "0000111010000100010100",
			652 => "0001100100110100001100",
			653 => "0011010111111100001000",
			654 => "0010100000001000000100",
			655 => "0000000000101001110101",
			656 => "0000000000101001110101",
			657 => "0000000000101001110101",
			658 => "0000011001011000000100",
			659 => "0000000000101001110101",
			660 => "0000000000101001110101",
			661 => "0001101011001100000100",
			662 => "0000000000101001110101",
			663 => "0000000000101001110101",
			664 => "0001011110010000000100",
			665 => "0000000000101001110101",
			666 => "0010100110011000000100",
			667 => "0000000000101001110101",
			668 => "0000000000101001110101",
			669 => "0000000001010100110000",
			670 => "0001011100100100011100",
			671 => "0011000100011000010000",
			672 => "0001111101100000000100",
			673 => "0000000000101100001001",
			674 => "0011100100001000000100",
			675 => "0000000000101100001001",
			676 => "0010100111101100000100",
			677 => "0000000000101100001001",
			678 => "0000000000101100001001",
			679 => "0001001100000000001000",
			680 => "0010011111000000000100",
			681 => "0000000000101100001001",
			682 => "0000000000101100001001",
			683 => "0000000000101100001001",
			684 => "0000011001011000000100",
			685 => "0000000000101100001001",
			686 => "0010010100111100001100",
			687 => "0011010010011100000100",
			688 => "0000000000101100001001",
			689 => "0011000100011000000100",
			690 => "0000000000101100001001",
			691 => "0000001000101100001001",
			692 => "0000000000101100001001",
			693 => "0010110101100100001000",
			694 => "0000000001110000000100",
			695 => "0000000000101100001001",
			696 => "1111111000101100001001",
			697 => "0010110110110100001000",
			698 => "0010010100111100000100",
			699 => "0000000000101100001001",
			700 => "0000000000101100001001",
			701 => "0001011110010000001000",
			702 => "0011000100011000000100",
			703 => "0000000000101100001001",
			704 => "0000000000101100001001",
			705 => "0000000000101100001001",
			706 => "0000000001010100101000",
			707 => "0000110110111100100100",
			708 => "0001101101111100011000",
			709 => "0001111101100000000100",
			710 => "0000000000101101111101",
			711 => "0010100100111100001100",
			712 => "0001010001101000001000",
			713 => "0011100100001000000100",
			714 => "0000000000101101111101",
			715 => "0000000000101101111101",
			716 => "0000000000101101111101",
			717 => "0011110000110100000100",
			718 => "0000000000101101111101",
			719 => "0000000000101101111101",
			720 => "0001101101111100001000",
			721 => "0010100000001000000100",
			722 => "0000000000101101111101",
			723 => "0000000000101101111101",
			724 => "0000000000101101111101",
			725 => "0000000000101101111101",
			726 => "0000111000001100001000",
			727 => "0000100110101100000100",
			728 => "0000000000101101111101",
			729 => "0000000000101101111101",
			730 => "0000010101011100001000",
			731 => "0010110101110100000100",
			732 => "0000000000101101111101",
			733 => "0000000000101101111101",
			734 => "0000000000101101111101",
			735 => "0000111000001100101100",
			736 => "0010001000100100101000",
			737 => "0011001100110000010000",
			738 => "0000010111100100001100",
			739 => "0000100100001000000100",
			740 => "0000000000101111110001",
			741 => "0000010010001100000100",
			742 => "0000000000101111110001",
			743 => "0000000000101111110001",
			744 => "0000000000101111110001",
			745 => "0000111100010000010000",
			746 => "0000010110101000000100",
			747 => "0000000000101111110001",
			748 => "0011001000000000001000",
			749 => "0011010010011100000100",
			750 => "0000000000101111110001",
			751 => "0000000000101111110001",
			752 => "0000000000101111110001",
			753 => "0000011001011000000100",
			754 => "0000000000101111110001",
			755 => "0000000000101111110001",
			756 => "0000000000101111110001",
			757 => "0001101000010000001100",
			758 => "0011001011000000000100",
			759 => "0000000000101111110001",
			760 => "0000011101111100000100",
			761 => "0000000000101111110001",
			762 => "0000000000101111110001",
			763 => "0000000000101111110001",
			764 => "0010101010100000110000",
			765 => "0011100101110100010100",
			766 => "0011000100000000001000",
			767 => "0001111001110000000100",
			768 => "1111111000110010011101",
			769 => "0000011000110010011101",
			770 => "0000100001101000000100",
			771 => "1111111000110010011101",
			772 => "0010011011111100000100",
			773 => "0000001000110010011101",
			774 => "1111111000110010011101",
			775 => "0010010100111100011000",
			776 => "0000110111010100010100",
			777 => "0001011111010000001100",
			778 => "0011101110101000000100",
			779 => "0000001000110010011101",
			780 => "0000100010000100000100",
			781 => "0000001000110010011101",
			782 => "0000010000110010011101",
			783 => "0000100010000100000100",
			784 => "0000001000110010011101",
			785 => "1111111000110010011101",
			786 => "0000011000110010011101",
			787 => "1111111000110010011101",
			788 => "0010100010101100010100",
			789 => "0000101010000100001100",
			790 => "0000111000001100000100",
			791 => "1111111000110010011101",
			792 => "0001111000011000000100",
			793 => "0000001000110010011101",
			794 => "1111111000110010011101",
			795 => "0000010101011100000100",
			796 => "0000011000110010011101",
			797 => "1111111000110010011101",
			798 => "0010100010101100001000",
			799 => "0011010100101000000100",
			800 => "1111111000110010011101",
			801 => "0000001000110010011101",
			802 => "0011010011000000000100",
			803 => "1111111000110010011101",
			804 => "0010110111111100000100",
			805 => "0000001000110010011101",
			806 => "1111111000110010011101",
			807 => "0001001111100100111000",
			808 => "0000111111010100101000",
			809 => "0010100000001000011100",
			810 => "0010110100001000001100",
			811 => "0000010110101000001000",
			812 => "0011100100001000000100",
			813 => "0000000000110100011001",
			814 => "0000000000110100011001",
			815 => "0000000000110100011001",
			816 => "0000010000111100001100",
			817 => "0011101110101000000100",
			818 => "0000000000110100011001",
			819 => "0011110010000100000100",
			820 => "0000000000110100011001",
			821 => "0000000000110100011001",
			822 => "0000000000110100011001",
			823 => "0000000101000100000100",
			824 => "0000000000110100011001",
			825 => "0001101101111100000100",
			826 => "0000000000110100011001",
			827 => "0000000000110100011001",
			828 => "0010110101110100001100",
			829 => "0010011000010000001000",
			830 => "0000010000111100000100",
			831 => "0000000000110100011001",
			832 => "0000000000110100011001",
			833 => "0000000000110100011001",
			834 => "0000000000110100011001",
			835 => "0011011111101000000100",
			836 => "0000000000110100011001",
			837 => "0000000000110100011001",
			838 => "0001001111100100111000",
			839 => "0001111100101000010000",
			840 => "0001111101100000000100",
			841 => "0000000000110110011101",
			842 => "0000010111100100001000",
			843 => "0011110001111100000100",
			844 => "0000000000110110011101",
			845 => "0000000000110110011101",
			846 => "0000000000110110011101",
			847 => "0000111001100000001000",
			848 => "0011110010000000000100",
			849 => "0000000000110110011101",
			850 => "0000000000110110011101",
			851 => "0001101101111100001000",
			852 => "0011010111111100000100",
			853 => "0000000000110110011101",
			854 => "0000000000110110011101",
			855 => "0000110110111100001100",
			856 => "0010100000001000000100",
			857 => "0000000000110110011101",
			858 => "0001110110100100000100",
			859 => "0000000000110110011101",
			860 => "0000000000110110011101",
			861 => "0010011111000000000100",
			862 => "0000000000110110011101",
			863 => "0000111000001100000100",
			864 => "0000000000110110011101",
			865 => "0000000000110110011101",
			866 => "0011110110001100001000",
			867 => "0001000110111000000100",
			868 => "0000000000110110011101",
			869 => "1111111000110110011101",
			870 => "0000000000110110011101",
			871 => "0000111100000000101000",
			872 => "0001101101111100100000",
			873 => "0011100110100100001000",
			874 => "0001101111001100000100",
			875 => "0000000000111000110001",
			876 => "0000000000111000110001",
			877 => "0011001110001100010000",
			878 => "0010110100001000000100",
			879 => "0000000000111000110001",
			880 => "0011111010011100000100",
			881 => "0000000000111000110001",
			882 => "0001111100101000000100",
			883 => "0000000000111000110001",
			884 => "0000000000111000110001",
			885 => "0010110110100100000100",
			886 => "0000000000111000110001",
			887 => "0000000000111000110001",
			888 => "0010100111101100000100",
			889 => "0000000000111000110001",
			890 => "1111111000111000110001",
			891 => "0010011100011000000100",
			892 => "0000000000111000110001",
			893 => "0010010100111100011000",
			894 => "0001111000011000001100",
			895 => "0001101101111100000100",
			896 => "0000000000111000110001",
			897 => "0000110111011000000100",
			898 => "0000000000111000110001",
			899 => "0000000000111000110001",
			900 => "0010110100010000001000",
			901 => "0010110010001000000100",
			902 => "0000000000111000110001",
			903 => "0000000000111000110001",
			904 => "0000000000111000110001",
			905 => "0000111000100000000100",
			906 => "0000000000111000110001",
			907 => "0000000000111000110001",
			908 => "0011000011011100001000",
			909 => "0001101101011100000100",
			910 => "0000000000111010110101",
			911 => "0000000000111010110101",
			912 => "0000111000100000101100",
			913 => "0010001000100100100000",
			914 => "0010110010001000010100",
			915 => "0000101101000100001100",
			916 => "0011000110000100001000",
			917 => "0001101001011000000100",
			918 => "0000000000111010110101",
			919 => "0000000000111010110101",
			920 => "0000000000111010110101",
			921 => "0000011001011000000100",
			922 => "0000000000111010110101",
			923 => "0000000000111010110101",
			924 => "0000111010000100001000",
			925 => "0000101110110100000100",
			926 => "0000000000111010110101",
			927 => "0000000000111010110101",
			928 => "0000000000111010110101",
			929 => "0000111011111000001000",
			930 => "0000101000100000000100",
			931 => "0000000000111010110101",
			932 => "0000000000111010110101",
			933 => "0000000000111010110101",
			934 => "0001101000010000001100",
			935 => "0011001000000000000100",
			936 => "0000000000111010110101",
			937 => "0000011101111100000100",
			938 => "0000000000111010110101",
			939 => "0000000000111010110101",
			940 => "0000000000111010110101",
			941 => "0001111101100000000100",
			942 => "1111111000111100111001",
			943 => "0000111010000100101000",
			944 => "0010001000100100011100",
			945 => "0000101101000100010000",
			946 => "0010010000111100001000",
			947 => "0011100100001000000100",
			948 => "0000000000111100111001",
			949 => "0000000000111100111001",
			950 => "0010011110010100000100",
			951 => "0000000000111100111001",
			952 => "0000000000111100111001",
			953 => "0010011111000000001000",
			954 => "0001101101111100000100",
			955 => "0000000000111100111001",
			956 => "0000000000111100111001",
			957 => "0000000000111100111001",
			958 => "0011001001110100001000",
			959 => "0011001011000000000100",
			960 => "0000000000111100111001",
			961 => "0000000000111100111001",
			962 => "0000000000111100111001",
			963 => "0001111111011100001000",
			964 => "0010011000010000000100",
			965 => "0000000000111100111001",
			966 => "0000000000111100111001",
			967 => "0001011110010000000100",
			968 => "0000000000111100111001",
			969 => "0001101000010000001000",
			970 => "0010011010100000000100",
			971 => "0000000000111100111001",
			972 => "0000000000111100111001",
			973 => "0000000000111100111001",
			974 => "0000001011010101000000",
			975 => "0010011111000000011000",
			976 => "0001111101100000000100",
			977 => "0000000000111111001101",
			978 => "0011001000000000010000",
			979 => "0001111000011000001100",
			980 => "0011101110101000001000",
			981 => "0011111001110100000100",
			982 => "0000000000111111001101",
			983 => "0000000000111111001101",
			984 => "0000000000111111001101",
			985 => "0000000000111111001101",
			986 => "0000000000111111001101",
			987 => "0010110010001000001100",
			988 => "0000011001011000000100",
			989 => "0000000000111111001101",
			990 => "0010000111110100000100",
			991 => "0000000000111111001101",
			992 => "0000000000111111001101",
			993 => "0010110100010000010000",
			994 => "0010101010100000001000",
			995 => "0001100100110100000100",
			996 => "0000000000111111001101",
			997 => "0000000000111111001101",
			998 => "0000100111011000000100",
			999 => "0000000000111111001101",
			1000 => "0000000000111111001101",
			1001 => "0001101010011000000100",
			1002 => "0000000000111111001101",
			1003 => "0010101010100100000100",
			1004 => "0000000000111111001101",
			1005 => "0000000000111111001101",
			1006 => "0011110110001100000100",
			1007 => "1111111000111111001101",
			1008 => "0001101000010000000100",
			1009 => "0000000000111111001101",
			1010 => "0000000000111111001101",
			1011 => "0010001000100100101100",
			1012 => "0011110001001000011100",
			1013 => "0011110010001000011000",
			1014 => "0011001000111100001000",
			1015 => "0011100100001000000100",
			1016 => "1100111001000010001001",
			1017 => "1101100001000010001001",
			1018 => "0011111011011100001100",
			1019 => "0011101011000000000100",
			1020 => "1100111001000010001001",
			1021 => "0010010001000100000100",
			1022 => "1101011001000010001001",
			1023 => "1100111001000010001001",
			1024 => "1101000001000010001001",
			1025 => "1101010001000010001001",
			1026 => "0010011111000000001000",
			1027 => "0000100111100000000100",
			1028 => "1110010001000010001001",
			1029 => "1111000001000010001001",
			1030 => "0011010100101000000100",
			1031 => "1100111001000010001001",
			1032 => "1110010001000010001001",
			1033 => "0010001000100100001100",
			1034 => "0010011111000000000100",
			1035 => "1110101001000010001001",
			1036 => "0011111100000000000100",
			1037 => "1100111001000010001001",
			1038 => "1101011001000010001001",
			1039 => "0010001001000100010100",
			1040 => "0000101010000100010000",
			1041 => "0010011111000000001000",
			1042 => "0000100111100000000100",
			1043 => "1100111001000010001001",
			1044 => "1101100001000010001001",
			1045 => "0000110000010000000100",
			1046 => "1100111001000010001001",
			1047 => "1101001001000010001001",
			1048 => "1101110001000010001001",
			1049 => "0010100010101100010000",
			1050 => "0001001101101100001000",
			1051 => "0010101010100100000100",
			1052 => "1101000001000010001001",
			1053 => "1100111001000010001001",
			1054 => "0010001010110000000100",
			1055 => "1101010001000010001001",
			1056 => "1100111001000010001001",
			1057 => "1100111001000010001001",
			1058 => "0000001011010101001000",
			1059 => "0001100100110100101000",
			1060 => "0011101110101000010100",
			1061 => "0001100001000100010000",
			1062 => "0011000110000100001100",
			1063 => "0011100100001000000100",
			1064 => "0000000001000100110101",
			1065 => "0010010101011100000100",
			1066 => "0000001001000100110101",
			1067 => "0000000001000100110101",
			1068 => "0000000001000100110101",
			1069 => "1111111001000100110101",
			1070 => "0010010100111100010000",
			1071 => "0001111111011100001100",
			1072 => "0010011111000000000100",
			1073 => "0000001001000100110101",
			1074 => "0001111000011000000100",
			1075 => "0000000001000100110101",
			1076 => "0000001001000100110101",
			1077 => "0000000001000100110101",
			1078 => "0000000001000100110101",
			1079 => "0000111000001100010100",
			1080 => "0000100010000100001100",
			1081 => "0001010001000000001000",
			1082 => "0010001000100100000100",
			1083 => "0000000001000100110101",
			1084 => "1111111001000100110101",
			1085 => "0000000001000100110101",
			1086 => "0000011001011000000100",
			1087 => "0000000001000100110101",
			1088 => "1111111001000100110101",
			1089 => "0000010101011100001000",
			1090 => "0011001001110100000100",
			1091 => "0000001001000100110101",
			1092 => "0000000001000100110101",
			1093 => "0000000001000100110101",
			1094 => "0011110110001100000100",
			1095 => "1111111001000100110101",
			1096 => "0001100101010000001000",
			1097 => "0000010100110100000100",
			1098 => "0000001001000100110101",
			1099 => "0000000001000100110101",
			1100 => "1111111001000100110101",
			1101 => "0001001111100101000100",
			1102 => "0010010101011100010000",
			1103 => "0000000011101000001100",
			1104 => "0011110001111100000100",
			1105 => "0000000001000111010001",
			1106 => "0000010111100100000100",
			1107 => "0000000001000111010001",
			1108 => "0000000001000111010001",
			1109 => "0000000001000111010001",
			1110 => "0000111001100000010100",
			1111 => "0000011101011100001000",
			1112 => "0010011110010100000100",
			1113 => "0000000001000111010001",
			1114 => "0000000001000111010001",
			1115 => "0010011101011000000100",
			1116 => "0000000001000111010001",
			1117 => "0000101110010000000100",
			1118 => "0000000001000111010001",
			1119 => "0000000001000111010001",
			1120 => "0001101101111100001000",
			1121 => "0011010111111100000100",
			1122 => "0000000001000111010001",
			1123 => "0000000001000111010001",
			1124 => "0000110110111100001100",
			1125 => "0010100000001000000100",
			1126 => "0000000001000111010001",
			1127 => "0011001010111000000100",
			1128 => "0000000001000111010001",
			1129 => "0000000001000111010001",
			1130 => "0010110101110100001000",
			1131 => "0001010111100000000100",
			1132 => "0000000001000111010001",
			1133 => "0000000001000111010001",
			1134 => "0000000001000111010001",
			1135 => "0011110110001100001000",
			1136 => "0001000110111000000100",
			1137 => "0000000001000111010001",
			1138 => "0000000001000111010001",
			1139 => "0000000001000111010001",
			1140 => "0000001101010001000000",
			1141 => "0011000001111100011100",
			1142 => "0001100001000100010100",
			1143 => "0000010111100100010000",
			1144 => "0011100100001000000100",
			1145 => "0000000001001001010101",
			1146 => "0011001100110000001000",
			1147 => "0001111101100000000100",
			1148 => "0000000001001001010101",
			1149 => "0000000001001001010101",
			1150 => "0000000001001001010101",
			1151 => "0000000001001001010101",
			1152 => "0001111000000000000100",
			1153 => "0000000001001001010101",
			1154 => "0000000001001001010101",
			1155 => "0000011001011000001000",
			1156 => "0010011100011000000100",
			1157 => "0000000001001001010101",
			1158 => "0000000001001001010101",
			1159 => "0000111111010100001100",
			1160 => "0000011001011000001000",
			1161 => "0001011101000100000100",
			1162 => "0000000001001001010101",
			1163 => "0000000001001001010101",
			1164 => "0000000001001001010101",
			1165 => "0000010000111100001000",
			1166 => "0001011111010000000100",
			1167 => "0000000001001001010101",
			1168 => "0000000001001001010101",
			1169 => "0001011100010000000100",
			1170 => "0000000001001001010101",
			1171 => "0000000001001001010101",
			1172 => "0000000001001001010101",
			1173 => "0001111101100000000100",
			1174 => "1111111001001011101001",
			1175 => "0000111010000100101000",
			1176 => "0000000101000100011000",
			1177 => "0000101101000100010000",
			1178 => "0010010000111100001000",
			1179 => "0011100100001000000100",
			1180 => "0000000001001011101001",
			1181 => "0000000001001011101001",
			1182 => "0010011110010100000100",
			1183 => "0000000001001011101001",
			1184 => "0000000001001011101001",
			1185 => "0001101101111100000100",
			1186 => "0000000001001011101001",
			1187 => "0000000001001011101001",
			1188 => "0010001000100100000100",
			1189 => "0000000001001011101001",
			1190 => "0010110110110100000100",
			1191 => "0000000001001011101001",
			1192 => "0000100111011000000100",
			1193 => "0000000001001011101001",
			1194 => "0000000001001011101001",
			1195 => "0001111111011100010000",
			1196 => "0010011000010000001100",
			1197 => "0000010000111100001000",
			1198 => "0001100100110100000100",
			1199 => "0000000001001011101001",
			1200 => "0000001001001011101001",
			1201 => "0000000001001011101001",
			1202 => "0000000001001011101001",
			1203 => "0011010110010000000100",
			1204 => "0000000001001011101001",
			1205 => "0001101000010000001000",
			1206 => "0000011101111100000100",
			1207 => "0000000001001011101001",
			1208 => "0000000001001011101001",
			1209 => "0000000001001011101001",
			1210 => "0000001011010101010100",
			1211 => "0010011111000000100100",
			1212 => "0000001010100100010000",
			1213 => "0010010000111100001100",
			1214 => "0011110001111100000100",
			1215 => "0000000001001110100101",
			1216 => "0001111101100000000100",
			1217 => "0000000001001110100101",
			1218 => "0000001001001110100101",
			1219 => "0000000001001110100101",
			1220 => "0000110000110100001000",
			1221 => "0010010101011100000100",
			1222 => "0000000001001110100101",
			1223 => "0000000001001110100101",
			1224 => "0011001000000000001000",
			1225 => "0001111000011000000100",
			1226 => "0000001001001110100101",
			1227 => "0000000001001110100101",
			1228 => "0000000001001110100101",
			1229 => "0000110111010100011000",
			1230 => "0000000101000100001100",
			1231 => "0011010101110000001000",
			1232 => "0011000100011000000100",
			1233 => "0000000001001110100101",
			1234 => "0000000001001110100101",
			1235 => "0000000001001110100101",
			1236 => "0001111111011100001000",
			1237 => "0011001011000000000100",
			1238 => "0000000001001110100101",
			1239 => "1111111001001110100101",
			1240 => "0000000001001110100101",
			1241 => "0011001001110100001100",
			1242 => "0010110010001000000100",
			1243 => "0000000001001110100101",
			1244 => "0000010101011100000100",
			1245 => "0000000001001110100101",
			1246 => "0000000001001110100101",
			1247 => "0001101010011000000100",
			1248 => "0000000001001110100101",
			1249 => "0011011110010000000100",
			1250 => "0000000001001110100101",
			1251 => "0000000001001110100101",
			1252 => "0011110110001100000100",
			1253 => "1111111001001110100101",
			1254 => "0001101000010000000100",
			1255 => "0000000001001110100101",
			1256 => "0000000001001110100101",
			1257 => "0010001000100100110100",
			1258 => "0011100101110100011100",
			1259 => "0001101101011100001000",
			1260 => "0000111010111100000100",
			1261 => "1111111001010001110001",
			1262 => "0000011001010001110001",
			1263 => "0011000100000000000100",
			1264 => "0000000001010001110001",
			1265 => "0010110100001000000100",
			1266 => "1111111001010001110001",
			1267 => "0010010001000100001000",
			1268 => "0011001100110000000100",
			1269 => "0000010001010001110001",
			1270 => "0000000001010001110001",
			1271 => "1111111001010001110001",
			1272 => "0010010100111100010100",
			1273 => "0000110111010100010000",
			1274 => "0011100010000100001100",
			1275 => "0001110100001000000100",
			1276 => "0000010001010001110001",
			1277 => "0011111111010000000100",
			1278 => "0000000001010001110001",
			1279 => "0000010001010001110001",
			1280 => "0000001001010001110001",
			1281 => "0000100001010001110001",
			1282 => "1111111001010001110001",
			1283 => "0010100010101100100000",
			1284 => "0000111000100000011100",
			1285 => "0000101010000100010100",
			1286 => "0000111000001100001100",
			1287 => "0010101010100000001000",
			1288 => "0011110111011000000100",
			1289 => "1111111001010001110001",
			1290 => "0000001001010001110001",
			1291 => "1111111001010001110001",
			1292 => "0011100111011000000100",
			1293 => "0000010001010001110001",
			1294 => "1111111001010001110001",
			1295 => "0000100111010100000100",
			1296 => "0000010001010001110001",
			1297 => "1111111001010001110001",
			1298 => "0000101001010001110001",
			1299 => "0010100010101100001000",
			1300 => "0011010100101000000100",
			1301 => "1111111001010001110001",
			1302 => "0000001001010001110001",
			1303 => "0011010011000000000100",
			1304 => "1111111001010001110001",
			1305 => "0010110111111100000100",
			1306 => "0000010001010001110001",
			1307 => "1111111001010001110001",
			1308 => "0000001011010100111100",
			1309 => "0011000001101000111000",
			1310 => "0010000111110100011100",
			1311 => "0000101100100100010100",
			1312 => "0000010111100100001100",
			1313 => "0011101011000000001000",
			1314 => "0011000110000100000100",
			1315 => "0000000001010100001101",
			1316 => "0000000001010100001101",
			1317 => "0000001001010100001101",
			1318 => "0011001100110000000100",
			1319 => "0000000001010100001101",
			1320 => "1111111001010100001101",
			1321 => "0010011001100100000100",
			1322 => "0000001001010100001101",
			1323 => "0000000001010100001101",
			1324 => "0000111100010000001000",
			1325 => "0010100111101100000100",
			1326 => "0000000001010100001101",
			1327 => "1111111001010100001101",
			1328 => "0010100000001000000100",
			1329 => "0000001001010100001101",
			1330 => "0000111010000100001000",
			1331 => "0010110010001000000100",
			1332 => "0000000001010100001101",
			1333 => "1111111001010100001101",
			1334 => "0000000001010100000100",
			1335 => "0000001001010100001101",
			1336 => "0000000001010100001101",
			1337 => "0000001001010100001101",
			1338 => "0010110101100100000100",
			1339 => "1111111001010100001101",
			1340 => "0010111011011100001000",
			1341 => "0011100110111100000100",
			1342 => "0000001001010100001101",
			1343 => "0000000001010100001101",
			1344 => "0001011111100100000100",
			1345 => "1111111001010100001101",
			1346 => "0000000001010100001101",
			1347 => "0010010100111101000100",
			1348 => "0011101010001000100000",
			1349 => "0000001100011100011000",
			1350 => "0001110000001100010000",
			1351 => "0011000011011100000100",
			1352 => "0000000001010110100001",
			1353 => "0011011000011000000100",
			1354 => "0000000001010110100001",
			1355 => "0011000110000100000100",
			1356 => "0000000001010110100001",
			1357 => "0000000001010110100001",
			1358 => "0011010000110100000100",
			1359 => "0000000001010110100001",
			1360 => "0000000001010110100001",
			1361 => "0010000011101000000100",
			1362 => "0000000001010110100001",
			1363 => "0000000001010110100001",
			1364 => "0001111111011100100000",
			1365 => "0001111000011000011000",
			1366 => "0010110110110100001100",
			1367 => "0001110001101000001000",
			1368 => "0000000010101000000100",
			1369 => "0000000001010110100001",
			1370 => "0000000001010110100001",
			1371 => "0000000001010110100001",
			1372 => "0000000101000100000100",
			1373 => "0000000001010110100001",
			1374 => "0011001011000000000100",
			1375 => "0000000001010110100001",
			1376 => "0000000001010110100001",
			1377 => "0000111100000000000100",
			1378 => "0000000001010110100001",
			1379 => "0000000001010110100001",
			1380 => "0000000001010110100001",
			1381 => "0000010000111100000100",
			1382 => "0000000001010110100001",
			1383 => "0000000001010110100001",
			1384 => "0000000011101000001100",
			1385 => "0000010111100100001000",
			1386 => "0011100100001000000100",
			1387 => "0000000001011000111101",
			1388 => "0000000001011000111101",
			1389 => "0000000001011000111101",
			1390 => "0001111000000000001100",
			1391 => "0001100001000100000100",
			1392 => "0000000001011000111101",
			1393 => "0011001010111100000100",
			1394 => "1111111001011000111101",
			1395 => "0000000001011000111101",
			1396 => "0000011001011000001100",
			1397 => "0001101011001100001000",
			1398 => "0011101110101000000100",
			1399 => "0000000001011000111101",
			1400 => "0000000001011000111101",
			1401 => "0000000001011000111101",
			1402 => "0000111100000000010000",
			1403 => "0001101101111100000100",
			1404 => "0000000001011000111101",
			1405 => "0001111001001000000100",
			1406 => "0000000001011000111101",
			1407 => "0011000100011000000100",
			1408 => "0000000001011000111101",
			1409 => "0000000001011000111101",
			1410 => "0011001000000000010000",
			1411 => "0001100100110100001000",
			1412 => "0010110101100100000100",
			1413 => "0000000001011000111101",
			1414 => "0000000001011000111101",
			1415 => "0011011010001000000100",
			1416 => "0000000001011000111101",
			1417 => "0000000001011000111101",
			1418 => "0000101110110100000100",
			1419 => "0000000001011000111101",
			1420 => "0001000000010000000100",
			1421 => "0000000001011000111101",
			1422 => "0000000001011000111101",
			1423 => "0000001101010001000000",
			1424 => "0001111000000000010100",
			1425 => "0000000110011100010000",
			1426 => "0011111011000000000100",
			1427 => "0000000001011011000001",
			1428 => "0000010111100100001000",
			1429 => "0011000011011100000100",
			1430 => "0000000001011011000001",
			1431 => "0000000001011011000001",
			1432 => "0000000001011011000001",
			1433 => "0000000001011011000001",
			1434 => "0000011001011000001100",
			1435 => "0001111111011100001000",
			1436 => "0011010111111100000100",
			1437 => "0000001001011011000001",
			1438 => "0000000001011011000001",
			1439 => "0000000001011011000001",
			1440 => "0011010100101000000100",
			1441 => "0000000001011011000001",
			1442 => "0001111000011000010000",
			1443 => "0011001000000000001000",
			1444 => "0010110100010000000100",
			1445 => "0000000001011011000001",
			1446 => "0000000001011011000001",
			1447 => "0001110001101000000100",
			1448 => "0000000001011011000001",
			1449 => "0000000001011011000001",
			1450 => "0010110010001000000100",
			1451 => "0000000001011011000001",
			1452 => "0000011101111100000100",
			1453 => "0000000001011011000001",
			1454 => "0000000001011011000001",
			1455 => "1111111001011011000001",
			1456 => "0001111101100000000100",
			1457 => "1111111001011101000101",
			1458 => "0010100111101100010000",
			1459 => "0000101101000100001100",
			1460 => "0010111110110000001000",
			1461 => "0000100100001000000100",
			1462 => "0000000001011101000101",
			1463 => "0000001001011101000101",
			1464 => "1111111001011101000101",
			1465 => "0000001001011101000101",
			1466 => "0001011110101000001100",
			1467 => "0010000111110100000100",
			1468 => "0000000001011101000101",
			1469 => "0010111011011100000100",
			1470 => "1111111001011101000101",
			1471 => "0000000001011101000101",
			1472 => "0010011100011000000100",
			1473 => "1111111001011101000101",
			1474 => "0001111000011000010000",
			1475 => "0010011111000000001000",
			1476 => "0000111111010100000100",
			1477 => "0000000001011101000101",
			1478 => "0000001001011101000101",
			1479 => "0011011010001000000100",
			1480 => "0000000001011101000101",
			1481 => "0000000001011101000101",
			1482 => "0000111000100000001000",
			1483 => "0010001000100100000100",
			1484 => "0000000001011101000101",
			1485 => "1111111001011101000101",
			1486 => "0010011010100000000100",
			1487 => "0000001001011101000101",
			1488 => "0000000001011101000101",
			1489 => "0010101010100101100000",
			1490 => "0010001000100100110000",
			1491 => "0000101101000100011100",
			1492 => "0000010111100100010000",
			1493 => "0011101010111000001000",
			1494 => "0001101111001100000100",
			1495 => "0000001001100000110001",
			1496 => "1111111001100000110001",
			1497 => "0011111011000000000100",
			1498 => "0000110001100000110001",
			1499 => "0000001001100000110001",
			1500 => "0010000000001000000100",
			1501 => "1111111001100000110001",
			1502 => "0001100001000100000100",
			1503 => "0000000001100000110001",
			1504 => "1111111001100000110001",
			1505 => "0000010000111100010000",
			1506 => "0001111000011000001100",
			1507 => "0010100000001000000100",
			1508 => "0000001001100000110001",
			1509 => "0011100110010000000100",
			1510 => "0000000001100000110001",
			1511 => "0000001001100000110001",
			1512 => "0000000001100000110001",
			1513 => "1111111001100000110001",
			1514 => "0000111010000100100000",
			1515 => "0010100000001000001000",
			1516 => "0000100110010000000100",
			1517 => "1111111001100000110001",
			1518 => "0000001001100000110001",
			1519 => "0001101101111100001000",
			1520 => "0000011111001100000100",
			1521 => "0000000001100000110001",
			1522 => "0000001001100000110001",
			1523 => "0011111100010000001000",
			1524 => "0001010001000000000100",
			1525 => "1111111001100000110001",
			1526 => "0000001001100000110001",
			1527 => "0001110001101000000100",
			1528 => "0000000001100000110001",
			1529 => "1111111001100000110001",
			1530 => "0001111111011100001100",
			1531 => "0010010100111100001000",
			1532 => "0000110111010100000100",
			1533 => "0000001001100000110001",
			1534 => "0000010001100000110001",
			1535 => "0000000001100000110001",
			1536 => "1111111001100000110001",
			1537 => "0010100111110100001100",
			1538 => "0000100110101100000100",
			1539 => "1111111001100000110001",
			1540 => "0000011110010100000100",
			1541 => "0000010001100000110001",
			1542 => "0000000001100000110001",
			1543 => "0001011111100100000100",
			1544 => "1111111001100000110001",
			1545 => "0011111011100100000100",
			1546 => "0000001001100000110001",
			1547 => "1111111001100000110001",
			1548 => "0000001001101001001100",
			1549 => "0011101110101000011100",
			1550 => "0001100001000100011000",
			1551 => "0000111001001000000100",
			1552 => "0000000001100011111101",
			1553 => "0011000110000100010000",
			1554 => "0011001100110000001000",
			1555 => "0001000111010000000100",
			1556 => "0000000001100011111101",
			1557 => "0000000001100011111101",
			1558 => "0000010111100100000100",
			1559 => "0000001001100011111101",
			1560 => "0000000001100011111101",
			1561 => "0000000001100011111101",
			1562 => "1111111001100011111101",
			1563 => "0001101101111100001000",
			1564 => "0011001000000000000100",
			1565 => "0000001001100011111101",
			1566 => "0000000001100011111101",
			1567 => "0000111100000000001000",
			1568 => "0011000100011000000100",
			1569 => "0000000001100011111101",
			1570 => "1111111001100011111101",
			1571 => "0011001000000000010000",
			1572 => "0001100100110100001000",
			1573 => "0010010100111100000100",
			1574 => "0000001001100011111101",
			1575 => "0000000001100011111101",
			1576 => "0000110111010100000100",
			1577 => "0000000001100011111101",
			1578 => "0000001001100011111101",
			1579 => "0011011010001000001000",
			1580 => "0000000101000100000100",
			1581 => "0000001001100011111101",
			1582 => "1111111001100011111101",
			1583 => "0011001001001000000100",
			1584 => "0000001001100011111101",
			1585 => "0000000001100011111101",
			1586 => "0000100010110000010000",
			1587 => "0010000110011100001100",
			1588 => "0011011111010000000100",
			1589 => "1111111001100011111101",
			1590 => "0011100110111100000100",
			1591 => "0000000001100011111101",
			1592 => "0000000001100011111101",
			1593 => "1111111001100011111101",
			1594 => "0010100001010000001000",
			1595 => "0001100101010000000100",
			1596 => "0000001001100011111101",
			1597 => "0000000001100011111101",
			1598 => "1111111001100011111101",
			1599 => "0010100010101101000100",
			1600 => "0000010000111101000000",
			1601 => "0011101110101000100000",
			1602 => "0000000110011000011100",
			1603 => "0011001100110000010000",
			1604 => "0011111011000000001000",
			1605 => "0001101111001100000100",
			1606 => "0000001001100110110001",
			1607 => "1111111001100110110001",
			1608 => "0000010111100100000100",
			1609 => "0000010001100110110001",
			1610 => "0000001001100110110001",
			1611 => "0000010111100100001000",
			1612 => "0011000110000100000100",
			1613 => "0000000001100110110001",
			1614 => "0000000001100110110001",
			1615 => "1111111001100110110001",
			1616 => "1111111001100110110001",
			1617 => "0000111000001100011000",
			1618 => "0001101101111100001100",
			1619 => "0010110010001000000100",
			1620 => "0000001001100110110001",
			1621 => "0011001011000000000100",
			1622 => "0000001001100110110001",
			1623 => "0000000001100110110001",
			1624 => "0000111100010000000100",
			1625 => "1111110001100110110001",
			1626 => "0000011001011000000100",
			1627 => "0000001001100110110001",
			1628 => "0000000001100110110001",
			1629 => "0010110101110100000100",
			1630 => "0000010001100110110001",
			1631 => "0000001001100110110001",
			1632 => "1111111001100110110001",
			1633 => "0010100011101000001100",
			1634 => "0001001111101000000100",
			1635 => "1111111001100110110001",
			1636 => "0010000110011100000100",
			1637 => "0000010001100110110001",
			1638 => "0000000001100110110001",
			1639 => "0001011111100100000100",
			1640 => "1111111001100110110001",
			1641 => "0010110111111100000100",
			1642 => "0000001001100110110001",
			1643 => "1111111001100110110001",
			1644 => "0000001100000101011000",
			1645 => "0010000111110100011100",
			1646 => "0000101101000100010100",
			1647 => "0001111100101000010000",
			1648 => "0011100100001000000100",
			1649 => "0000000001101010010101",
			1650 => "0010010000111100000100",
			1651 => "0000001001101010010101",
			1652 => "0011010100000100000100",
			1653 => "1111111001101010010101",
			1654 => "0000001001101010010101",
			1655 => "1111111001101010010101",
			1656 => "0001101101111100000100",
			1657 => "0000001001101010010101",
			1658 => "0000000001101010010101",
			1659 => "0000111110110100001100",
			1660 => "0010110101100100001000",
			1661 => "0000100011001000000100",
			1662 => "1111111001101010010101",
			1663 => "0000000001101010010101",
			1664 => "1111110001101010010101",
			1665 => "0000101110110100010000",
			1666 => "0010100000001000001000",
			1667 => "0010010100111100000100",
			1668 => "0000001001101010010101",
			1669 => "0000000001101010010101",
			1670 => "0000110110111100000100",
			1671 => "1111111001101010010101",
			1672 => "0000000001101010010101",
			1673 => "0000111010000100010000",
			1674 => "0010110110110100001000",
			1675 => "0010011111000000000100",
			1676 => "0000000001101010010101",
			1677 => "0000000001101010010101",
			1678 => "0000000001010100000100",
			1679 => "1111111001101010010101",
			1680 => "0000000001101010010101",
			1681 => "0011011001011100001000",
			1682 => "0000000001110000000100",
			1683 => "0000001001101010010101",
			1684 => "0000000001101010010101",
			1685 => "0000100110111100000100",
			1686 => "1111111001101010010101",
			1687 => "0000001001101010010101",
			1688 => "0000100010110000010000",
			1689 => "0010100011101000001100",
			1690 => "0001001101101100000100",
			1691 => "1111111001101010010101",
			1692 => "0001011101000100000100",
			1693 => "0000000001101010010101",
			1694 => "0000000001101010010101",
			1695 => "1111111001101010010101",
			1696 => "0001101000010000000100",
			1697 => "0000001001101010010101",
			1698 => "0010001001101000000100",
			1699 => "0000000001101010010101",
			1700 => "1111111001101010010101",
			1701 => "0000001100000101010000",
			1702 => "0010000111110100011000",
			1703 => "0011100100001000000100",
			1704 => "0000000001101101100001",
			1705 => "0000010000111100010000",
			1706 => "0000010110101000000100",
			1707 => "0000001001101101100001",
			1708 => "0010110100001000000100",
			1709 => "1111111001101101100001",
			1710 => "0011110010001000000100",
			1711 => "0000000001101101100001",
			1712 => "0000001001101101100001",
			1713 => "0000000001101101100001",
			1714 => "0000111100010000001000",
			1715 => "0001001100000000000100",
			1716 => "1111111001101101100001",
			1717 => "0000000001101101100001",
			1718 => "0011001000000000100000",
			1719 => "0011110111011000010000",
			1720 => "0010001000100100001000",
			1721 => "0000111100000000000100",
			1722 => "0000000001101101100001",
			1723 => "0000001001101101100001",
			1724 => "0011100010000100000100",
			1725 => "0000000001101101100001",
			1726 => "1111111001101101100001",
			1727 => "0000000001110000001000",
			1728 => "0010110010001000000100",
			1729 => "0000000001101101100001",
			1730 => "0000001001101101100001",
			1731 => "0011001011000000000100",
			1732 => "0000000001101101100001",
			1733 => "0000000001101101100001",
			1734 => "0000000101000100000100",
			1735 => "0000001001101101100001",
			1736 => "0001011001010000000100",
			1737 => "1111111001101101100001",
			1738 => "0011001001001000000100",
			1739 => "0000001001101101100001",
			1740 => "0000000001101101100001",
			1741 => "0000011111001100000100",
			1742 => "1111111001101101100001",
			1743 => "0010010100111100001100",
			1744 => "0011011111010000000100",
			1745 => "1111111001101101100001",
			1746 => "0000110010010100000100",
			1747 => "0000001001101101100001",
			1748 => "0000000001101101100001",
			1749 => "0001010000010000000100",
			1750 => "1111111001101101100001",
			1751 => "0000001001101101100001",
			1752 => "0000001100000101011000",
			1753 => "0011001000000000110100",
			1754 => "0011111100100100010100",
			1755 => "0001100001000100010000",
			1756 => "0011000110000100001100",
			1757 => "0011100100001000000100",
			1758 => "0000000001110001000101",
			1759 => "0010010000111100000100",
			1760 => "0000001001110001000101",
			1761 => "0000000001110001000101",
			1762 => "0000000001110001000101",
			1763 => "1111111001110001000101",
			1764 => "0010011111000000000100",
			1765 => "0000001001110001000101",
			1766 => "0001111000011000010000",
			1767 => "0011001011000000001000",
			1768 => "0001011110101000000100",
			1769 => "0000000001110001000101",
			1770 => "0000001001110001000101",
			1771 => "0010100000001000000100",
			1772 => "0000000001110001000101",
			1773 => "1111111001110001000101",
			1774 => "0001111000011000001000",
			1775 => "0010010100111100000100",
			1776 => "0000001001110001000101",
			1777 => "0000000001110001000101",
			1778 => "0000000001110001000101",
			1779 => "0011101010001000000100",
			1780 => "1111111001110001000101",
			1781 => "0011111100010000001000",
			1782 => "0010100000001000000100",
			1783 => "0000001001110001000101",
			1784 => "0000000001110001000101",
			1785 => "0011001000000000001000",
			1786 => "0010001000100100000100",
			1787 => "0000001001110001000101",
			1788 => "0000000001110001000101",
			1789 => "0010001000010100001000",
			1790 => "0011001001110100000100",
			1791 => "1111111001110001000101",
			1792 => "0000000001110001000101",
			1793 => "0011001001110100000100",
			1794 => "0000001001110001000101",
			1795 => "0000000001110001000101",
			1796 => "0011110110001100010000",
			1797 => "0010100011101000001100",
			1798 => "0001001101101100000100",
			1799 => "1111111001110001000101",
			1800 => "0001011101000100000100",
			1801 => "0000000001110001000101",
			1802 => "0000000001110001000101",
			1803 => "1111111001110001000101",
			1804 => "0001100101010000001000",
			1805 => "0000001101010000000100",
			1806 => "0000000001110001000101",
			1807 => "0000001001110001000101",
			1808 => "1111111001110001000101",
			1809 => "0001011110110000000100",
			1810 => "1111111001110011110001",
			1811 => "0000000001010100110100",
			1812 => "0000110110111100101100",
			1813 => "0011000100011000011000",
			1814 => "0011111100100100001100",
			1815 => "0001100001000100001000",
			1816 => "0010110100001000000100",
			1817 => "0000000001110011110001",
			1818 => "0000000001110011110001",
			1819 => "1111111001110011110001",
			1820 => "0001100100110100001000",
			1821 => "0010010100111100000100",
			1822 => "0000001001110011110001",
			1823 => "0000000001110011110001",
			1824 => "0000000001110011110001",
			1825 => "0001101101111100000100",
			1826 => "0000000001110011110001",
			1827 => "0001011100100100001000",
			1828 => "0010011001100100000100",
			1829 => "0000000001110011110001",
			1830 => "1111111001110011110001",
			1831 => "0000000101000100000100",
			1832 => "0000000001110011110001",
			1833 => "1111111001110011110001",
			1834 => "0001011110000100000100",
			1835 => "0000000001110011110001",
			1836 => "0000001001110011110001",
			1837 => "0000111000001100001000",
			1838 => "0011110000010000000100",
			1839 => "1111111001110011110001",
			1840 => "0000000001110011110001",
			1841 => "0001101011001100001100",
			1842 => "0010011000010000001000",
			1843 => "0001010010011100000100",
			1844 => "0000001001110011110001",
			1845 => "0000000001110011110001",
			1846 => "0000000001110011110001",
			1847 => "0011010011000000000100",
			1848 => "1111111001110011110001",
			1849 => "0000001010111000000100",
			1850 => "0000000001110011110001",
			1851 => "0000000001110011110001",
			1852 => "0001111101100000000100",
			1853 => "1111111001110110110101",
			1854 => "0001111000011000111000",
			1855 => "0010100000001000100100",
			1856 => "0000111100010000011100",
			1857 => "0010000111110100010000",
			1858 => "0000101101000100001000",
			1859 => "0010010000111100000100",
			1860 => "0000000001110110110101",
			1861 => "0000000001110110110101",
			1862 => "0010011001100100000100",
			1863 => "0000001001110110110101",
			1864 => "0000000001110110110101",
			1865 => "0000000110011100000100",
			1866 => "0000000001110110110101",
			1867 => "0011010010011100000100",
			1868 => "1111111001110110110101",
			1869 => "0000000001110110110101",
			1870 => "0010010100111100000100",
			1871 => "0000001001110110110101",
			1872 => "0000000001110110110101",
			1873 => "0000111010000100001000",
			1874 => "0011111010000100000100",
			1875 => "1111111001110110110101",
			1876 => "0000000001110110110101",
			1877 => "0000101100000000000100",
			1878 => "0000000001110110110101",
			1879 => "0011000100011000000100",
			1880 => "0000000001110110110101",
			1881 => "0000000001110110110101",
			1882 => "0001111111011100010000",
			1883 => "0010011000010000001100",
			1884 => "0000100110010000000100",
			1885 => "0000000001110110110101",
			1886 => "0011010101110000000100",
			1887 => "0000000001110110110101",
			1888 => "0000001001110110110101",
			1889 => "0000000001110110110101",
			1890 => "0011011100010100001000",
			1891 => "0011001011000000000100",
			1892 => "0000000001110110110101",
			1893 => "0000000001110110110101",
			1894 => "0010011010100000001100",
			1895 => "0010001001101000001000",
			1896 => "0001100101010000000100",
			1897 => "0000000001110110110101",
			1898 => "0000000001110110110101",
			1899 => "0000000001110110110101",
			1900 => "0000000001110110110101",
			1901 => "0001111101100000000100",
			1902 => "1111111001111001010011",
			1903 => "0010100111101100001000",
			1904 => "0011100100001000000100",
			1905 => "0000000001111001010011",
			1906 => "0000000001111001010011",
			1907 => "0000111010000100101000",
			1908 => "0000111100010000010000",
			1909 => "0000001100011100000100",
			1910 => "0000000001111001010011",
			1911 => "0001110001101000001000",
			1912 => "0011010010011100000100",
			1913 => "1111111001111001010011",
			1914 => "0000000001111001010011",
			1915 => "0000000001111001010011",
			1916 => "0011010111111100001100",
			1917 => "0000010000111100001000",
			1918 => "0001111111011100000100",
			1919 => "0000000001111001010011",
			1920 => "0000000001111001010011",
			1921 => "0000000001111001010011",
			1922 => "0001111111011100001000",
			1923 => "0011001001001000000100",
			1924 => "1111111001111001010011",
			1925 => "0000000001111001010011",
			1926 => "0000000001111001010011",
			1927 => "0011000100011000000100",
			1928 => "0000000001111001010011",
			1929 => "0010010100111100001000",
			1930 => "0001111111011100000100",
			1931 => "0000001001111001010011",
			1932 => "0000000001111001010011",
			1933 => "0000111000100000001000",
			1934 => "0001110001101000000100",
			1935 => "0000000001111001010011",
			1936 => "0000000001111001010011",
			1937 => "0000011101111100000100",
			1938 => "0000000001111001010011",
			1939 => "0000000001111001010011",
			1940 => "0000000001111001010101",
			1941 => "0000000001111001011001",
			1942 => "0000000001111001011101",
			1943 => "0000000001111001100001",
			1944 => "0000000001111001100101",
			1945 => "0000000001111001101001",
			1946 => "0000000001111001101101",
			1947 => "0000000001111001110001",
			1948 => "0011001100110000000100",
			1949 => "0000000001111010000101",
			1950 => "0011000001101000000100",
			1951 => "0000000001111010000101",
			1952 => "0000000001111010000101",
			1953 => "0000110111010100001000",
			1954 => "0000111101010100000100",
			1955 => "0000000001111010100001",
			1956 => "0000000001111010100001",
			1957 => "0000110010100100000100",
			1958 => "0000000001111010100001",
			1959 => "0000000001111010100001",
			1960 => "0000000001010100001100",
			1961 => "0001111101100000000100",
			1962 => "0000000001111010111101",
			1963 => "0001000111001000000100",
			1964 => "0000000001111010111101",
			1965 => "0000000001111010111101",
			1966 => "0000000001111010111101",
			1967 => "0000110111010100001100",
			1968 => "0010010000111100000100",
			1969 => "0000000001111011011001",
			1970 => "0000101010000100000100",
			1971 => "0000000001111011011001",
			1972 => "0000000001111011011001",
			1973 => "0000000001111011011001",
			1974 => "0001011111010000001100",
			1975 => "0001110001101000000100",
			1976 => "0000000001111011111101",
			1977 => "0001011101000100000100",
			1978 => "0000000001111011111101",
			1979 => "0000000001111011111101",
			1980 => "0001110001001000000100",
			1981 => "0000000001111011111101",
			1982 => "0000000001111011111101",
			1983 => "0010010101011100001100",
			1984 => "0011100100001000000100",
			1985 => "0000000001111100100001",
			1986 => "0000001100011100000100",
			1987 => "0000000001111100100001",
			1988 => "0000000001111100100001",
			1989 => "0001101101111100000100",
			1990 => "0000000001111100100001",
			1991 => "0000000001111100100001",
			1992 => "0010110101100100001100",
			1993 => "0011001100110000000100",
			1994 => "0000000001111101001101",
			1995 => "0011001000000000000100",
			1996 => "0000000001111101001101",
			1997 => "0000000001111101001101",
			1998 => "0000010000111100001000",
			1999 => "0001110111010000000100",
			2000 => "0000000001111101001101",
			2001 => "0000000001111101001101",
			2002 => "0000000001111101001101",
			2003 => "0000111010000100001100",
			2004 => "0001110001101000001000",
			2005 => "0001110110000100000100",
			2006 => "0000000001111101111001",
			2007 => "0000000001111101111001",
			2008 => "0000000001111101111001",
			2009 => "0001111000011000000100",
			2010 => "0000000001111101111001",
			2011 => "0001111111011100000100",
			2012 => "0000000001111101111001",
			2013 => "0000000001111101111001",
			2014 => "0010100010101100010000",
			2015 => "0011101110101000000100",
			2016 => "0000000001111110011101",
			2017 => "0010110101110100001000",
			2018 => "0000010000111100000100",
			2019 => "0000000001111110011101",
			2020 => "0000000001111110011101",
			2021 => "0000000001111110011101",
			2022 => "0000000001111110011101",
			2023 => "0010110100010000010000",
			2024 => "0010111000011000000100",
			2025 => "0000000001111111000001",
			2026 => "0000010000111100001000",
			2027 => "0000011111001100000100",
			2028 => "0000000001111111000001",
			2029 => "0000000001111111000001",
			2030 => "0000000001111111000001",
			2031 => "0000000001111111000001",
			2032 => "0000000001010100010000",
			2033 => "0000010000111100001100",
			2034 => "0001111101100000000100",
			2035 => "0000000001111111100101",
			2036 => "0001000111001000000100",
			2037 => "0000000001111111100101",
			2038 => "0000000001111111100101",
			2039 => "0000000001111111100101",
			2040 => "0000000001111111100101",
			2041 => "0001100100110100010000",
			2042 => "0010101010100000001100",
			2043 => "0001100111101000000100",
			2044 => "0000000010000000010001",
			2045 => "0010100000001000000100",
			2046 => "0000000010000000010001",
			2047 => "0000000010000000010001",
			2048 => "0000000010000000010001",
			2049 => "0010100000001000000100",
			2050 => "0000000010000000010001",
			2051 => "0000000010000000010001",
			2052 => "0011100110100100000100",
			2053 => "0000000010000000111101",
			2054 => "0001011111010000001100",
			2055 => "0001010100000100000100",
			2056 => "0000000010000000111101",
			2057 => "0001010101001000000100",
			2058 => "0000000010000000111101",
			2059 => "0000000010000000111101",
			2060 => "0001011111100100000100",
			2061 => "0000000010000000111101",
			2062 => "0000000010000000111101",
			2063 => "0000000110011100010000",
			2064 => "0011011010011100001100",
			2065 => "0001000111001000000100",
			2066 => "0000000010000001110001",
			2067 => "0001111110001100000100",
			2068 => "0000000010000001110001",
			2069 => "0000000010000001110001",
			2070 => "0000000010000001110001",
			2071 => "0001111000011000001000",
			2072 => "0011011110010000000100",
			2073 => "0000000010000001110001",
			2074 => "0000000010000001110001",
			2075 => "0000000010000001110001",
			2076 => "0001100100110100010000",
			2077 => "0010101010100000001100",
			2078 => "0000100111100000000100",
			2079 => "0000000010000010100101",
			2080 => "0010100000001000000100",
			2081 => "0000000010000010100101",
			2082 => "0000000010000010100101",
			2083 => "0000000010000010100101",
			2084 => "0000101110111000001000",
			2085 => "0010100000001000000100",
			2086 => "0000000010000010100101",
			2087 => "0000000010000010100101",
			2088 => "0000000010000010100101",
			2089 => "0001011110010000010100",
			2090 => "0010000111110100001100",
			2091 => "0010100100111100000100",
			2092 => "0000000010000011100001",
			2093 => "0000000110011100000100",
			2094 => "0000000010000011100001",
			2095 => "0000000010000011100001",
			2096 => "0010100111101100000100",
			2097 => "0000000010000011100001",
			2098 => "0000000010000011100001",
			2099 => "0001101000010000001000",
			2100 => "0000011101111100000100",
			2101 => "0000000010000011100001",
			2102 => "0000000010000011100001",
			2103 => "0000000010000011100001",
			2104 => "0011100110100100001000",
			2105 => "0001101101011100000100",
			2106 => "0000000010000100010101",
			2107 => "0000000010000100010101",
			2108 => "0010100000001000010000",
			2109 => "0001100100110100001100",
			2110 => "0010010100111100001000",
			2111 => "0011111010011100000100",
			2112 => "0000000010000100010101",
			2113 => "0000000010000100010101",
			2114 => "0000000010000100010101",
			2115 => "0000000010000100010101",
			2116 => "0000000010000100010101",
			2117 => "0011101110101000001000",
			2118 => "0010001001111100000100",
			2119 => "0000000010000101001001",
			2120 => "0000000010000101001001",
			2121 => "0000010101011100010000",
			2122 => "0001110111010000001100",
			2123 => "0001101010011000001000",
			2124 => "0011000110000100000100",
			2125 => "0000000010000101001001",
			2126 => "0000000010000101001001",
			2127 => "0000000010000101001001",
			2128 => "0000000010000101001001",
			2129 => "0000000010000101001001",
			2130 => "0000000001010100010100",
			2131 => "0000010000111100010000",
			2132 => "0001111101100000000100",
			2133 => "0000000010000101110101",
			2134 => "0011001000000000001000",
			2135 => "0001000111001000000100",
			2136 => "0000000010000101110101",
			2137 => "0000000010000101110101",
			2138 => "0000000010000101110101",
			2139 => "0000000010000101110101",
			2140 => "0000000010000101110101",
			2141 => "0011001100110000001100",
			2142 => "0000001010110000001000",
			2143 => "0000100100001000000100",
			2144 => "0000000010000110111001",
			2145 => "0000000010000110111001",
			2146 => "0000000010000110111001",
			2147 => "0001111000000000001100",
			2148 => "0011001100110000000100",
			2149 => "0000000010000110111001",
			2150 => "0011000100011000000100",
			2151 => "0000000010000110111001",
			2152 => "0000000010000110111001",
			2153 => "0001100100110100001000",
			2154 => "0011001000000000000100",
			2155 => "0000000010000110111001",
			2156 => "0000000010000110111001",
			2157 => "0000000010000110111001",
			2158 => "0000111100010000011000",
			2159 => "0010010000111100001100",
			2160 => "0011100100001000000100",
			2161 => "0000000010001000000101",
			2162 => "0000000101000100000100",
			2163 => "0000000010001000000101",
			2164 => "0000000010001000000101",
			2165 => "0000010110101000000100",
			2166 => "0000000010001000000101",
			2167 => "0011010010011100000100",
			2168 => "0000000010001000000101",
			2169 => "0000000010001000000101",
			2170 => "0010100001010000001100",
			2171 => "0001011110101000000100",
			2172 => "0000000010001000000101",
			2173 => "0000011101111100000100",
			2174 => "0000000010001000000101",
			2175 => "0000000010001000000101",
			2176 => "0000000010001000000101",
			2177 => "0011001100110000001100",
			2178 => "0000101101000100001000",
			2179 => "0011100100001000000100",
			2180 => "0000000010001001010001",
			2181 => "0000000010001001010001",
			2182 => "0000000010001001010001",
			2183 => "0000111010000100010000",
			2184 => "0011001001110100001100",
			2185 => "0000101010000100001000",
			2186 => "0011101100010000000100",
			2187 => "0000000010001001010001",
			2188 => "0000000010001001010001",
			2189 => "0000000010001001010001",
			2190 => "0000000010001001010001",
			2191 => "0010011000010000001000",
			2192 => "0000101101001000000100",
			2193 => "0000000010001001010001",
			2194 => "0000000010001001010001",
			2195 => "0000000010001001010001",
			2196 => "0010011100011000001100",
			2197 => "0010010000111100000100",
			2198 => "0000000010001010011101",
			2199 => "0000010110101000000100",
			2200 => "0000000010001010011101",
			2201 => "0000000010001010011101",
			2202 => "0001000110111100001100",
			2203 => "0011000100011000000100",
			2204 => "0000000010001010011101",
			2205 => "0011001001001000000100",
			2206 => "0000000010001010011101",
			2207 => "0000000010001010011101",
			2208 => "0000010000111100001100",
			2209 => "0011001001110100001000",
			2210 => "0011000111001000000100",
			2211 => "0000000010001010011101",
			2212 => "0000000010001010011101",
			2213 => "0000000010001010011101",
			2214 => "0000000010001010011101",
			2215 => "0001010111100000011100",
			2216 => "0000000110011100001100",
			2217 => "0011111010011100000100",
			2218 => "0000000010001011110001",
			2219 => "0000111001010100000100",
			2220 => "0000000010001011110001",
			2221 => "0000000010001011110001",
			2222 => "0010110010001000001100",
			2223 => "0010100111101100000100",
			2224 => "0000000010001011110001",
			2225 => "0011001001110100000100",
			2226 => "0000000010001011110001",
			2227 => "0000000010001011110001",
			2228 => "0000000010001011110001",
			2229 => "0001101000010000001100",
			2230 => "0000011101111100001000",
			2231 => "0010110101100100000100",
			2232 => "0000000010001011110001",
			2233 => "0000000010001011110001",
			2234 => "0000000010001011110001",
			2235 => "0000000010001011110001",
			2236 => "0000111100010000011000",
			2237 => "0010010000111100001100",
			2238 => "0011100100001000000100",
			2239 => "0000000010001101000101",
			2240 => "0000000101000100000100",
			2241 => "0000000010001101000101",
			2242 => "0000000010001101000101",
			2243 => "0001110101101100000100",
			2244 => "0000000010001101000101",
			2245 => "0011010010011100000100",
			2246 => "0000000010001101000101",
			2247 => "0000000010001101000101",
			2248 => "0010100001010000010000",
			2249 => "0010011010100000001100",
			2250 => "0011011111010000000100",
			2251 => "0000000010001101000101",
			2252 => "0011101100010100000100",
			2253 => "0000000010001101000101",
			2254 => "0000000010001101000101",
			2255 => "0000000010001101000101",
			2256 => "0000000010001101000101",
			2257 => "0010011100011000010100",
			2258 => "0001101101011100000100",
			2259 => "0000000010001110010001",
			2260 => "0001010110100100000100",
			2261 => "0000000010001110010001",
			2262 => "0001111100101000001000",
			2263 => "0001110110000100000100",
			2264 => "0000000010001110010001",
			2265 => "0000000010001110010001",
			2266 => "0000000010001110010001",
			2267 => "0000010000111100010000",
			2268 => "0001111111011100001100",
			2269 => "0001110001111100000100",
			2270 => "0000000010001110010001",
			2271 => "0001101011001100000100",
			2272 => "0000000010001110010001",
			2273 => "0000000010001110010001",
			2274 => "0000000010001110010001",
			2275 => "0000000010001110010001",
			2276 => "0001011111010000011000",
			2277 => "0000000101000100010000",
			2278 => "0011001100110000001100",
			2279 => "0000000110011000001000",
			2280 => "0011001100110000000100",
			2281 => "0000000010001111100101",
			2282 => "0000000010001111100101",
			2283 => "0000000010001111100101",
			2284 => "0000000010001111100101",
			2285 => "0010001000100100000100",
			2286 => "0000000010001111100101",
			2287 => "0000000010001111100101",
			2288 => "0001100101010000010000",
			2289 => "0011001011000000000100",
			2290 => "0000000010001111100101",
			2291 => "0000011101011100000100",
			2292 => "0000000010001111100101",
			2293 => "0000011101111100000100",
			2294 => "0000000010001111100101",
			2295 => "0000000010001111100101",
			2296 => "0000000010001111100101",
			2297 => "0010001001101000011000",
			2298 => "0011100100001000000100",
			2299 => "0000000010010000011001",
			2300 => "0010011111000000010000",
			2301 => "0001111000011000001100",
			2302 => "0001111101100000000100",
			2303 => "0000000010010000011001",
			2304 => "0001101011001100000100",
			2305 => "0000000010010000011001",
			2306 => "0000000010010000011001",
			2307 => "0000000010010000011001",
			2308 => "0000000010010000011001",
			2309 => "0000000010010000011001",
			2310 => "0000000001010100100000",
			2311 => "0011110000011100001100",
			2312 => "0000010110101000001000",
			2313 => "0011100100001000000100",
			2314 => "0000000010010001100101",
			2315 => "0000000010010001100101",
			2316 => "0000000010010001100101",
			2317 => "0011001000000000010000",
			2318 => "0001100100110100001100",
			2319 => "0000010000111100001000",
			2320 => "0010100100111100000100",
			2321 => "0000000010010001100101",
			2322 => "0000000010010001100101",
			2323 => "0000000010010001100101",
			2324 => "0000000010010001100101",
			2325 => "0000000010010001100101",
			2326 => "0001101101111100000100",
			2327 => "0000000010010001100101",
			2328 => "0000000010010001100101",
			2329 => "0001011100100100011100",
			2330 => "0000000110011100001100",
			2331 => "0011111010011100000100",
			2332 => "0000000010010011000001",
			2333 => "0000101010010100000100",
			2334 => "0000000010010011000001",
			2335 => "0000000010010011000001",
			2336 => "0011111100010000001100",
			2337 => "0011010101110000001000",
			2338 => "0010000111110100000100",
			2339 => "0000000010010011000001",
			2340 => "0000000010010011000001",
			2341 => "0000000010010011000001",
			2342 => "0000000010010011000001",
			2343 => "0001101000010000010000",
			2344 => "0001010111100000000100",
			2345 => "0000000010010011000001",
			2346 => "0000011101111100001000",
			2347 => "0010110101100100000100",
			2348 => "0000000010010011000001",
			2349 => "0000000010010011000001",
			2350 => "0000000010010011000001",
			2351 => "0000000010010011000001",
			2352 => "0000111100010000011000",
			2353 => "0010010000111100001100",
			2354 => "0001000110110100001000",
			2355 => "0011100100001000000100",
			2356 => "0000000010010100011101",
			2357 => "0000000010010100011101",
			2358 => "0000000010010100011101",
			2359 => "0011001100110000000100",
			2360 => "0000000010010100011101",
			2361 => "0011101010001000000100",
			2362 => "0000000010010100011101",
			2363 => "0000000010010100011101",
			2364 => "0010011100011000000100",
			2365 => "0000000010010100011101",
			2366 => "0010011010100000010000",
			2367 => "0010100001010000001100",
			2368 => "0011011111010000000100",
			2369 => "0000000010010100011101",
			2370 => "0011000111001000000100",
			2371 => "0000000010010100011101",
			2372 => "0000000010010100011101",
			2373 => "0000000010010100011101",
			2374 => "0000000010010100011101",
			2375 => "0010011100011000001000",
			2376 => "0010010000111100000100",
			2377 => "0000000010010101110001",
			2378 => "0000000010010101110001",
			2379 => "0001000110111100010100",
			2380 => "0011000100011000000100",
			2381 => "0000000010010101110001",
			2382 => "0011001001001000001100",
			2383 => "0010011001100100000100",
			2384 => "0000000010010101110001",
			2385 => "0010100111101100000100",
			2386 => "0000000010010101110001",
			2387 => "0000000010010101110001",
			2388 => "0000000010010101110001",
			2389 => "0010100001010000001100",
			2390 => "0011000111001000000100",
			2391 => "0000000010010101110001",
			2392 => "0010011010100000000100",
			2393 => "0000000010010101110001",
			2394 => "0000000010010101110001",
			2395 => "0000000010010101110001",
			2396 => "0010100000001000011000",
			2397 => "0010010101011100010000",
			2398 => "0000010110101000001100",
			2399 => "0000100100001000000100",
			2400 => "0000000010010111011101",
			2401 => "0000000011101000000100",
			2402 => "0000000010010111011101",
			2403 => "0000000010010111011101",
			2404 => "0000000010010111011101",
			2405 => "0000101101000100000100",
			2406 => "0000000010010111011101",
			2407 => "0000000010010111011101",
			2408 => "0000111010000100001100",
			2409 => "0011111111010100001000",
			2410 => "0000010000111100000100",
			2411 => "0000000010010111011101",
			2412 => "0000000010010111011101",
			2413 => "0000000010010111011101",
			2414 => "0011001011000000000100",
			2415 => "0000000010010111011101",
			2416 => "0001010010011100001100",
			2417 => "0000010000111100001000",
			2418 => "0001111111011100000100",
			2419 => "0000000010010111011101",
			2420 => "0000000010010111011101",
			2421 => "0000000010010111011101",
			2422 => "0000000010010111011101",
			2423 => "0011101100010000100000",
			2424 => "0011000100011000010100",
			2425 => "0011000110000100000100",
			2426 => "0000000010011001000001",
			2427 => "0010010100111100001100",
			2428 => "0010011001011000000100",
			2429 => "0000000010011001000001",
			2430 => "0000000110001000000100",
			2431 => "0000000010011001000001",
			2432 => "0000000010011001000001",
			2433 => "0000000010011001000001",
			2434 => "0001110001101000000100",
			2435 => "0000000010011001000001",
			2436 => "0000000110011100000100",
			2437 => "0000000010011001000001",
			2438 => "0000000010011001000001",
			2439 => "0010110101100100000100",
			2440 => "0000000010011001000001",
			2441 => "0010100001010000001100",
			2442 => "0000011101111100001000",
			2443 => "0001010111100000000100",
			2444 => "0000000010011001000001",
			2445 => "0000000010011001000001",
			2446 => "0000000010011001000001",
			2447 => "0000000010011001000001",
			2448 => "0011010111111100011100",
			2449 => "0000111001001000000100",
			2450 => "0000000010011010001101",
			2451 => "0010101010100000010100",
			2452 => "0011000011011100000100",
			2453 => "0000000010011010001101",
			2454 => "0000010000111100001100",
			2455 => "0001110110000100000100",
			2456 => "0000000010011010001101",
			2457 => "0001111000011000000100",
			2458 => "0000000010011010001101",
			2459 => "0000000010011010001101",
			2460 => "0000000010011010001101",
			2461 => "0000000010011010001101",
			2462 => "0010101010100000001000",
			2463 => "0000101100000000000100",
			2464 => "0000000010011010001101",
			2465 => "0000000010011010001101",
			2466 => "0000000010011010001101",
			2467 => "0000111000011000001000",
			2468 => "0001101101011100000100",
			2469 => "0000000010011011010001",
			2470 => "0000000010011011010001",
			2471 => "0010100000001000011000",
			2472 => "0001100100110100010100",
			2473 => "0001100000111100000100",
			2474 => "0000000010011011010001",
			2475 => "0010110100001000000100",
			2476 => "0000000010011011010001",
			2477 => "0010010100111100001000",
			2478 => "0011111010011100000100",
			2479 => "0000000010011011010001",
			2480 => "0000000010011011010001",
			2481 => "0000000010011011010001",
			2482 => "0000000010011011010001",
			2483 => "0000000010011011010001",
			2484 => "0001010101001000010000",
			2485 => "0001100001000100000100",
			2486 => "0000000010011100100101",
			2487 => "0000011001011000001000",
			2488 => "0011001001110100000100",
			2489 => "0000000010011100100101",
			2490 => "0000000010011100100101",
			2491 => "0000000010011100100101",
			2492 => "0001111000011000000100",
			2493 => "0000000010011100100101",
			2494 => "0001100101010000010100",
			2495 => "0011001011000000000100",
			2496 => "0000000010011100100101",
			2497 => "0010110010001000000100",
			2498 => "0000000010011100100101",
			2499 => "0000011101111100001000",
			2500 => "0000011101011100000100",
			2501 => "0000000010011100100101",
			2502 => "0000000010011100100101",
			2503 => "0000000010011100100101",
			2504 => "0000000010011100100101",
			2505 => "0011010111111100011100",
			2506 => "0000111001001000000100",
			2507 => "0000000010011101100001",
			2508 => "0010010100111100010100",
			2509 => "0011000011011100000100",
			2510 => "0000000010011101100001",
			2511 => "0011001011000000001100",
			2512 => "0001100000111100000100",
			2513 => "0000000010011101100001",
			2514 => "0011111010011100000100",
			2515 => "0000000010011101100001",
			2516 => "0000000010011101100001",
			2517 => "0000000010011101100001",
			2518 => "0000000010011101100001",
			2519 => "0000000010011101100001",
			2520 => "0000111000001100101100",
			2521 => "0010100000001000100000",
			2522 => "0011111001001000001100",
			2523 => "0000010110101000001000",
			2524 => "0011100100001000000100",
			2525 => "0000000010011111001101",
			2526 => "0000000010011111001101",
			2527 => "0000000010011111001101",
			2528 => "0000101110110100010000",
			2529 => "0000010000111100001100",
			2530 => "0011101011000000000100",
			2531 => "0000000010011111001101",
			2532 => "0010110100001000000100",
			2533 => "0000000010011111001101",
			2534 => "0000000010011111001101",
			2535 => "0000000010011111001101",
			2536 => "0000000010011111001101",
			2537 => "0011110000010000001000",
			2538 => "0010110100010000000100",
			2539 => "0000000010011111001101",
			2540 => "0000000010011111001101",
			2541 => "0000000010011111001101",
			2542 => "0000010101011100001000",
			2543 => "0001110111010000000100",
			2544 => "0000000010011111001101",
			2545 => "0000000010011111001101",
			2546 => "0000000010011111001101",
			2547 => "0001010110100100001100",
			2548 => "0011000110000100001000",
			2549 => "0001101101011100000100",
			2550 => "0000000010100001000001",
			2551 => "1111111010100001000001",
			2552 => "0000000010100001000001",
			2553 => "0000111111010100011100",
			2554 => "0000011001011000010000",
			2555 => "0000110000110100000100",
			2556 => "0000000010100001000001",
			2557 => "0011001000000000001000",
			2558 => "0011000011011100000100",
			2559 => "0000000010100001000001",
			2560 => "0000000010100001000001",
			2561 => "0000000010100001000001",
			2562 => "0011000100011000000100",
			2563 => "0000000010100001000001",
			2564 => "0011001001110100000100",
			2565 => "0000000010100001000001",
			2566 => "0000000010100001000001",
			2567 => "0010010100111100010000",
			2568 => "0000110010010100001100",
			2569 => "0011001001110100001000",
			2570 => "0000111010000100000100",
			2571 => "0000000010100001000001",
			2572 => "0000000010100001000001",
			2573 => "0000000010100001000001",
			2574 => "0000000010100001000001",
			2575 => "0000000010100001000001",
			2576 => "0000000001010100110100",
			2577 => "0000101110010000100000",
			2578 => "0000011101011100011000",
			2579 => "0011000011011100001000",
			2580 => "0010110101101100000100",
			2581 => "0000000010100011001101",
			2582 => "0000000010100011001101",
			2583 => "0001101001011000000100",
			2584 => "0000000010100011001101",
			2585 => "0001110110000100000100",
			2586 => "0000000010100011001101",
			2587 => "0001110000001100000100",
			2588 => "0000000010100011001101",
			2589 => "0000000010100011001101",
			2590 => "0000111001100000000100",
			2591 => "0000000010100011001101",
			2592 => "0000000010100011001101",
			2593 => "0011111100000000001100",
			2594 => "0001100100110100001000",
			2595 => "0000010000111100000100",
			2596 => "0000000010100011001101",
			2597 => "0000000010100011001101",
			2598 => "0000000010100011001101",
			2599 => "0001111000011000000100",
			2600 => "0000000010100011001101",
			2601 => "0000000010100011001101",
			2602 => "0011111111010100001000",
			2603 => "0000111000001100000100",
			2604 => "0000000010100011001101",
			2605 => "0000000010100011001101",
			2606 => "0000010000111100001000",
			2607 => "0000011111001100000100",
			2608 => "0000000010100011001101",
			2609 => "0000000010100011001101",
			2610 => "0000000010100011001101",
			2611 => "0001100100110100100100",
			2612 => "0001000010010100100000",
			2613 => "0011001001110100011100",
			2614 => "0000100110010000010100",
			2615 => "0001111100101000001100",
			2616 => "0010000010101100001000",
			2617 => "0000100100001000000100",
			2618 => "0000000010100100101001",
			2619 => "0000000010100100101001",
			2620 => "0000000010100100101001",
			2621 => "0011001000000000000100",
			2622 => "0000000010100100101001",
			2623 => "0000000010100100101001",
			2624 => "0000010000111100000100",
			2625 => "0000000010100100101001",
			2626 => "0000000010100100101001",
			2627 => "0000000010100100101001",
			2628 => "0000000010100100101001",
			2629 => "0011110110001100001000",
			2630 => "0010001000100100000100",
			2631 => "0000000010100100101001",
			2632 => "0000000010100100101001",
			2633 => "0000000010100100101001",
			2634 => "0010110010001000101100",
			2635 => "0010100111101100100000",
			2636 => "0000001010100100010000",
			2637 => "0000010110101000001100",
			2638 => "0000100100001000000100",
			2639 => "0000000010100110101101",
			2640 => "0010010000111100000100",
			2641 => "0000000010100110101101",
			2642 => "0000000010100110101101",
			2643 => "0000000010100110101101",
			2644 => "0010100100111100000100",
			2645 => "0000000010100110101101",
			2646 => "0011110010001000000100",
			2647 => "0000000010100110101101",
			2648 => "0001101101111100000100",
			2649 => "0000000010100110101101",
			2650 => "0000000010100110101101",
			2651 => "0000111100000000001000",
			2652 => "0000000110011100000100",
			2653 => "0000000010100110101101",
			2654 => "0000000010100110101101",
			2655 => "0000000010100110101101",
			2656 => "0010010100111100010100",
			2657 => "0010111011110100010000",
			2658 => "0011001011000000000100",
			2659 => "0000000010100110101101",
			2660 => "0011100110010000000100",
			2661 => "0000000010100110101101",
			2662 => "0011001001110100000100",
			2663 => "0000000010100110101101",
			2664 => "0000000010100110101101",
			2665 => "0000000010100110101101",
			2666 => "0000000010100110101101",
			2667 => "0010001001000100101100",
			2668 => "0011101000011000001100",
			2669 => "0011101011000000000100",
			2670 => "1111111010101001001001",
			2671 => "0011011111011100000100",
			2672 => "0000010010101001001001",
			2673 => "1111111010101001001001",
			2674 => "0000010000111100011000",
			2675 => "0001111111011100010100",
			2676 => "0010110101110100010000",
			2677 => "0011101100010000001000",
			2678 => "0001100100110100000100",
			2679 => "0000001010101001001001",
			2680 => "0000000010101001001001",
			2681 => "0011001000000000000100",
			2682 => "0000010010101001001001",
			2683 => "0000001010101001001001",
			2684 => "1111111010101001001001",
			2685 => "1111111010101001001001",
			2686 => "0011010011001000000100",
			2687 => "1111111010101001001001",
			2688 => "0000000010101001001001",
			2689 => "0010000001010000010000",
			2690 => "0001001101101100001100",
			2691 => "0000010000111100001000",
			2692 => "0001001000001100000100",
			2693 => "1111111010101001001001",
			2694 => "0000001010101001001001",
			2695 => "1111111010101001001001",
			2696 => "0000010010101001001001",
			2697 => "0011010011000000001100",
			2698 => "0010001100011100001000",
			2699 => "0010001010110000000100",
			2700 => "1111111010101001001001",
			2701 => "0000000010101001001001",
			2702 => "1111111010101001001001",
			2703 => "0010001110111100000100",
			2704 => "0000010010101001001001",
			2705 => "1111111010101001001001",
			2706 => "0011000011011100001100",
			2707 => "0011011010001100001000",
			2708 => "0010101100011000000100",
			2709 => "0000000010101011010101",
			2710 => "1111111010101011010101",
			2711 => "0000000010101011010101",
			2712 => "0000111111010100100100",
			2713 => "0011001011000000011000",
			2714 => "0011011110101000010000",
			2715 => "0001111101111000001100",
			2716 => "0001110110000100000100",
			2717 => "0000000010101011010101",
			2718 => "0011000110000100000100",
			2719 => "0000000010101011010101",
			2720 => "0000000010101011010101",
			2721 => "0000000010101011010101",
			2722 => "0010010100111100000100",
			2723 => "0000000010101011010101",
			2724 => "0000000010101011010101",
			2725 => "0000011001011000001000",
			2726 => "0010000111110100000100",
			2727 => "0000000010101011010101",
			2728 => "0000000010101011010101",
			2729 => "0000000010101011010101",
			2730 => "0000010000111100001000",
			2731 => "0001111111011100000100",
			2732 => "0000000010101011010101",
			2733 => "0000000010101011010101",
			2734 => "0011010110010000000100",
			2735 => "0000000010101011010101",
			2736 => "0011001011011100001000",
			2737 => "0011100000010100000100",
			2738 => "0000000010101011010101",
			2739 => "0000000010101011010101",
			2740 => "0000000010101011010101",
			2741 => "0010101010100000110000",
			2742 => "0011100101110100011000",
			2743 => "0001101101011100001000",
			2744 => "0011100100001000000100",
			2745 => "1111111010101110001001",
			2746 => "0000010010101110001001",
			2747 => "0010110100001000000100",
			2748 => "1111111010101110001001",
			2749 => "0010010001000100001000",
			2750 => "0001010001101000000100",
			2751 => "0000000010101110001001",
			2752 => "0000010010101110001001",
			2753 => "1111111010101110001001",
			2754 => "0010010100111100010100",
			2755 => "0001111111011100010000",
			2756 => "0000111010000100001100",
			2757 => "0001011111010000001000",
			2758 => "0011101110101000000100",
			2759 => "0000001010101110001001",
			2760 => "0000001010101110001001",
			2761 => "0000000010101110001001",
			2762 => "0000010010101110001001",
			2763 => "0000000010101110001001",
			2764 => "1111111010101110001001",
			2765 => "0010100010101100011000",
			2766 => "0000101010000100001100",
			2767 => "0000111000001100000100",
			2768 => "1111111010101110001001",
			2769 => "0001111000011000000100",
			2770 => "0000001010101110001001",
			2771 => "1111111010101110001001",
			2772 => "0010010101010000001000",
			2773 => "0001001000100000000100",
			2774 => "0000001010101110001001",
			2775 => "0000010010101110001001",
			2776 => "1111111010101110001001",
			2777 => "0010100010101100001000",
			2778 => "0011010100101000000100",
			2779 => "1111111010101110001001",
			2780 => "0000001010101110001001",
			2781 => "0011010011000000000100",
			2782 => "1111111010101110001001",
			2783 => "0010110111111100000100",
			2784 => "0000001010101110001001",
			2785 => "1111111010101110001001",
			2786 => "0001010110100100001100",
			2787 => "0001000001101000000100",
			2788 => "0000000010110000001101",
			2789 => "0011101000011000000100",
			2790 => "0000000010110000001101",
			2791 => "0000000010110000001101",
			2792 => "0010100000001000010000",
			2793 => "0011101011000000000100",
			2794 => "0000000010110000001101",
			2795 => "0010110100001000000100",
			2796 => "0000000010110000001101",
			2797 => "0010010100111100000100",
			2798 => "0000000010110000001101",
			2799 => "0000000010110000001101",
			2800 => "0000111000001100010100",
			2801 => "0001010111100000000100",
			2802 => "0000000010110000001101",
			2803 => "0010101010100100001100",
			2804 => "0011010101110000000100",
			2805 => "0000000010110000001101",
			2806 => "0010110101110100000100",
			2807 => "0000000010110000001101",
			2808 => "0000000010110000001101",
			2809 => "0000000010110000001101",
			2810 => "0011101000101000010000",
			2811 => "0001010111100000000100",
			2812 => "0000000010110000001101",
			2813 => "0010110001001000001000",
			2814 => "0010100001010000000100",
			2815 => "0000000010110000001101",
			2816 => "0000000010110000001101",
			2817 => "0000000010110000001101",
			2818 => "0000000010110000001101",
			2819 => "0000111100010000101000",
			2820 => "0010100111101100011100",
			2821 => "0011000110000100010100",
			2822 => "0011111010011100001000",
			2823 => "0010110101101100000100",
			2824 => "0000000010110010110001",
			2825 => "0000000010110010110001",
			2826 => "0011001000111100000100",
			2827 => "0000000010110010110001",
			2828 => "0001111100101000000100",
			2829 => "0000000010110010110001",
			2830 => "0000000010110010110001",
			2831 => "0000101100100100000100",
			2832 => "0000000010110010110001",
			2833 => "0000000010110010110001",
			2834 => "0010000111110100000100",
			2835 => "0000000010110010110001",
			2836 => "0001110001101000000100",
			2837 => "0000000010110010110001",
			2838 => "0000000010110010110001",
			2839 => "0010011100011000000100",
			2840 => "0000000010110010110001",
			2841 => "0010010100111100011100",
			2842 => "0011001000000000001100",
			2843 => "0001100100110100001000",
			2844 => "0001000010000100000100",
			2845 => "0000000010110010110001",
			2846 => "0000000010110010110001",
			2847 => "0000000010110010110001",
			2848 => "0011011010001000001000",
			2849 => "0011010111111100000100",
			2850 => "0000000010110010110001",
			2851 => "0000000010110010110001",
			2852 => "0011011100000000000100",
			2853 => "0000000010110010110001",
			2854 => "0000000010110010110001",
			2855 => "0000111000100000000100",
			2856 => "0000000010110010110001",
			2857 => "0011011010001000000100",
			2858 => "0000000010110010110001",
			2859 => "0000000010110010110001",
			2860 => "0010101010100000110000",
			2861 => "0011101000011000001100",
			2862 => "0011101011000000000100",
			2863 => "1111111010110101010101",
			2864 => "0011011111011100000100",
			2865 => "0000011010110101010101",
			2866 => "1111111010110101010101",
			2867 => "0010010100111100100000",
			2868 => "0010110101110100011100",
			2869 => "0011101100010000010000",
			2870 => "0010100000001000001000",
			2871 => "0010011110010100000100",
			2872 => "0000010010110101010101",
			2873 => "0000001010110101010101",
			2874 => "0010011111000000000100",
			2875 => "0000001010110101010101",
			2876 => "0000000010110101010101",
			2877 => "0011001001110100001000",
			2878 => "0011001000000000000100",
			2879 => "0000011010110101010101",
			2880 => "0000010010110101010101",
			2881 => "0000000010110101010101",
			2882 => "1111111010110101010101",
			2883 => "1111111010110101010101",
			2884 => "0010100010101100010000",
			2885 => "0000101010000100001000",
			2886 => "0010110101110100000100",
			2887 => "1111111010110101010101",
			2888 => "0000000010110101010101",
			2889 => "0000010101011100000100",
			2890 => "0000010010110101010101",
			2891 => "1111111010110101010101",
			2892 => "0011010011000000001100",
			2893 => "0010100011101000001000",
			2894 => "0010100011101000000100",
			2895 => "1111111010110101010101",
			2896 => "0000000010110101010101",
			2897 => "1111111010110101010101",
			2898 => "0000100011111000000100",
			2899 => "0000011010110101010101",
			2900 => "1111111010110101010101",
			2901 => "0011000011011100001000",
			2902 => "0001101101011100000100",
			2903 => "0000000010110111100001",
			2904 => "0000000010110111100001",
			2905 => "0011010111111100100100",
			2906 => "0001100100110100011000",
			2907 => "0011111100100100010000",
			2908 => "0011000110000100001100",
			2909 => "0001101001011000000100",
			2910 => "0000000010110111100001",
			2911 => "0001110110000100000100",
			2912 => "0000000010110111100001",
			2913 => "0000000010110111100001",
			2914 => "0000000010110111100001",
			2915 => "0010010100111100000100",
			2916 => "0000000010110111100001",
			2917 => "0000000010110111100001",
			2918 => "0001011111010000001000",
			2919 => "0010100000001000000100",
			2920 => "0000000010110111100001",
			2921 => "0000000010110111100001",
			2922 => "0000000010110111100001",
			2923 => "0000111000001100001000",
			2924 => "0011011010001000000100",
			2925 => "0000000010110111100001",
			2926 => "0000000010110111100001",
			2927 => "0001101000010000010000",
			2928 => "0011001011000000000100",
			2929 => "0000000010110111100001",
			2930 => "0001101010011000000100",
			2931 => "0000000010110111100001",
			2932 => "0010011010100000000100",
			2933 => "0000000010110111100001",
			2934 => "0000000010110111100001",
			2935 => "0000000010110111100001",
			2936 => "0001110110000100010000",
			2937 => "0011111011000000000100",
			2938 => "0000000010111001110101",
			2939 => "0001011010011100001000",
			2940 => "0001101001011000000100",
			2941 => "0000000010111001110101",
			2942 => "0000000010111001110101",
			2943 => "0000000010111001110101",
			2944 => "0001110001101000010100",
			2945 => "0000001100000100010000",
			2946 => "0001100000111100000100",
			2947 => "0000000010111001110101",
			2948 => "0010011111000000001000",
			2949 => "0011111010011100000100",
			2950 => "0000000010111001110101",
			2951 => "0000000010111001110101",
			2952 => "0000000010111001110101",
			2953 => "0000000010111001110101",
			2954 => "0001111000011000010100",
			2955 => "0011000100011000000100",
			2956 => "0000000010111001110101",
			2957 => "0001001000110100001100",
			2958 => "0001101101111100000100",
			2959 => "0000000010111001110101",
			2960 => "0011011001010000000100",
			2961 => "0000000010111001110101",
			2962 => "0000000010111001110101",
			2963 => "0000000010111001110101",
			2964 => "0011001011000000000100",
			2965 => "0000000010111001110101",
			2966 => "0011010100101000000100",
			2967 => "0000000010111001110101",
			2968 => "0001101000010000001000",
			2969 => "0001010001000000000100",
			2970 => "0000000010111001110101",
			2971 => "0000000010111001110101",
			2972 => "0000000010111001110101",
			2973 => "0010101010100100110100",
			2974 => "0001110110000100010000",
			2975 => "0010111100101000001100",
			2976 => "0010110000001100000100",
			2977 => "1111111010111100100001",
			2978 => "0001011001110100000100",
			2979 => "0000000010111100100001",
			2980 => "0000000010111100100001",
			2981 => "1111110010111100100001",
			2982 => "0000010110101000000100",
			2983 => "0000110010111100100001",
			2984 => "0010010100111100011100",
			2985 => "0011111011011100001100",
			2986 => "0000010111100100001000",
			2987 => "0000010111100100000100",
			2988 => "0000000010111100100001",
			2989 => "0000000010111100100001",
			2990 => "1111111010111100100001",
			2991 => "0011001001110100001000",
			2992 => "0011111111010100000100",
			2993 => "0000001010111100100001",
			2994 => "0000010010111100100001",
			2995 => "0010001000100100000100",
			2996 => "0000001010111100100001",
			2997 => "1111111010111100100001",
			2998 => "1111111010111100100001",
			2999 => "0010100111110100010000",
			3000 => "0000101000100000001100",
			3001 => "0010110101100100000100",
			3002 => "1111111010111100100001",
			3003 => "0010111011011100000100",
			3004 => "0000001010111100100001",
			3005 => "1111111010111100100001",
			3006 => "0000010010111100100001",
			3007 => "0001011111100100001100",
			3008 => "0000100010110000000100",
			3009 => "1111111010111100100001",
			3010 => "0000101000001000000100",
			3011 => "0000011010111100100001",
			3012 => "1111111010111100100001",
			3013 => "0011001011011100000100",
			3014 => "0000010010111100100001",
			3015 => "1111111010111100100001",
			3016 => "0010001001000100101100",
			3017 => "0011101011000000000100",
			3018 => "1111111010111110111101",
			3019 => "0000010000111100100000",
			3020 => "0001111111011100011100",
			3021 => "0011101110101000010000",
			3022 => "0011001100110000001000",
			3023 => "0010110100001000000100",
			3024 => "0000000010111110111101",
			3025 => "0000010010111110111101",
			3026 => "0001111101111000000100",
			3027 => "0000000010111110111101",
			3028 => "1111111010111110111101",
			3029 => "0010110101110100001000",
			3030 => "0011101100010000000100",
			3031 => "0000001010111110111101",
			3032 => "0000010010111110111101",
			3033 => "1111111010111110111101",
			3034 => "1111111010111110111101",
			3035 => "0011010011001000000100",
			3036 => "1111111010111110111101",
			3037 => "0000000010111110111101",
			3038 => "0010100010101100001100",
			3039 => "0011111010000100000100",
			3040 => "1111111010111110111101",
			3041 => "0000010101011100000100",
			3042 => "0000010010111110111101",
			3043 => "1111111010111110111101",
			3044 => "0011010011000000010000",
			3045 => "0010100011101000001100",
			3046 => "0010100011101000000100",
			3047 => "1111111010111110111101",
			3048 => "0010001010110000000100",
			3049 => "1111111010111110111101",
			3050 => "0000001010111110111101",
			3051 => "1111111010111110111101",
			3052 => "0011100011010100000100",
			3053 => "0000010010111110111101",
			3054 => "1111111010111110111101",
			3055 => "0010001000100100110100",
			3056 => "0011110010001000011100",
			3057 => "0011100110100100010100",
			3058 => "0001101101011100001000",
			3059 => "0001011110110000000100",
			3060 => "1111111011000010010001",
			3061 => "0000100011000010010001",
			3062 => "0011101011000000000100",
			3063 => "1111111011000010010001",
			3064 => "0011011111011100000100",
			3065 => "0000010011000010010001",
			3066 => "1111111011000010010001",
			3067 => "0001100000111100000100",
			3068 => "0001010011000010010001",
			3069 => "1111111011000010010001",
			3070 => "0010010100111100010100",
			3071 => "0010111110110000000100",
			3072 => "0000110011000010010001",
			3073 => "0000101100100100000100",
			3074 => "1111111011000010010001",
			3075 => "0000111010000100001000",
			3076 => "0000100010000100000100",
			3077 => "0000011011000010010001",
			3078 => "0000001011000010010001",
			3079 => "0000100011000010010001",
			3080 => "1111111011000010010001",
			3081 => "0000001001101000011000",
			3082 => "0000010000111100001100",
			3083 => "0000100111011000001000",
			3084 => "0010011111000000000100",
			3085 => "0000010011000010010001",
			3086 => "1111111011000010010001",
			3087 => "0000111011000010010001",
			3088 => "0000110000010000000100",
			3089 => "1111111011000010010001",
			3090 => "0010110101110100000100",
			3091 => "0000100011000010010001",
			3092 => "1111111011000010010001",
			3093 => "0010100010101100001100",
			3094 => "0011011111010000000100",
			3095 => "1111111011000010010001",
			3096 => "0000001001101000000100",
			3097 => "1111111011000010010001",
			3098 => "0000011011000010010001",
			3099 => "0011010011000000000100",
			3100 => "1111111011000010010001",
			3101 => "0011010010010100001100",
			3102 => "0001011000100000001000",
			3103 => "0001011111100100000100",
			3104 => "0000000011000010010001",
			3105 => "0000001011000010010001",
			3106 => "1111111011000010010001",
			3107 => "1111111011000010010001",
			3108 => "0010010100111100111100",
			3109 => "0011101010001000011100",
			3110 => "0000001100011100011000",
			3111 => "0001110000001100010000",
			3112 => "0011000011011100000100",
			3113 => "0000000011000100010101",
			3114 => "0011011000011000000100",
			3115 => "0000000011000100010101",
			3116 => "0011000110000100000100",
			3117 => "0000000011000100010101",
			3118 => "0000000011000100010101",
			3119 => "0011010000110100000100",
			3120 => "0000000011000100010101",
			3121 => "0000000011000100010101",
			3122 => "0000000011000100010101",
			3123 => "0001111111011100011100",
			3124 => "0001111000011000010100",
			3125 => "0001110001101000001100",
			3126 => "0011010111111100001000",
			3127 => "0000000010101000000100",
			3128 => "0000000011000100010101",
			3129 => "0000000011000100010101",
			3130 => "0000000011000100010101",
			3131 => "0000011001011000000100",
			3132 => "0000000011000100010101",
			3133 => "0000000011000100010101",
			3134 => "0000111100000000000100",
			3135 => "0000000011000100010101",
			3136 => "0000000011000100010101",
			3137 => "0000000011000100010101",
			3138 => "0000010000111100000100",
			3139 => "0000000011000100010101",
			3140 => "0000000011000100010101",
			3141 => "0000000001010100110000",
			3142 => "0000010000111100101100",
			3143 => "0001111000011000101000",
			3144 => "0010100100111100011000",
			3145 => "0010010101011100001100",
			3146 => "0011100100001000000100",
			3147 => "0000000011000110101001",
			3148 => "0000010110101000000100",
			3149 => "0000000011000110101001",
			3150 => "0000000011000110101001",
			3151 => "0001101001011000000100",
			3152 => "0000000011000110101001",
			3153 => "0010101001100100000100",
			3154 => "0000000011000110101001",
			3155 => "0000000011000110101001",
			3156 => "0000010111100100000100",
			3157 => "0000000011000110101001",
			3158 => "0010010100111100001000",
			3159 => "0011110010001000000100",
			3160 => "0000000011000110101001",
			3161 => "0000000011000110101001",
			3162 => "0000000011000110101001",
			3163 => "0000000011000110101001",
			3164 => "0000000011000110101001",
			3165 => "0010110101100100001000",
			3166 => "0000000001110000000100",
			3167 => "0000000011000110101001",
			3168 => "1111111011000110101001",
			3169 => "0010110110110100001000",
			3170 => "0010010100111100000100",
			3171 => "0000000011000110101001",
			3172 => "0000000011000110101001",
			3173 => "0001011110010000001000",
			3174 => "0011000100011000000100",
			3175 => "0000000011000110101001",
			3176 => "0000000011000110101001",
			3177 => "0000000011000110101001",
			3178 => "0000001011010101001100",
			3179 => "0001100100110100101000",
			3180 => "0011101110101000010100",
			3181 => "0001100001000100010000",
			3182 => "0011000110000100001100",
			3183 => "0011100100001000000100",
			3184 => "0000000011001001011101",
			3185 => "0000010110101000000100",
			3186 => "0000001011001001011101",
			3187 => "0000000011001001011101",
			3188 => "0000000011001001011101",
			3189 => "1111111011001001011101",
			3190 => "0010101010100000010000",
			3191 => "0000010000111100001100",
			3192 => "0011000100011000000100",
			3193 => "0000001011001001011101",
			3194 => "0011000100011000000100",
			3195 => "0000000011001001011101",
			3196 => "0000001011001001011101",
			3197 => "0000000011001001011101",
			3198 => "0000000011001001011101",
			3199 => "0000111000001100011000",
			3200 => "0001000111011000010000",
			3201 => "0001010111100000001000",
			3202 => "0011001010111000000100",
			3203 => "0000000011001001011101",
			3204 => "0000000011001001011101",
			3205 => "0000010000111100000100",
			3206 => "0000001011001001011101",
			3207 => "0000000011001001011101",
			3208 => "0000011001011000000100",
			3209 => "0000000011001001011101",
			3210 => "1111111011001001011101",
			3211 => "0000010101011100001000",
			3212 => "0011001001110100000100",
			3213 => "0000001011001001011101",
			3214 => "0000000011001001011101",
			3215 => "0000000011001001011101",
			3216 => "0000100010110000000100",
			3217 => "1111111011001001011101",
			3218 => "0001100101010000001000",
			3219 => "0000011101011100000100",
			3220 => "0000000011001001011101",
			3221 => "0000001011001001011101",
			3222 => "1111111011001001011101",
			3223 => "0011011000011000001000",
			3224 => "0001101101011100000100",
			3225 => "0000000011001100000001",
			3226 => "1111111011001100000001",
			3227 => "0010101010100000100000",
			3228 => "0001100100110100010100",
			3229 => "0011000011011100000100",
			3230 => "0000000011001100000001",
			3231 => "0000110110100100000100",
			3232 => "0000000011001100000001",
			3233 => "0011001001110100001000",
			3234 => "0010010100111100000100",
			3235 => "0000000011001100000001",
			3236 => "0000000011001100000001",
			3237 => "0000000011001100000001",
			3238 => "0000111010000100001000",
			3239 => "0001110001101000000100",
			3240 => "0000000011001100000001",
			3241 => "0000000011001100000001",
			3242 => "0000000011001100000001",
			3243 => "0000111000001100010000",
			3244 => "0010011111000000001100",
			3245 => "0010011010011000000100",
			3246 => "0000000011001100000001",
			3247 => "0000101011101100000100",
			3248 => "0000000011001100000001",
			3249 => "0000000011001100000001",
			3250 => "0000000011001100000001",
			3251 => "0001101010011000010000",
			3252 => "0001110111010000001100",
			3253 => "0010010101010000001000",
			3254 => "0010001000010100000100",
			3255 => "0000000011001100000001",
			3256 => "0000000011001100000001",
			3257 => "0000000011001100000001",
			3258 => "0000000011001100000001",
			3259 => "0011011111101000000100",
			3260 => "0000000011001100000001",
			3261 => "0011000010001000000100",
			3262 => "0000000011001100000001",
			3263 => "0000000011001100000001",
			3264 => "0000001101010001001100",
			3265 => "0010101010100000101000",
			3266 => "0001100100110100011000",
			3267 => "0001101001011000001000",
			3268 => "0000010110101000000100",
			3269 => "0000000011001110011101",
			3270 => "0000000011001110011101",
			3271 => "0011000011011100000100",
			3272 => "0000000011001110011101",
			3273 => "0001110110000100000100",
			3274 => "0000000011001110011101",
			3275 => "0000010000111100000100",
			3276 => "0000000011001110011101",
			3277 => "0000000011001110011101",
			3278 => "0000111010000100001100",
			3279 => "0000011001011000000100",
			3280 => "0000000011001110011101",
			3281 => "0010001000100100000100",
			3282 => "0000000011001110011101",
			3283 => "0000000011001110011101",
			3284 => "0000000011001110011101",
			3285 => "0000111000001100010000",
			3286 => "0000100110101100001100",
			3287 => "0011111100000000001000",
			3288 => "0011111100010000000100",
			3289 => "0000000011001110011101",
			3290 => "0000000011001110011101",
			3291 => "0000000011001110011101",
			3292 => "0000000011001110011101",
			3293 => "0000010101011100001100",
			3294 => "0001110111010000001000",
			3295 => "0010001000010100000100",
			3296 => "0000000011001110011101",
			3297 => "0000000011001110011101",
			3298 => "0000000011001110011101",
			3299 => "0001110111110000000100",
			3300 => "0000000011001110011101",
			3301 => "0000000011001110011101",
			3302 => "1111111011001110011101",
			3303 => "0000001011010101001100",
			3304 => "0010011111000000011000",
			3305 => "0001111101100000000100",
			3306 => "0000000011010001001001",
			3307 => "0001011111010000010000",
			3308 => "0001111111011100001100",
			3309 => "0011101110101000001000",
			3310 => "0011111001110100000100",
			3311 => "0000001011010001001001",
			3312 => "0000000011010001001001",
			3313 => "0000001011010001001001",
			3314 => "0000000011010001001001",
			3315 => "0000000011010001001001",
			3316 => "0001010101001000010100",
			3317 => "0000000101000100001000",
			3318 => "0011010101110000000100",
			3319 => "0000000011010001001001",
			3320 => "0000000011010001001001",
			3321 => "0001000110111100001000",
			3322 => "0001110110100100000100",
			3323 => "0000000011010001001001",
			3324 => "1111111011010001001001",
			3325 => "0000000011010001001001",
			3326 => "0001111000011000010100",
			3327 => "0001001010000100001000",
			3328 => "0011010111111100000100",
			3329 => "0000000011010001001001",
			3330 => "0000000011010001001001",
			3331 => "0001111000011000001000",
			3332 => "0001111000011000000100",
			3333 => "0000000011010001001001",
			3334 => "0000000011010001001001",
			3335 => "0000000011010001001001",
			3336 => "0001110111010000001000",
			3337 => "0000010101011100000100",
			3338 => "0000000011010001001001",
			3339 => "0000000011010001001001",
			3340 => "0000000011010001001001",
			3341 => "0011110110001100000100",
			3342 => "1111111011010001001001",
			3343 => "0001101000010000000100",
			3344 => "0000000011010001001001",
			3345 => "0000000011010001001001",
			3346 => "0000001001101001000100",
			3347 => "0011101110101000011000",
			3348 => "0000100000110100010100",
			3349 => "0000011101101000010000",
			3350 => "0011100001101000001100",
			3351 => "0000010110101000001000",
			3352 => "0011010110100100000100",
			3353 => "0000000011010100001101",
			3354 => "0000001011010100001101",
			3355 => "1111111011010100001101",
			3356 => "0000001011010100001101",
			3357 => "1111111011010100001101",
			3358 => "1111111011010100001101",
			3359 => "0010011111000000001000",
			3360 => "0010110010001000000100",
			3361 => "0000001011010100001101",
			3362 => "0000000011010100001101",
			3363 => "0000111100000000001000",
			3364 => "0010100000001000000100",
			3365 => "0000000011010100001101",
			3366 => "1111111011010100001101",
			3367 => "0011001000000000010000",
			3368 => "0000000001110000001000",
			3369 => "0000110110111100000100",
			3370 => "0000000011010100001101",
			3371 => "0000001011010100001101",
			3372 => "0011101111010100000100",
			3373 => "0000000011010100001101",
			3374 => "0000000011010100001101",
			3375 => "0010011111000000000100",
			3376 => "1111111011010100001101",
			3377 => "0011011010001000000100",
			3378 => "0000000011010100001101",
			3379 => "0000001011010100001101",
			3380 => "0000100010110000010100",
			3381 => "0010000110011100010000",
			3382 => "0011011111010000000100",
			3383 => "1111111011010100001101",
			3384 => "0010111011011100001000",
			3385 => "0011100110111100000100",
			3386 => "0000001011010100001101",
			3387 => "0000000011010100001101",
			3388 => "0000000011010100001101",
			3389 => "1111111011010100001101",
			3390 => "0010100001010000001000",
			3391 => "0000011101011000000100",
			3392 => "0000010011010100001101",
			3393 => "0000000011010100001101",
			3394 => "1111111011010100001101",
			3395 => "0010001001000101001000",
			3396 => "0010010100111101000000",
			3397 => "0011101110101000101000",
			3398 => "0011001100110000011000",
			3399 => "0010110100001000010000",
			3400 => "0001101101011100001000",
			3401 => "0000110100001000000100",
			3402 => "0000000011010111010001",
			3403 => "0000010011010111010001",
			3404 => "0011011111011100000100",
			3405 => "1111111011010111010001",
			3406 => "0000000011010111010001",
			3407 => "0001100101011100000100",
			3408 => "0000011011010111010001",
			3409 => "0000001011010111010001",
			3410 => "0001100101011100001100",
			3411 => "0001111110001100001000",
			3412 => "0010111010111100000100",
			3413 => "0000000011010111010001",
			3414 => "0000001011010111010001",
			3415 => "1111111011010111010001",
			3416 => "1111111011010111010001",
			3417 => "0000111000001100010100",
			3418 => "0000000001010100001100",
			3419 => "0010010100111100001000",
			3420 => "0011100010000100000100",
			3421 => "0000001011010111010001",
			3422 => "0000001011010111010001",
			3423 => "1111111011010111010001",
			3424 => "0010011111000000000100",
			3425 => "0000001011010111010001",
			3426 => "1111111011010111010001",
			3427 => "0000010011010111010001",
			3428 => "0000001100000100000100",
			3429 => "1111111011010111010001",
			3430 => "0000001011010111010001",
			3431 => "0010100011101000010000",
			3432 => "0000100110101100001100",
			3433 => "0010110101100100000100",
			3434 => "1111111011010111010001",
			3435 => "0011101100000000000100",
			3436 => "0000001011010111010001",
			3437 => "1111111011010111010001",
			3438 => "0000010011010111010001",
			3439 => "0001011111100100000100",
			3440 => "1111111011010111010001",
			3441 => "0001011000100000000100",
			3442 => "0000000011010111010001",
			3443 => "1111111011010111010001",
			3444 => "0000001011010101000100",
			3445 => "0010000111110100100000",
			3446 => "0000101101000100011100",
			3447 => "0000010111100100010000",
			3448 => "0011100100001000000100",
			3449 => "0000000011011010001101",
			3450 => "0001111110001100001000",
			3451 => "0010010000111100000100",
			3452 => "0000001011011010001101",
			3453 => "0000000011011010001101",
			3454 => "0000000011011010001101",
			3455 => "0011001100110000001000",
			3456 => "0001111110001100000100",
			3457 => "0000000011011010001101",
			3458 => "0000000011011010001101",
			3459 => "1111111011011010001101",
			3460 => "0000001011011010001101",
			3461 => "0011101110010000000100",
			3462 => "1111111011011010001101",
			3463 => "0010100000001000000100",
			3464 => "0000001011011010001101",
			3465 => "0000101100000000010000",
			3466 => "0011010111111100001000",
			3467 => "0001001100010000000100",
			3468 => "1111111011011010001101",
			3469 => "0000000011011010001101",
			3470 => "0011001001110100000100",
			3471 => "1111111011011010001101",
			3472 => "0000000011011010001101",
			3473 => "0010101010100000000100",
			3474 => "0000001011011010001101",
			3475 => "0000010101011100000100",
			3476 => "0000000011011010001101",
			3477 => "1111111011011010001101",
			3478 => "0011010011000000010100",
			3479 => "0010100111110100010000",
			3480 => "0011000100011000000100",
			3481 => "1111111011011010001101",
			3482 => "0000001111001000001000",
			3483 => "0011001000000000000100",
			3484 => "0000000011011010001101",
			3485 => "0000000011011010001101",
			3486 => "0000001011011010001101",
			3487 => "1111111011011010001101",
			3488 => "0011100011110100000100",
			3489 => "0000001011011010001101",
			3490 => "0000000011011010001101",
			3491 => "0001111101100000000100",
			3492 => "1111111011011100011001",
			3493 => "0000000110011100001100",
			3494 => "0000011001011000001000",
			3495 => "0011100100001000000100",
			3496 => "0000000011011100011001",
			3497 => "0000001011011100011001",
			3498 => "0000000011011100011001",
			3499 => "0010110101100100001100",
			3500 => "0010000111110100000100",
			3501 => "0000000011011100011001",
			3502 => "0011111111100100000100",
			3503 => "1111111011011100011001",
			3504 => "0000000011011100011001",
			3505 => "0000111111010100010000",
			3506 => "0010001000100100001000",
			3507 => "0011011001010000000100",
			3508 => "0000000011011100011001",
			3509 => "0000001011011100011001",
			3510 => "0000011001011000000100",
			3511 => "0000000011011100011001",
			3512 => "1111111011011100011001",
			3513 => "0001111111011100001100",
			3514 => "0000010000111100001000",
			3515 => "0000111000001100000100",
			3516 => "0000000011011100011001",
			3517 => "0000001011011100011001",
			3518 => "0000000011011100011001",
			3519 => "0011010011000000001000",
			3520 => "0011001011000000000100",
			3521 => "0000000011011100011001",
			3522 => "1111111011011100011001",
			3523 => "0001110000110100000100",
			3524 => "0000001011011100011001",
			3525 => "0000000011011100011001",
			3526 => "0000001011010101010100",
			3527 => "0010000111110100100000",
			3528 => "0011111100100100011100",
			3529 => "0000010111100100010000",
			3530 => "0000110110100100001000",
			3531 => "0001101111001100000100",
			3532 => "0000001011011111110101",
			3533 => "1111111011011111110101",
			3534 => "0001111110001100000100",
			3535 => "0000001011011111110101",
			3536 => "0000000011011111110101",
			3537 => "0011001100110000001000",
			3538 => "0001111110001100000100",
			3539 => "0000000011011111110101",
			3540 => "0000000011011111110101",
			3541 => "1111111011011111110101",
			3542 => "0000001011011111110101",
			3543 => "0000111001100000001100",
			3544 => "0001110001101000001000",
			3545 => "0011110010000000000100",
			3546 => "1111111011011111110101",
			3547 => "0000000011011111110101",
			3548 => "1111110011011111110101",
			3549 => "0010100000001000001100",
			3550 => "0000111100010000001000",
			3551 => "0001101101111100000100",
			3552 => "0000001011011111110101",
			3553 => "1111111011011111110101",
			3554 => "0000001011011111110101",
			3555 => "0000110111010100010000",
			3556 => "0010110100010000001000",
			3557 => "0011111100000000000100",
			3558 => "0000000011011111110101",
			3559 => "1111111011011111110101",
			3560 => "0011001000000000000100",
			3561 => "0000000011011111110101",
			3562 => "1111110011011111110101",
			3563 => "0011001001110100001000",
			3564 => "0010010100111100000100",
			3565 => "0000001011011111110101",
			3566 => "0000000011011111110101",
			3567 => "1111111011011111110101",
			3568 => "0011010011000000010100",
			3569 => "0010100111110100010000",
			3570 => "0011000100011000000100",
			3571 => "1111111011011111110101",
			3572 => "0010111011011100001000",
			3573 => "0010110101100100000100",
			3574 => "0000000011011111110101",
			3575 => "0000001011011111110101",
			3576 => "0000000011011111110101",
			3577 => "1111111011011111110101",
			3578 => "0001110000110100000100",
			3579 => "0000001011011111110101",
			3580 => "1111111011011111110101",
			3581 => "0010001001000101010000",
			3582 => "0010000111110100100000",
			3583 => "0000101101000100011100",
			3584 => "0000010111100100010000",
			3585 => "0011100100001000000100",
			3586 => "0000000011100011001001",
			3587 => "0001111110001100001000",
			3588 => "0001111101100000000100",
			3589 => "0000000011100011001001",
			3590 => "0000001011100011001001",
			3591 => "0000000011100011001001",
			3592 => "0011001100110000001000",
			3593 => "0001111110001100000100",
			3594 => "0000000011100011001001",
			3595 => "0000000011100011001001",
			3596 => "1111111011100011001001",
			3597 => "0000001011100011001001",
			3598 => "0000101110010000001000",
			3599 => "0010100111101100000100",
			3600 => "1111101011100011001001",
			3601 => "0000000011100011001001",
			3602 => "0010100000001000001100",
			3603 => "0000111100010000001000",
			3604 => "0010011111000000000100",
			3605 => "0000001011100011001001",
			3606 => "1111110011100011001001",
			3607 => "0000001011100011001001",
			3608 => "0000101100000000010000",
			3609 => "0011010111111100001000",
			3610 => "0000110110111100000100",
			3611 => "0000000011100011001001",
			3612 => "0000001011100011001001",
			3613 => "0011001001110100000100",
			3614 => "1111111011100011001001",
			3615 => "0000000011100011001001",
			3616 => "0010110100010000001000",
			3617 => "0010101010100000000100",
			3618 => "0000001011100011001001",
			3619 => "0000000011100011001001",
			3620 => "1111111011100011001001",
			3621 => "0011010011000000010100",
			3622 => "0010100111110100010000",
			3623 => "0000101000100000001100",
			3624 => "0011001000000000000100",
			3625 => "1111111011100011001001",
			3626 => "0011001001001000000100",
			3627 => "0000000011100011001001",
			3628 => "1111111011100011001001",
			3629 => "0000001011100011001001",
			3630 => "1111111011100011001001",
			3631 => "0010011010011000000100",
			3632 => "1111111011100011001001",
			3633 => "0000001011100011001001",
			3634 => "0010100111110100111100",
			3635 => "0010011000010000111000",
			3636 => "0011111111010100110000",
			3637 => "0000000001010100100000",
			3638 => "0001010111100000010000",
			3639 => "0011001011000000001000",
			3640 => "0000110000110100000100",
			3641 => "0000000011100101010101",
			3642 => "0000000011100101010101",
			3643 => "0010000111110100000100",
			3644 => "0000000011100101010101",
			3645 => "1111111011100101010101",
			3646 => "0010001000100100001000",
			3647 => "0000111100000000000100",
			3648 => "0000000011100101010101",
			3649 => "0000001011100101010101",
			3650 => "0011001011000000000100",
			3651 => "0000000011100101010101",
			3652 => "0000000011100101010101",
			3653 => "0000111000001100001100",
			3654 => "0001010111100000001000",
			3655 => "0001010010110100000100",
			3656 => "0000000011100101010101",
			3657 => "0000000011100101010101",
			3658 => "1111111011100101010101",
			3659 => "0000000011100101010101",
			3660 => "0010110101110100000100",
			3661 => "0000001011100101010101",
			3662 => "0000000011100101010101",
			3663 => "0000000011100101010101",
			3664 => "0011010011000000000100",
			3665 => "1111111011100101010101",
			3666 => "0001110000110100000100",
			3667 => "0000000011100101010101",
			3668 => "0000000011100101010101",
			3669 => "0001111101100000000100",
			3670 => "1111111011100111101001",
			3671 => "0010100111101100001000",
			3672 => "0011100100001000000100",
			3673 => "0000000011100111101001",
			3674 => "0000000011100111101001",
			3675 => "0000111010000100100000",
			3676 => "0000111100010000001100",
			3677 => "0010000111110100000100",
			3678 => "0000000011100111101001",
			3679 => "0010100111101100000100",
			3680 => "0000000011100111101001",
			3681 => "1111111011100111101001",
			3682 => "0011010111111100001100",
			3683 => "0000010000111100001000",
			3684 => "0001111111011100000100",
			3685 => "0000000011100111101001",
			3686 => "0000000011100111101001",
			3687 => "0000000011100111101001",
			3688 => "0001111111011100000100",
			3689 => "0000000011100111101001",
			3690 => "0000000011100111101001",
			3691 => "0010110010001000001000",
			3692 => "0011010111111100000100",
			3693 => "0000000011100111101001",
			3694 => "0000000011100111101001",
			3695 => "0001110111010000001100",
			3696 => "0000010101011100001000",
			3697 => "0001111000011000000100",
			3698 => "0000000011100111101001",
			3699 => "0000001011100111101001",
			3700 => "0000000011100111101001",
			3701 => "0011011111101000000100",
			3702 => "0000000011100111101001",
			3703 => "0001111110101100000100",
			3704 => "0000000011100111101001",
			3705 => "0000000011100111101001",
			3706 => "0001111101100000000100",
			3707 => "1111111011101010010101",
			3708 => "0010100111101100010100",
			3709 => "0000010111100100001000",
			3710 => "0011110001111100000100",
			3711 => "0000000011101010010101",
			3712 => "0000000011101010010101",
			3713 => "0000101101000100001000",
			3714 => "0011001100110000000100",
			3715 => "0000000011101010010101",
			3716 => "0000000011101010010101",
			3717 => "0000000011101010010101",
			3718 => "0001010101001000100000",
			3719 => "0011001000000000010100",
			3720 => "0001111000000000000100",
			3721 => "1111111011101010010101",
			3722 => "0011000100011000001000",
			3723 => "0000001100000100000100",
			3724 => "0000000011101010010101",
			3725 => "0000000011101010010101",
			3726 => "0010001000100100000100",
			3727 => "0000000011101010010101",
			3728 => "0000000011101010010101",
			3729 => "0001110001101000000100",
			3730 => "0000000011101010010101",
			3731 => "0011001001110100000100",
			3732 => "1111111011101010010101",
			3733 => "0000000011101010010101",
			3734 => "0000010000111100010100",
			3735 => "0001111111011100010000",
			3736 => "0000111010000100001000",
			3737 => "0011111100000000000100",
			3738 => "0000000011101010010101",
			3739 => "0000000011101010010101",
			3740 => "0010001000100100000100",
			3741 => "0000000011101010010101",
			3742 => "0000001011101010010101",
			3743 => "0000000011101010010101",
			3744 => "0000111111100000001000",
			3745 => "0010110100010000000100",
			3746 => "0000000011101010010101",
			3747 => "0000000011101010010101",
			3748 => "0000000011101010010101",
			3749 => "0001111101100000000100",
			3750 => "1111111011101101000001",
			3751 => "0000000001010100111000",
			3752 => "0000110110111100110000",
			3753 => "0011000100011000011000",
			3754 => "0011111100100100001100",
			3755 => "0011000110000100001000",
			3756 => "0010110100001000000100",
			3757 => "0000000011101101000001",
			3758 => "0000000011101101000001",
			3759 => "0000000011101101000001",
			3760 => "0000010000111100001000",
			3761 => "0011000100011000000100",
			3762 => "0000001011101101000001",
			3763 => "0000000011101101000001",
			3764 => "0000000011101101000001",
			3765 => "0001110001101000001000",
			3766 => "0010011111000000000100",
			3767 => "0000000011101101000001",
			3768 => "0000000011101101000001",
			3769 => "0000011001011000001000",
			3770 => "0010011001100100000100",
			3771 => "0000000011101101000001",
			3772 => "1111111011101101000001",
			3773 => "0000010000111100000100",
			3774 => "0000000011101101000001",
			3775 => "0000000011101101000001",
			3776 => "0001011110000100000100",
			3777 => "0000000011101101000001",
			3778 => "0000001011101101000001",
			3779 => "0000111000001100001000",
			3780 => "0011110000010000000100",
			3781 => "0000000011101101000001",
			3782 => "0000000011101101000001",
			3783 => "0000010101011100001100",
			3784 => "0001111111011100000100",
			3785 => "0000001011101101000001",
			3786 => "0011001001110100000100",
			3787 => "0000000011101101000001",
			3788 => "0000000011101101000001",
			3789 => "0001010111010100000100",
			3790 => "1111111011101101000001",
			3791 => "0000000011101101000001",
			3792 => "0001111101100000000100",
			3793 => "1111111011101111110101",
			3794 => "0010100111101100010000",
			3795 => "0000011101011100001100",
			3796 => "0011110001111100000100",
			3797 => "0000000011101111110101",
			3798 => "0001001001100000000100",
			3799 => "0000000011101111110101",
			3800 => "0000000011101111110101",
			3801 => "0000000011101111110101",
			3802 => "0000110110111100011100",
			3803 => "0001110001101000001100",
			3804 => "0000110110010000000100",
			3805 => "0000000011101111110101",
			3806 => "0001100100110100000100",
			3807 => "0000000011101111110101",
			3808 => "0000000011101111110101",
			3809 => "0001101101111100000100",
			3810 => "0000000011101111110101",
			3811 => "0011000100011000000100",
			3812 => "0000000011101111110101",
			3813 => "0011001001110100000100",
			3814 => "1111111011101111110101",
			3815 => "0000000011101111110101",
			3816 => "0001111000011000011000",
			3817 => "0011110111011000001100",
			3818 => "0001110001101000001000",
			3819 => "0010010100111100000100",
			3820 => "0000000011101111110101",
			3821 => "0000000011101111110101",
			3822 => "0000000011101111110101",
			3823 => "0011010111111100000100",
			3824 => "0000000011101111110101",
			3825 => "0011011110010000000100",
			3826 => "1111111011101111110101",
			3827 => "0000000011101111110101",
			3828 => "0000010000111100001100",
			3829 => "0001111111011100001000",
			3830 => "0011010100101000000100",
			3831 => "0000000011101111110101",
			3832 => "0000000011101111110101",
			3833 => "0000000011101111110101",
			3834 => "0000111111100000000100",
			3835 => "0000000011101111110101",
			3836 => "0000000011101111110101",
			3837 => "0001111101100000000100",
			3838 => "1111111011110010011011",
			3839 => "0010100001010001001100",
			3840 => "0001111000011000110000",
			3841 => "0010100111101100010100",
			3842 => "0000101101000100010000",
			3843 => "0000010110101000001000",
			3844 => "0011001000111000000100",
			3845 => "0000001011110010011011",
			3846 => "0000000011110010011011",
			3847 => "0011001100110000000100",
			3848 => "0000000011110010011011",
			3849 => "0000000011110010011011",
			3850 => "0000001011110010011011",
			3851 => "0000111100010000001100",
			3852 => "0000000110011100000100",
			3853 => "0000000011110010011011",
			3854 => "0001110001101000000100",
			3855 => "1111111011110010011011",
			3856 => "0000000011110010011011",
			3857 => "0010100000001000001000",
			3858 => "0010010100111100000100",
			3859 => "0000001011110010011011",
			3860 => "0000000011110010011011",
			3861 => "0001101101111100000100",
			3862 => "0000000011110010011011",
			3863 => "0000000011110010011011",
			3864 => "0001111111011100001100",
			3865 => "0000010000111100001000",
			3866 => "0000100110010000000100",
			3867 => "0000000011110010011011",
			3868 => "0000001011110010011011",
			3869 => "0000000011110010011011",
			3870 => "0011101011111000000100",
			3871 => "0000000011110010011011",
			3872 => "0000011101111100001000",
			3873 => "0010001001101000000100",
			3874 => "0000000011110010011011",
			3875 => "0000000011110010011011",
			3876 => "0000000011110010011011",
			3877 => "0000000011110010011011",
			3878 => "0000000011110010011101",
			3879 => "0000000011110010100001",
			3880 => "0000000011110010100101",
			3881 => "0000000011110010101001",
			3882 => "0000000011110010101101",
			3883 => "0000000011110010110001",
			3884 => "0000000011110010110101",
			3885 => "0000000011110010111001",
			3886 => "0010001001111100001000",
			3887 => "0011110001111100000100",
			3888 => "0000000011110011010101",
			3889 => "0000000011110011010101",
			3890 => "0011111100010100000100",
			3891 => "0000000011110011010101",
			3892 => "0000000011110011010101",
			3893 => "0000110111010100001000",
			3894 => "0000111101010100000100",
			3895 => "0000000011110011110001",
			3896 => "0000000011110011110001",
			3897 => "0000110010100100000100",
			3898 => "0000000011110011110001",
			3899 => "0000000011110011110001",
			3900 => "0000010110101000000100",
			3901 => "0000000011110100001101",
			3902 => "0011011010001000001000",
			3903 => "0001010101001000000100",
			3904 => "0000000011110100001101",
			3905 => "0000000011110100001101",
			3906 => "0000000011110100001101",
			3907 => "0000110111010100001100",
			3908 => "0010010000111100000100",
			3909 => "0000000011110100101001",
			3910 => "0011011010001000000100",
			3911 => "0000000011110100101001",
			3912 => "0000000011110100101001",
			3913 => "0000000011110100101001",
			3914 => "0001011111010000001100",
			3915 => "0001110001101000000100",
			3916 => "0000000011110101001101",
			3917 => "0001011101000100000100",
			3918 => "0000000011110101001101",
			3919 => "0000000011110101001101",
			3920 => "0001110001001000000100",
			3921 => "0000000011110101001101",
			3922 => "0000000011110101001101",
			3923 => "0010010101011100001100",
			3924 => "0011100100001000000100",
			3925 => "0000000011110101110001",
			3926 => "0000001100011100000100",
			3927 => "0000000011110101110001",
			3928 => "0000000011110101110001",
			3929 => "0001101101111100000100",
			3930 => "0000000011110101110001",
			3931 => "0000000011110101110001",
			3932 => "0010110101100100001100",
			3933 => "0011001100110000000100",
			3934 => "0000000011110110011101",
			3935 => "0011001000000000000100",
			3936 => "0000000011110110011101",
			3937 => "0000000011110110011101",
			3938 => "0000010000111100001000",
			3939 => "0001110111010000000100",
			3940 => "0000000011110110011101",
			3941 => "0000000011110110011101",
			3942 => "0000000011110110011101",
			3943 => "0010100000001000001100",
			3944 => "0000000010101100000100",
			3945 => "0000000011110111001001",
			3946 => "0000000001110000000100",
			3947 => "0000000011110111001001",
			3948 => "0000000011110111001001",
			3949 => "0010100110011000001000",
			3950 => "0000000001010100000100",
			3951 => "0000000011110111001001",
			3952 => "0000000011110111001001",
			3953 => "0000000011110111001001",
			3954 => "0010110100010000010000",
			3955 => "0010111000011000000100",
			3956 => "0000000011110111101101",
			3957 => "0001100100110100001000",
			3958 => "0000010000111100000100",
			3959 => "0000000011110111101101",
			3960 => "0000000011110111101101",
			3961 => "0000000011110111101101",
			3962 => "0000000011110111101101",
			3963 => "0001001111100100010000",
			3964 => "0000101100010000000100",
			3965 => "0000000011111000010001",
			3966 => "0000101010000100001000",
			3967 => "0010001001000100000100",
			3968 => "0000000011111000010001",
			3969 => "0000000011111000010001",
			3970 => "0000000011111000010001",
			3971 => "0000000011111000010001",
			3972 => "0001111000011000010000",
			3973 => "0001110001101000000100",
			3974 => "0000000011111000110101",
			3975 => "0001101101111100000100",
			3976 => "0000000011111000110101",
			3977 => "0011011001010000000100",
			3978 => "0000000011111000110101",
			3979 => "0000000011111000110101",
			3980 => "0000000011111000110101",
			3981 => "0001100100110100010000",
			3982 => "0010101010100000001100",
			3983 => "0001100111101000000100",
			3984 => "0000000011111001100001",
			3985 => "0010100000001000000100",
			3986 => "0000000011111001100001",
			3987 => "0000000011111001100001",
			3988 => "0000000011111001100001",
			3989 => "0010100000001000000100",
			3990 => "0000000011111001100001",
			3991 => "0000000011111001100001",
			3992 => "0010001001111100001100",
			3993 => "0010010000111100001000",
			3994 => "0011110001111100000100",
			3995 => "0000000011111010010101",
			3996 => "0000000011111010010101",
			3997 => "0000000011111010010101",
			3998 => "0010110101100100000100",
			3999 => "0000000011111010010101",
			4000 => "0010110100010000000100",
			4001 => "0000000011111010010101",
			4002 => "0010110111111100000100",
			4003 => "0000000011111010010101",
			4004 => "0000000011111010010101",
			4005 => "0010100000001000010000",
			4006 => "0010100100110100000100",
			4007 => "0000000011111011001001",
			4008 => "0000000001010100001000",
			4009 => "0010100111101100000100",
			4010 => "0000000011111011001001",
			4011 => "0000000011111011001001",
			4012 => "0000000011111011001001",
			4013 => "0000000101000100000100",
			4014 => "0000000011111011001001",
			4015 => "0010100110011000000100",
			4016 => "0000000011111011001001",
			4017 => "0000000011111011001001",
			4018 => "0000111110110100001100",
			4019 => "0010010000111100000100",
			4020 => "0000000011111011111101",
			4021 => "0000010110101000000100",
			4022 => "0000000011111011111101",
			4023 => "0000000011111011111101",
			4024 => "0000100111010100001100",
			4025 => "0001111111011100001000",
			4026 => "0000010000111100000100",
			4027 => "0000000011111011111101",
			4028 => "0000000011111011111101",
			4029 => "0000000011111011111101",
			4030 => "0000000011111011111101",
			4031 => "0010001001111100001100",
			4032 => "0000010110101000001000",
			4033 => "0011100100001000000100",
			4034 => "0000000011111100111001",
			4035 => "0000000011111100111001",
			4036 => "0000000011111100111001",
			4037 => "0000011001011000001100",
			4038 => "0001010101001000001000",
			4039 => "0011110000010000000100",
			4040 => "0000000011111100111001",
			4041 => "0000000011111100111001",
			4042 => "0000000011111100111001",
			4043 => "0000010000111100000100",
			4044 => "0000000011111100111001",
			4045 => "0000000011111100111001",
			4046 => "0010011100011000001000",
			4047 => "0011001100110000000100",
			4048 => "0000000011111101101101",
			4049 => "0000000011111101101101",
			4050 => "0010011111000000010000",
			4051 => "0011001000011000001100",
			4052 => "0000011111001100000100",
			4053 => "0000000011111101101101",
			4054 => "0011000110000100000100",
			4055 => "0000000011111101101101",
			4056 => "0000000011111101101101",
			4057 => "0000000011111101101101",
			4058 => "0000000011111101101101",
			4059 => "0011101110101000001000",
			4060 => "0010001001111100000100",
			4061 => "0000000011111110100001",
			4062 => "0000000011111110100001",
			4063 => "0000010101011100010000",
			4064 => "0001110111010000001100",
			4065 => "0001101010011000001000",
			4066 => "0011000110000100000100",
			4067 => "0000000011111110100001",
			4068 => "0000000011111110100001",
			4069 => "0000000011111110100001",
			4070 => "0000000011111110100001",
			4071 => "0000000011111110100001",
			4072 => "0000010110101000000100",
			4073 => "0000000011111111001101",
			4074 => "0011011010001000010000",
			4075 => "0011001100110000000100",
			4076 => "0000000011111111001101",
			4077 => "0011001001001000001000",
			4078 => "0001111111011100000100",
			4079 => "0000000011111111001101",
			4080 => "0000000011111111001101",
			4081 => "0000000011111111001101",
			4082 => "0000000011111111001101",
			4083 => "0000111110110100001100",
			4084 => "0011011010011100000100",
			4085 => "0000000100000000001001",
			4086 => "0000010110101000000100",
			4087 => "0000000100000000001001",
			4088 => "0000000100000000001001",
			4089 => "0000011111001100000100",
			4090 => "0000000100000000001001",
			4091 => "0010110101110100001100",
			4092 => "0000010000111100001000",
			4093 => "0001101011001100000100",
			4094 => "0000000100000000001001",
			4095 => "0000000100000000001001",
			4096 => "0000000100000000001001",
			4097 => "0000000100000000001001",
			4098 => "0010110101100100010000",
			4099 => "0000100000110100000100",
			4100 => "0000000100000001001101",
			4101 => "0011001000000000001000",
			4102 => "0001111000011000000100",
			4103 => "0000000100000001001101",
			4104 => "0000000100000001001101",
			4105 => "0000000100000001001101",
			4106 => "0001101101111100000100",
			4107 => "0000000100000001001101",
			4108 => "0000011101111100001100",
			4109 => "0001011100100100000100",
			4110 => "0000000100000001001101",
			4111 => "0001100101010000000100",
			4112 => "0000000100000001001101",
			4113 => "0000000100000001001101",
			4114 => "0000000100000001001101",
			4115 => "0000111100010000010100",
			4116 => "0010010000111100001100",
			4117 => "0000000011101000001000",
			4118 => "0011100100001000000100",
			4119 => "0000000100000010011001",
			4120 => "0000000100000010011001",
			4121 => "0000000100000010011001",
			4122 => "0000010110101000000100",
			4123 => "0000000100000010011001",
			4124 => "0000000100000010011001",
			4125 => "0000011111001100000100",
			4126 => "0000000100000010011001",
			4127 => "0000011101111100001100",
			4128 => "0001011110101000000100",
			4129 => "0000000100000010011001",
			4130 => "0010100001010000000100",
			4131 => "0000000100000010011001",
			4132 => "0000000100000010011001",
			4133 => "0000000100000010011001",
			4134 => "0011101010001000010100",
			4135 => "0010100111101100010000",
			4136 => "0000010110101000001000",
			4137 => "0011100100001000000100",
			4138 => "0000000100000011100101",
			4139 => "0000000100000011100101",
			4140 => "0001100000111100000100",
			4141 => "0000000100000011100101",
			4142 => "0000000100000011100101",
			4143 => "0000000100000011100101",
			4144 => "0010010100111100010000",
			4145 => "0001111000011000001100",
			4146 => "0001111011000000000100",
			4147 => "0000000100000011100101",
			4148 => "0010110100000100000100",
			4149 => "0000000100000011100101",
			4150 => "0000000100000011100101",
			4151 => "0000000100000011100101",
			4152 => "0000000100000011100101",
			4153 => "0000111010000100011100",
			4154 => "0011001100110000010000",
			4155 => "0011100100001000000100",
			4156 => "0000000100000100111001",
			4157 => "0011000100000000000100",
			4158 => "0000000100000100111001",
			4159 => "0011100101110000000100",
			4160 => "0000000100000100111001",
			4161 => "0000000100000100111001",
			4162 => "0011001001110100001000",
			4163 => "0011101100010000000100",
			4164 => "0000000100000100111001",
			4165 => "0000000100000100111001",
			4166 => "0000000100000100111001",
			4167 => "0011001011011100001100",
			4168 => "0011000111001000000100",
			4169 => "0000000100000100111001",
			4170 => "0011100000010100000100",
			4171 => "0000000100000100111001",
			4172 => "0000000100000100111001",
			4173 => "0000000100000100111001",
			4174 => "0001110110000100001100",
			4175 => "0011111010111100000100",
			4176 => "0000000100000101111101",
			4177 => "0001011010011100000100",
			4178 => "0000000100000101111101",
			4179 => "0000000100000101111101",
			4180 => "0010011111000000010100",
			4181 => "0001110111010000010000",
			4182 => "0000001100000100001100",
			4183 => "0001011111010000001000",
			4184 => "0011111001001000000100",
			4185 => "0000000100000101111101",
			4186 => "0000000100000101111101",
			4187 => "0000000100000101111101",
			4188 => "0000000100000101111101",
			4189 => "0000000100000101111101",
			4190 => "0000000100000101111101",
			4191 => "0000011111001100010100",
			4192 => "0011001100110000010000",
			4193 => "0001111101100000000100",
			4194 => "0000000100000111001001",
			4195 => "0011100100001000000100",
			4196 => "0000000100000111001001",
			4197 => "0000000101000100000100",
			4198 => "0000000100000111001001",
			4199 => "0000000100000111001001",
			4200 => "0000000100000111001001",
			4201 => "0000010000111100010000",
			4202 => "0001111111011100001100",
			4203 => "0011010010110100000100",
			4204 => "0000000100000111001001",
			4205 => "0011000000001100000100",
			4206 => "0000000100000111001001",
			4207 => "0000000100000111001001",
			4208 => "0000000100000111001001",
			4209 => "0000000100000111001001",
			4210 => "0010110010001000011100",
			4211 => "0000000110011100010000",
			4212 => "0010010000111100001000",
			4213 => "0011100100001000000100",
			4214 => "0000000100001000100101",
			4215 => "0000000100001000100101",
			4216 => "0011100101100100000100",
			4217 => "0000000100001000100101",
			4218 => "0000000100001000100101",
			4219 => "0000111100000000001000",
			4220 => "0001011100100100000100",
			4221 => "0000000100001000100101",
			4222 => "0000000100001000100101",
			4223 => "0000000100001000100101",
			4224 => "0001110111010000010000",
			4225 => "0000010101011100001100",
			4226 => "0011001011000000000100",
			4227 => "0000000100001000100101",
			4228 => "0011001001110100000100",
			4229 => "0000000100001000100101",
			4230 => "0000000100001000100101",
			4231 => "0000000100001000100101",
			4232 => "0000000100001000100101",
			4233 => "0000010000111100011100",
			4234 => "0011101110101000001000",
			4235 => "0001100001000100000100",
			4236 => "0000000100001001100001",
			4237 => "0000000100001001100001",
			4238 => "0001111000011000010000",
			4239 => "0010010100111100001100",
			4240 => "0011011001011100001000",
			4241 => "0001101100011000000100",
			4242 => "0000000100001001100001",
			4243 => "0000000100001001100001",
			4244 => "0000000100001001100001",
			4245 => "0000000100001001100001",
			4246 => "0000000100001001100001",
			4247 => "0000000100001001100001",
			4248 => "0001010101001000010000",
			4249 => "0000100000110100000100",
			4250 => "0000000100001010101101",
			4251 => "0000011001011000001000",
			4252 => "0011001001110100000100",
			4253 => "0000000100001010101101",
			4254 => "0000000100001010101101",
			4255 => "0000000100001010101101",
			4256 => "0010110100010000000100",
			4257 => "0000000100001010101101",
			4258 => "0001100101010000010000",
			4259 => "0011001011000000000100",
			4260 => "0000000100001010101101",
			4261 => "0000011101111100001000",
			4262 => "0000011101011100000100",
			4263 => "0000000100001010101101",
			4264 => "0000000100001010101101",
			4265 => "0000000100001010101101",
			4266 => "0000000100001010101101",
			4267 => "0011001100110000010100",
			4268 => "0011100100001000000100",
			4269 => "0000000100001100001001",
			4270 => "0010011101111100001100",
			4271 => "0011000100000000000100",
			4272 => "0000000100001100001001",
			4273 => "0010011011101000000100",
			4274 => "0000000100001100001001",
			4275 => "0000000100001100001001",
			4276 => "0000000100001100001001",
			4277 => "0000111010000100001100",
			4278 => "0011001001110100001000",
			4279 => "0011101100010000000100",
			4280 => "0000000100001100001001",
			4281 => "0000000100001100001001",
			4282 => "0000000100001100001001",
			4283 => "0010011000010000001100",
			4284 => "0010011100011000000100",
			4285 => "0000000100001100001001",
			4286 => "0011001000011000000100",
			4287 => "0000000100001100001001",
			4288 => "0000000100001100001001",
			4289 => "0000000100001100001001",
			4290 => "0000111010000100011100",
			4291 => "0010100000001000001100",
			4292 => "0000101110010000001000",
			4293 => "0001011110101000000100",
			4294 => "0000000100001101110101",
			4295 => "0000000100001101110101",
			4296 => "0000000100001101110101",
			4297 => "0011111111010100001100",
			4298 => "0000000101000100000100",
			4299 => "0000000100001101110101",
			4300 => "0001101101111100000100",
			4301 => "0000000100001101110101",
			4302 => "0000000100001101110101",
			4303 => "0000000100001101110101",
			4304 => "0011001001001000010000",
			4305 => "0000001011010100001100",
			4306 => "0001111000011000000100",
			4307 => "0000000100001101110101",
			4308 => "0000010101011100000100",
			4309 => "0000000100001101110101",
			4310 => "0000000100001101110101",
			4311 => "0000000100001101110101",
			4312 => "0010110111111100001000",
			4313 => "0001110001101000000100",
			4314 => "0000000100001101110101",
			4315 => "0000000100001101110101",
			4316 => "0000000100001101110101",
			4317 => "0001011111010000100100",
			4318 => "0000000101000100010100",
			4319 => "0011111001001000001000",
			4320 => "0000011001111000000100",
			4321 => "0000000100001111100001",
			4322 => "0000000100001111100001",
			4323 => "0000011101101000001000",
			4324 => "0010110100001000000100",
			4325 => "0000000100001111100001",
			4326 => "0000000100001111100001",
			4327 => "0000000100001111100001",
			4328 => "0011011010001000001100",
			4329 => "0001011100100100000100",
			4330 => "0000000100001111100001",
			4331 => "0011010010011100000100",
			4332 => "0000000100001111100001",
			4333 => "0000000100001111100001",
			4334 => "0000000100001111100001",
			4335 => "0010100001010000010000",
			4336 => "0010110010001000000100",
			4337 => "0000000100001111100001",
			4338 => "0001111000011000000100",
			4339 => "0000000100001111100001",
			4340 => "0010011010100000000100",
			4341 => "0000000100001111100001",
			4342 => "0000000100001111100001",
			4343 => "0000000100001111100001",
			4344 => "0001011100100100011100",
			4345 => "0000000110011100001100",
			4346 => "0011111010011100000100",
			4347 => "0000000100010001000101",
			4348 => "0011111110101000000100",
			4349 => "0000000100010001000101",
			4350 => "0000000100010001000101",
			4351 => "0011111100010000001100",
			4352 => "0011010101110000001000",
			4353 => "0010000111110100000100",
			4354 => "0000000100010001000101",
			4355 => "0000000100010001000101",
			4356 => "0000000100010001000101",
			4357 => "0000000100010001000101",
			4358 => "0010100001010000010100",
			4359 => "0000011101111100010000",
			4360 => "0011000111001000000100",
			4361 => "0000000100010001000101",
			4362 => "0000111100010000000100",
			4363 => "0000000100010001000101",
			4364 => "0001101000010000000100",
			4365 => "0000000100010001000101",
			4366 => "0000000100010001000101",
			4367 => "0000000100010001000101",
			4368 => "0000000100010001000101",
			4369 => "0001011111010000011100",
			4370 => "0011001011000000010000",
			4371 => "0000001100000100001100",
			4372 => "0010101101011000000100",
			4373 => "0000000100010010101001",
			4374 => "0011000011011100000100",
			4375 => "0000000100010010101001",
			4376 => "0000000100010010101001",
			4377 => "0000000100010010101001",
			4378 => "0010000111110100000100",
			4379 => "0000000100010010101001",
			4380 => "0000001011010100000100",
			4381 => "0000000100010010101001",
			4382 => "0000000100010010101001",
			4383 => "0001100101010000010100",
			4384 => "0011001011000000000100",
			4385 => "0000000100010010101001",
			4386 => "0010011010100000001100",
			4387 => "0010100001010000001000",
			4388 => "0010110010001000000100",
			4389 => "0000000100010010101001",
			4390 => "0000000100010010101001",
			4391 => "0000000100010010101001",
			4392 => "0000000100010010101001",
			4393 => "0000000100010010101001",
			4394 => "0001111000000000011100",
			4395 => "0000100000110100010100",
			4396 => "0000010110101000010000",
			4397 => "0000100100001000000100",
			4398 => "0000000100010100011101",
			4399 => "0011000100000000000100",
			4400 => "0000000100010100011101",
			4401 => "0001000111001000000100",
			4402 => "0000000100010100011101",
			4403 => "0000000100010100011101",
			4404 => "0000000100010100011101",
			4405 => "0011000100011000000100",
			4406 => "0000000100010100011101",
			4407 => "0000000100010100011101",
			4408 => "0000111111010100010100",
			4409 => "0011001011000000001000",
			4410 => "0000011001011000000100",
			4411 => "0000000100010100011101",
			4412 => "0000000100010100011101",
			4413 => "0010000111110100000100",
			4414 => "0000000100010100011101",
			4415 => "0001110110100100000100",
			4416 => "0000000100010100011101",
			4417 => "0000000100010100011101",
			4418 => "0010010100111100001000",
			4419 => "0001111111011100000100",
			4420 => "0000000100010100011101",
			4421 => "0000000100010100011101",
			4422 => "0000000100010100011101",
			4423 => "0000111000011000001000",
			4424 => "0001101101011100000100",
			4425 => "0000000100010101100001",
			4426 => "0000000100010101100001",
			4427 => "0010100000001000011000",
			4428 => "0001100100110100010100",
			4429 => "0001100000111100000100",
			4430 => "0000000100010101100001",
			4431 => "0010110100001000000100",
			4432 => "0000000100010101100001",
			4433 => "0011111010011100000100",
			4434 => "0000000100010101100001",
			4435 => "0000010000111100000100",
			4436 => "0000000100010101100001",
			4437 => "0000000100010101100001",
			4438 => "0000000100010101100001",
			4439 => "0000000100010101100001",
			4440 => "0010100000001000010100",
			4441 => "0010010101011100001100",
			4442 => "0000010110101000001000",
			4443 => "0011100100001000000100",
			4444 => "0000000100010111001101",
			4445 => "0000000100010111001101",
			4446 => "0000000100010111001101",
			4447 => "0000101101000100000100",
			4448 => "0000000100010111001101",
			4449 => "0000000100010111001101",
			4450 => "0000111010000100001100",
			4451 => "0000010000111100001000",
			4452 => "0000101010000100000100",
			4453 => "0000000100010111001101",
			4454 => "0000000100010111001101",
			4455 => "0000000100010111001101",
			4456 => "0011001011000000000100",
			4457 => "0000000100010111001101",
			4458 => "0000011101111100010000",
			4459 => "0001110001101000000100",
			4460 => "0000000100010111001101",
			4461 => "0000011111001100000100",
			4462 => "0000000100010111001101",
			4463 => "0001010010011100000100",
			4464 => "0000000100010111001101",
			4465 => "0000000100010111001101",
			4466 => "0000000100010111001101",
			4467 => "0001011111010000100000",
			4468 => "0000000101000100011000",
			4469 => "0011001000000000010100",
			4470 => "0010101101011000000100",
			4471 => "0000000100011000110001",
			4472 => "0011000011011100000100",
			4473 => "0000000100011000110001",
			4474 => "0010100000001000001000",
			4475 => "0011001011000000000100",
			4476 => "0000000100011000110001",
			4477 => "0000000100011000110001",
			4478 => "0000000100011000110001",
			4479 => "0000000100011000110001",
			4480 => "0010100000001000000100",
			4481 => "0000000100011000110001",
			4482 => "0000000100011000110001",
			4483 => "0010100001010000010000",
			4484 => "0011001011000000000100",
			4485 => "0000000100011000110001",
			4486 => "0000011101111100001000",
			4487 => "0001111000011000000100",
			4488 => "0000000100011000110001",
			4489 => "0000000100011000110001",
			4490 => "0000000100011000110001",
			4491 => "0000000100011000110001",
			4492 => "0000000001010100101100",
			4493 => "0011101000011000001100",
			4494 => "0000010110101000001000",
			4495 => "0011100100001000000100",
			4496 => "0000000100011010010101",
			4497 => "0000000100011010010101",
			4498 => "1111111100011010010101",
			4499 => "0011001000000000010100",
			4500 => "0001100100110100010000",
			4501 => "0001100000111100000100",
			4502 => "0000000100011010010101",
			4503 => "0010010100111100001000",
			4504 => "0011100101100100000100",
			4505 => "0000000100011010010101",
			4506 => "0000000100011010010101",
			4507 => "0000000100011010010101",
			4508 => "0000000100011010010101",
			4509 => "0000101110110100000100",
			4510 => "0000000100011010010101",
			4511 => "0000101100010000000100",
			4512 => "0000000100011010010101",
			4513 => "0000000100011010010101",
			4514 => "0001101101111100000100",
			4515 => "0000000100011010010101",
			4516 => "0000000100011010010101",
			4517 => "0000111000001100101100",
			4518 => "0010001000100100100100",
			4519 => "0011001100110000010000",
			4520 => "0000010111100100001100",
			4521 => "0011110001111100000100",
			4522 => "0000000100011100001001",
			4523 => "0000010010001100000100",
			4524 => "0000000100011100001001",
			4525 => "0000000100011100001001",
			4526 => "0000000100011100001001",
			4527 => "0000111100010000001100",
			4528 => "0000010110101000000100",
			4529 => "0000000100011100001001",
			4530 => "0010000100101100000100",
			4531 => "0000000100011100001001",
			4532 => "0000000100011100001001",
			4533 => "0000011001011000000100",
			4534 => "0000000100011100001001",
			4535 => "0000000100011100001001",
			4536 => "0011111111100100000100",
			4537 => "0000000100011100001001",
			4538 => "0000000100011100001001",
			4539 => "0001101000010000001100",
			4540 => "0011001011000000000100",
			4541 => "0000000100011100001001",
			4542 => "0000011101111100000100",
			4543 => "0000000100011100001001",
			4544 => "0000000100011100001001",
			4545 => "0000000100011100001001",
			4546 => "0001101001011000010000",
			4547 => "0000010110101000001100",
			4548 => "0011100100001000000100",
			4549 => "0000000100011110000101",
			4550 => "0001111101100000000100",
			4551 => "0000000100011110000101",
			4552 => "0000000100011110000101",
			4553 => "0000000100011110000101",
			4554 => "0001010101001000011100",
			4555 => "0010000111110100000100",
			4556 => "0000000100011110000101",
			4557 => "0000111100010000001000",
			4558 => "0010100111101100000100",
			4559 => "0000000100011110000101",
			4560 => "0000000100011110000101",
			4561 => "0010100000001000000100",
			4562 => "0000000100011110000101",
			4563 => "0011101001100000000100",
			4564 => "0000000100011110000101",
			4565 => "0000101000100000000100",
			4566 => "0000000100011110000101",
			4567 => "0000000100011110000101",
			4568 => "0001111000011000001100",
			4569 => "0000010000111100001000",
			4570 => "0010001000100100000100",
			4571 => "0000000100011110000101",
			4572 => "0000000100011110000101",
			4573 => "0000000100011110000101",
			4574 => "0011010110010000000100",
			4575 => "0000000100011110000101",
			4576 => "0000000100011110000101",
			4577 => "0010110010001000110000",
			4578 => "0010100111101100100000",
			4579 => "0000001010100100010000",
			4580 => "0000010110101000001100",
			4581 => "0000100100001000000100",
			4582 => "0000000100100000001001",
			4583 => "0001111101100000000100",
			4584 => "0000000100100000001001",
			4585 => "0000000100100000001001",
			4586 => "0000000100100000001001",
			4587 => "0010100100111100000100",
			4588 => "0000000100100000001001",
			4589 => "0011110010001000000100",
			4590 => "0000000100100000001001",
			4591 => "0001101101111100000100",
			4592 => "0000000100100000001001",
			4593 => "0000000100100000001001",
			4594 => "0000111100000000001100",
			4595 => "0000000110011100000100",
			4596 => "0000000100100000001001",
			4597 => "0001011100100100000100",
			4598 => "0000000100100000001001",
			4599 => "0000000100100000001001",
			4600 => "0000000100100000001001",
			4601 => "0001110111010000010000",
			4602 => "0000010101011100001100",
			4603 => "0011001011000000000100",
			4604 => "0000000100100000001001",
			4605 => "0011001001110100000100",
			4606 => "0000000100100000001001",
			4607 => "0000000100100000001001",
			4608 => "0000000100100000001001",
			4609 => "0000000100100000001001",
			4610 => "0000000001010100110100",
			4611 => "0001011100100100100100",
			4612 => "0000011101011100010000",
			4613 => "0011000100011000001100",
			4614 => "0000100100001000000100",
			4615 => "0000000100100010000101",
			4616 => "0010100111101100000100",
			4617 => "0000000100100010000101",
			4618 => "0000000100100010000101",
			4619 => "0000000100100010000101",
			4620 => "0010011101011000000100",
			4621 => "0000000100100010000101",
			4622 => "0000101001100000001100",
			4623 => "0011000100001000000100",
			4624 => "0000000100100010000101",
			4625 => "0011001000000000000100",
			4626 => "0000000100100010000101",
			4627 => "0000000100100010000101",
			4628 => "0000000100100010000101",
			4629 => "0001011111010000001100",
			4630 => "0011000100011000000100",
			4631 => "0000000100100010000101",
			4632 => "0010010100111100000100",
			4633 => "0000000100100010000101",
			4634 => "0000000100100010000101",
			4635 => "0000000100100010000101",
			4636 => "0011110110001100001000",
			4637 => "0010100000001000000100",
			4638 => "0000000100100010000101",
			4639 => "0000000100100010000101",
			4640 => "0000000100100010000101",
			4641 => "0001010111100000110100",
			4642 => "0001101101111100100000",
			4643 => "0011100110100100001000",
			4644 => "0001101111001100000100",
			4645 => "0000000100100100101001",
			4646 => "0000000100100100101001",
			4647 => "0011001110001100010000",
			4648 => "0010110100001000000100",
			4649 => "0000000100100100101001",
			4650 => "0011111010011100000100",
			4651 => "0000000100100100101001",
			4652 => "0001111100101000000100",
			4653 => "0000000100100100101001",
			4654 => "0000000100100100101001",
			4655 => "0001011001010100000100",
			4656 => "0000000100100100101001",
			4657 => "0000000100100100101001",
			4658 => "0000111100000000010000",
			4659 => "0000001100011100000100",
			4660 => "0000000100100100101001",
			4661 => "0001011100100100001000",
			4662 => "0011010010011100000100",
			4663 => "0000000100100100101001",
			4664 => "0000000100100100101001",
			4665 => "0000000100100100101001",
			4666 => "0000000100100100101001",
			4667 => "0001101101111100001100",
			4668 => "0000101110110100000100",
			4669 => "0000000100100100101001",
			4670 => "0010011111000000000100",
			4671 => "0000000100100100101001",
			4672 => "0000000100100100101001",
			4673 => "0001111000011000001000",
			4674 => "0010010100111100000100",
			4675 => "0000000100100100101001",
			4676 => "0000000100100100101001",
			4677 => "0000111000100000000100",
			4678 => "0000000100100100101001",
			4679 => "0000110010100100000100",
			4680 => "0000000100100100101001",
			4681 => "0000000100100100101001",
			4682 => "0011101010001000011100",
			4683 => "0000001100011100011000",
			4684 => "0010100100111100010000",
			4685 => "0001010001101000001100",
			4686 => "0000110110100100000100",
			4687 => "0000000100100111000101",
			4688 => "0001100000111100000100",
			4689 => "0000000100100111000101",
			4690 => "0000000100100111000101",
			4691 => "0000000100100111000101",
			4692 => "0011110010001000000100",
			4693 => "0000000100100111000101",
			4694 => "0000000100100111000101",
			4695 => "1111111100100111000101",
			4696 => "0010010100111100100100",
			4697 => "0011001000000000001100",
			4698 => "0001100100110100001000",
			4699 => "0000111110110100000100",
			4700 => "0000000100100111000101",
			4701 => "0000000100100111000101",
			4702 => "0000000100100111000101",
			4703 => "0011101100010000001100",
			4704 => "0000000101000100000100",
			4705 => "0000000100100111000101",
			4706 => "0010110101110100000100",
			4707 => "0000000100100111000101",
			4708 => "0000000100100111000101",
			4709 => "0010011101011000000100",
			4710 => "0000000100100111000101",
			4711 => "0011001001110100000100",
			4712 => "0000000100100111000101",
			4713 => "0000000100100111000101",
			4714 => "0011011010001000000100",
			4715 => "0000000100100111000101",
			4716 => "0000111000001100000100",
			4717 => "0000000100100111000101",
			4718 => "0001011111010000000100",
			4719 => "0000000100100111000101",
			4720 => "0000000100100111000101",
			4721 => "0010000110011100110100",
			4722 => "0000010000111100101100",
			4723 => "0000110111010100100000",
			4724 => "0000000001010100010100",
			4725 => "0011111100000000010000",
			4726 => "0000111110110100001000",
			4727 => "0010000111110100000100",
			4728 => "0000000100101001000001",
			4729 => "0000000100101001000001",
			4730 => "0010010100111100000100",
			4731 => "0000001100101001000001",
			4732 => "0000000100101001000001",
			4733 => "0000000100101001000001",
			4734 => "0000011001011000001000",
			4735 => "0010110100000100000100",
			4736 => "0000000100101001000001",
			4737 => "0000000100101001000001",
			4738 => "0000000100101001000001",
			4739 => "0000101100000000000100",
			4740 => "0000000100101001000001",
			4741 => "0001111111011100000100",
			4742 => "0000001100101001000001",
			4743 => "0000000100101001000001",
			4744 => "0010010100111100000100",
			4745 => "0000000100101001000001",
			4746 => "0000000100101001000001",
			4747 => "0011010011000000000100",
			4748 => "1111111100101001000001",
			4749 => "0001110000110100000100",
			4750 => "0000000100101001000001",
			4751 => "0000000100101001000001",
			4752 => "0001111000011000111000",
			4753 => "0010110010001000101100",
			4754 => "0010100111101100011000",
			4755 => "0011000110000100010000",
			4756 => "0000001010110000001100",
			4757 => "0011100100001000000100",
			4758 => "0000000100101011001101",
			4759 => "0001111101100000000100",
			4760 => "0000000100101011001101",
			4761 => "0000000100101011001101",
			4762 => "0000000100101011001101",
			4763 => "0000101100100100000100",
			4764 => "0000000100101011001101",
			4765 => "0000000100101011001101",
			4766 => "0001010001000000010000",
			4767 => "0011111111100100001100",
			4768 => "0001111000011000001000",
			4769 => "0000000110011100000100",
			4770 => "0000000100101011001101",
			4771 => "0000000100101011001101",
			4772 => "0000000100101011001101",
			4773 => "0000000100101011001101",
			4774 => "0000000100101011001101",
			4775 => "0001110001101000000100",
			4776 => "0000000100101011001101",
			4777 => "0000010000111100000100",
			4778 => "0000000100101011001101",
			4779 => "0000000100101011001101",
			4780 => "0011010110010000001100",
			4781 => "0000000101000100000100",
			4782 => "0000000100101011001101",
			4783 => "0010111010010100000100",
			4784 => "0000000100101011001101",
			4785 => "0000000100101011001101",
			4786 => "0000000100101011001101",
			4787 => "0011000011011100001000",
			4788 => "0001101101011100000100",
			4789 => "0000000100101101001001",
			4790 => "0000000100101101001001",
			4791 => "0000111000100000101000",
			4792 => "0010001000100100100000",
			4793 => "0010110010001000011000",
			4794 => "0011111100100100001100",
			4795 => "0011000110000100001000",
			4796 => "0001101001011000000100",
			4797 => "0000000100101101001001",
			4798 => "0000000100101101001001",
			4799 => "0000000100101101001001",
			4800 => "0010011111000000001000",
			4801 => "0001111000011000000100",
			4802 => "0000000100101101001001",
			4803 => "0000000100101101001001",
			4804 => "0000000100101101001001",
			4805 => "0000010000111100000100",
			4806 => "0000000100101101001001",
			4807 => "0000000100101101001001",
			4808 => "0011111111100100000100",
			4809 => "0000000100101101001001",
			4810 => "0000000100101101001001",
			4811 => "0001101000010000001100",
			4812 => "0011001000000000000100",
			4813 => "0000000100101101001001",
			4814 => "0000011101111100000100",
			4815 => "0000000100101101001001",
			4816 => "0000000100101101001001",
			4817 => "0000000100101101001001",
			4818 => "0011011010011100001000",
			4819 => "0001101101011100000100",
			4820 => "0000000100101110110101",
			4821 => "1111111100101110110101",
			4822 => "0000010101011100101100",
			4823 => "0000110111010100100000",
			4824 => "0010110010001000011000",
			4825 => "0001100100110100010000",
			4826 => "0000111100010000001000",
			4827 => "0001101101111100000100",
			4828 => "0000000100101110110101",
			4829 => "0000000100101110110101",
			4830 => "0001100100110100000100",
			4831 => "0000001100101110110101",
			4832 => "0000000100101110110101",
			4833 => "0000110110111100000100",
			4834 => "0000000100101110110101",
			4835 => "0000000100101110110101",
			4836 => "0000101110110100000100",
			4837 => "0000000100101110110101",
			4838 => "1111111100101110110101",
			4839 => "0001110111010000001000",
			4840 => "0010110010001000000100",
			4841 => "0000000100101110110101",
			4842 => "0000001100101110110101",
			4843 => "0000000100101110110101",
			4844 => "0000000100101110110101",
			4845 => "0011001100110000001100",
			4846 => "0000001010110000001000",
			4847 => "0011100100001000000100",
			4848 => "0000000100110001000001",
			4849 => "0000000100110001000001",
			4850 => "0000000100110001000001",
			4851 => "0001111000000000001100",
			4852 => "0011001100110000000100",
			4853 => "0000000100110001000001",
			4854 => "0011000100011000000100",
			4855 => "0000000100110001000001",
			4856 => "0000000100110001000001",
			4857 => "0001100100110100010000",
			4858 => "0011001000000000001100",
			4859 => "0010010100111100001000",
			4860 => "0011011110101000000100",
			4861 => "0000000100110001000001",
			4862 => "0000000100110001000001",
			4863 => "0000000100110001000001",
			4864 => "0000000100110001000001",
			4865 => "0011101111010100010000",
			4866 => "0011001011000000000100",
			4867 => "0000000100110001000001",
			4868 => "0000101110110100000100",
			4869 => "0000000100110001000001",
			4870 => "0001010010011100000100",
			4871 => "0000000100110001000001",
			4872 => "0000000100110001000001",
			4873 => "0011001000000000000100",
			4874 => "0000000100110001000001",
			4875 => "0010001001101000001000",
			4876 => "0010001000010100000100",
			4877 => "0000000100110001000001",
			4878 => "0000000100110001000001",
			4879 => "0000000100110001000001",
			4880 => "0010101010100100101100",
			4881 => "0001110110000100001100",
			4882 => "0001101101011100001000",
			4883 => "0001111101100000000100",
			4884 => "0000000100110011011101",
			4885 => "0000000100110011011101",
			4886 => "1111111100110011011101",
			4887 => "0010010100111100011100",
			4888 => "0011001001110100010100",
			4889 => "0000010110101000000100",
			4890 => "0000100100110011011101",
			4891 => "0010100100111100001000",
			4892 => "0000010111100100000100",
			4893 => "0000000100110011011101",
			4894 => "1111111100110011011101",
			4895 => "0000110111010100000100",
			4896 => "0000001100110011011101",
			4897 => "0000001100110011011101",
			4898 => "0010001000100100000100",
			4899 => "0000001100110011011101",
			4900 => "1111111100110011011101",
			4901 => "1111111100110011011101",
			4902 => "0000011111001100000100",
			4903 => "1111111100110011011101",
			4904 => "0010011101011000010000",
			4905 => "0000101101101100001000",
			4906 => "0011100010011100000100",
			4907 => "0000000100110011011101",
			4908 => "0000001100110011011101",
			4909 => "0001110010110100000100",
			4910 => "0000101100110011011101",
			4911 => "0000000100110011011101",
			4912 => "0010111001010000001100",
			4913 => "0000010101011100001000",
			4914 => "0010001100011100000100",
			4915 => "0000001100110011011101",
			4916 => "1111111100110011011101",
			4917 => "1111111100110011011101",
			4918 => "0000010100110011011101",
			4919 => "0011011010011100001000",
			4920 => "0010101100011000000100",
			4921 => "0000000100110101010001",
			4922 => "1111111100110101010001",
			4923 => "0010010101010000110000",
			4924 => "0000110111010100100000",
			4925 => "0010110010001000011000",
			4926 => "0000000001010100001100",
			4927 => "0000110111011000001000",
			4928 => "0001110001101000000100",
			4929 => "0000000100110101010001",
			4930 => "0000000100110101010001",
			4931 => "0000001100110101010001",
			4932 => "0000111111010100001000",
			4933 => "0011010100101000000100",
			4934 => "0000000100110101010001",
			4935 => "0000000100110101010001",
			4936 => "0000000100110101010001",
			4937 => "0000101110110100000100",
			4938 => "0000000100110101010001",
			4939 => "1111111100110101010001",
			4940 => "0001111111011100001000",
			4941 => "0010011000010000000100",
			4942 => "0000001100110101010001",
			4943 => "0000000100110101010001",
			4944 => "0011001001110100000100",
			4945 => "0000000100110101010001",
			4946 => "0000000100110101010001",
			4947 => "0000000100110101010001",
			4948 => "0010101010100100101100",
			4949 => "0001110110000100001100",
			4950 => "0001101101011100001000",
			4951 => "0001101111001100000100",
			4952 => "0000000100110111101101",
			4953 => "0000000100110111101101",
			4954 => "1111111100110111101101",
			4955 => "0010010100111100011100",
			4956 => "0001111111011100010100",
			4957 => "0011111111010100010000",
			4958 => "0000000001010100001000",
			4959 => "0011000011011100000100",
			4960 => "0000000100110111101101",
			4961 => "0000001100110111101101",
			4962 => "0001111000011000000100",
			4963 => "0000000100110111101101",
			4964 => "0000001100110111101101",
			4965 => "0000010100110111101101",
			4966 => "0000100010000100000100",
			4967 => "0000000100110111101101",
			4968 => "1111111100110111101101",
			4969 => "1111111100110111101101",
			4970 => "0000011111001100000100",
			4971 => "1111111100110111101101",
			4972 => "0000011101011100001100",
			4973 => "0001011101000100000100",
			4974 => "0000000100110111101101",
			4975 => "0011000100010000000100",
			4976 => "0000010100110111101101",
			4977 => "0000000100110111101101",
			4978 => "0010111001010000010000",
			4979 => "0000010101011100001100",
			4980 => "0011111011101100000100",
			4981 => "1111111100110111101101",
			4982 => "0001001000001000000100",
			4983 => "0000001100110111101101",
			4984 => "0000000100110111101101",
			4985 => "1111111100110111101101",
			4986 => "0000001100110111101101",
			4987 => "0001111101100000000100",
			4988 => "1111111100111001110001",
			4989 => "0000000110011100011000",
			4990 => "0000011101011100010000",
			4991 => "0011000100011000001000",
			4992 => "0011100100001000000100",
			4993 => "0000000100111001110001",
			4994 => "0000001100111001110001",
			4995 => "0000100010011100000100",
			4996 => "0000000100111001110001",
			4997 => "0000000100111001110001",
			4998 => "0000110010000000000100",
			4999 => "0000000100111001110001",
			5000 => "0000001100111001110001",
			5001 => "0001011110101000001100",
			5002 => "0010000111110100000100",
			5003 => "0000000100111001110001",
			5004 => "0010111011011100000100",
			5005 => "1111111100111001110001",
			5006 => "0000000100111001110001",
			5007 => "0000011111001100000100",
			5008 => "1111111100111001110001",
			5009 => "0000010000111100001100",
			5010 => "0000101010000100001000",
			5011 => "0001111000011000000100",
			5012 => "0000000100111001110001",
			5013 => "1111111100111001110001",
			5014 => "0000001100111001110001",
			5015 => "0011001011011100000100",
			5016 => "1111111100111001110001",
			5017 => "0001101001111100000100",
			5018 => "0000000100111001110001",
			5019 => "0000000100111001110001",
			5020 => "0010101010100101001100",
			5021 => "0011101110101000100000",
			5022 => "0000010111100100010000",
			5023 => "0011101010111000001000",
			5024 => "0001101111001100000100",
			5025 => "0000001100111100110101",
			5026 => "1111111100111100110101",
			5027 => "0011000011011100000100",
			5028 => "0000001100111100110101",
			5029 => "0000011100111100110101",
			5030 => "0011000110000100001100",
			5031 => "0010110001111100000100",
			5032 => "1111111100111100110101",
			5033 => "0001000111010000000100",
			5034 => "0000000100111100110101",
			5035 => "0000001100111100110101",
			5036 => "1111111100111100110101",
			5037 => "0000010000111100100100",
			5038 => "0001111000011000010100",
			5039 => "0001001010000100010000",
			5040 => "0001101101111100001000",
			5041 => "0010100000001000000100",
			5042 => "0000001100111100110101",
			5043 => "0000001100111100110101",
			5044 => "0000111100010000000100",
			5045 => "1111110100111100110101",
			5046 => "0000000100111100110101",
			5047 => "0000010100111100110101",
			5048 => "0010110100010000001000",
			5049 => "0000000001010100000100",
			5050 => "0000001100111100110101",
			5051 => "1111111100111100110101",
			5052 => "0011101100010000000100",
			5053 => "1111110100111100110101",
			5054 => "1111111100111100110101",
			5055 => "0011010011001000000100",
			5056 => "1111111100111100110101",
			5057 => "0000001100111100110101",
			5058 => "0010100111110100001100",
			5059 => "0000100110101100000100",
			5060 => "1111111100111100110101",
			5061 => "0000011110010100000100",
			5062 => "0000010100111100110101",
			5063 => "0000000100111100110101",
			5064 => "0001011111100100000100",
			5065 => "1111111100111100110101",
			5066 => "0000101101000000000100",
			5067 => "0000001100111100110101",
			5068 => "1111111100111100110101",
			5069 => "0010100111110100111100",
			5070 => "0000010000111100110100",
			5071 => "0000110111010100101000",
			5072 => "0000000001010100011100",
			5073 => "0001010111100000010000",
			5074 => "0001110001101000001000",
			5075 => "0000110000110100000100",
			5076 => "0000000100111111000001",
			5077 => "0000000100111111000001",
			5078 => "0001101101111100000100",
			5079 => "0000000100111111000001",
			5080 => "1111111100111111000001",
			5081 => "0010001000100100001000",
			5082 => "0000111100000000000100",
			5083 => "0000000100111111000001",
			5084 => "0000001100111111000001",
			5085 => "0000000100111111000001",
			5086 => "0001010111100000001000",
			5087 => "0011011110101100000100",
			5088 => "0000000100111111000001",
			5089 => "0000000100111111000001",
			5090 => "0000000100111111000001",
			5091 => "0000101100000000000100",
			5092 => "0000000100111111000001",
			5093 => "0001111111011100000100",
			5094 => "0000001100111111000001",
			5095 => "0000000100111111000001",
			5096 => "0010010100111100000100",
			5097 => "0000000100111111000001",
			5098 => "0000000100111111000001",
			5099 => "0011010011000000000100",
			5100 => "1111111100111111000001",
			5101 => "0001110000110100000100",
			5102 => "0000000100111111000001",
			5103 => "0000000100111111000001",
			5104 => "0001111101100000000100",
			5105 => "1111111101000001000101",
			5106 => "0010100111101100010000",
			5107 => "0000011101011100001100",
			5108 => "0011100100001000000100",
			5109 => "0000000101000001000101",
			5110 => "0001001001100000000100",
			5111 => "0000000101000001000101",
			5112 => "0000000101000001000101",
			5113 => "0000000101000001000101",
			5114 => "0001010101001000011000",
			5115 => "0001110001101000010000",
			5116 => "0001111000000000000100",
			5117 => "0000000101000001000101",
			5118 => "0010001100011100001000",
			5119 => "0010000111110100000100",
			5120 => "0000000101000001000101",
			5121 => "0000000101000001000101",
			5122 => "0000000101000001000101",
			5123 => "0001111111011100000100",
			5124 => "0000000101000001000101",
			5125 => "0000000101000001000101",
			5126 => "0000010000111100010000",
			5127 => "0010110010001000000100",
			5128 => "0000000101000001000101",
			5129 => "0001111111011100001000",
			5130 => "0000111010000100000100",
			5131 => "0000000101000001000101",
			5132 => "0000000101000001000101",
			5133 => "0000000101000001000101",
			5134 => "0000111111100000000100",
			5135 => "0000000101000001000101",
			5136 => "0000000101000001000101",
			5137 => "0000001011010100111100",
			5138 => "0011000001101000111000",
			5139 => "0010100111101100011000",
			5140 => "0000101100100100010100",
			5141 => "0000010111100100001100",
			5142 => "0011111011000000000100",
			5143 => "0000000101000011100001",
			5144 => "0000011001111000000100",
			5145 => "0000000101000011100001",
			5146 => "0000001101000011100001",
			5147 => "0011001100110000000100",
			5148 => "0000000101000011100001",
			5149 => "1111111101000011100001",
			5150 => "0000001101000011100001",
			5151 => "0000111100010000010000",
			5152 => "0001101101111100001000",
			5153 => "0000011111001100000100",
			5154 => "0000000101000011100001",
			5155 => "0000000101000011100001",
			5156 => "0011000100011000000100",
			5157 => "0000000101000011100001",
			5158 => "1111111101000011100001",
			5159 => "0010100000001000000100",
			5160 => "0000001101000011100001",
			5161 => "0001101101111100000100",
			5162 => "1111111101000011100001",
			5163 => "0001111000011000000100",
			5164 => "0000000101000011100001",
			5165 => "0000000101000011100001",
			5166 => "0000100101000011100001",
			5167 => "0010110101100100000100",
			5168 => "1111111101000011100001",
			5169 => "0010111011011100001000",
			5170 => "0010010100101100000100",
			5171 => "0000001101000011100001",
			5172 => "0000000101000011100001",
			5173 => "0001011111100100000100",
			5174 => "1111111101000011100001",
			5175 => "0000000101000011100001",
			5176 => "0010001000100100110100",
			5177 => "0011101000011000010100",
			5178 => "0001101101011100001000",
			5179 => "0010100100110100000100",
			5180 => "1111111101000110110101",
			5181 => "0000100101000110110101",
			5182 => "0011101011000000000100",
			5183 => "1111111101000110110101",
			5184 => "0000010111100100000100",
			5185 => "0000011101000110110101",
			5186 => "1111111101000110110101",
			5187 => "0000010000111100011000",
			5188 => "0001111101111000000100",
			5189 => "0000101101000110110101",
			5190 => "0011100111110000000100",
			5191 => "1111111101000110110101",
			5192 => "0011010111111100001000",
			5193 => "0001111111011100000100",
			5194 => "0000010101000110110101",
			5195 => "0000001101000110110101",
			5196 => "0011001000000000000100",
			5197 => "0000010101000110110101",
			5198 => "0000001101000110110101",
			5199 => "0001101101111100000100",
			5200 => "0000001101000110110101",
			5201 => "1111111101000110110101",
			5202 => "0000001001101000011000",
			5203 => "0000010000111100010100",
			5204 => "0000110000010000010000",
			5205 => "0011001011000000000100",
			5206 => "0000010101000110110101",
			5207 => "0010101010100000000100",
			5208 => "1111111101000110110101",
			5209 => "0001111000011000000100",
			5210 => "0000010101000110110101",
			5211 => "1111111101000110110101",
			5212 => "0000101101000110110101",
			5213 => "1111111101000110110101",
			5214 => "0010100010101100001100",
			5215 => "0001001101101100000100",
			5216 => "1111111101000110110101",
			5217 => "0000011100110100000100",
			5218 => "1111111101000110110101",
			5219 => "0000011101000110110101",
			5220 => "0011010011000000000100",
			5221 => "1111111101000110110101",
			5222 => "0011010010010100001100",
			5223 => "0001011000100000001000",
			5224 => "0001011111100100000100",
			5225 => "0000000101000110110101",
			5226 => "0000001101000110110101",
			5227 => "1111111101000110110101",
			5228 => "1111111101000110110101",
			5229 => "0010001001000101001100",
			5230 => "0001100100110100101000",
			5231 => "0011101110101000010100",
			5232 => "0001100001000100010000",
			5233 => "0011000110000100001100",
			5234 => "0011100100001000000100",
			5235 => "0000000101001001111001",
			5236 => "0010010101011100000100",
			5237 => "0000001101001001111001",
			5238 => "0000000101001001111001",
			5239 => "0000000101001001111001",
			5240 => "1111111101001001111001",
			5241 => "0010010100111100010000",
			5242 => "0001111111011100001100",
			5243 => "0001111000011000001000",
			5244 => "0001110001101000000100",
			5245 => "0000001101001001111001",
			5246 => "0000000101001001111001",
			5247 => "0000001101001001111001",
			5248 => "0000000101001001111001",
			5249 => "0000000101001001111001",
			5250 => "0000111000001100011100",
			5251 => "0001000111011000010100",
			5252 => "0010110110110100001100",
			5253 => "0011101001100000001000",
			5254 => "0010001000100100000100",
			5255 => "0000000101001001111001",
			5256 => "0000000101001001111001",
			5257 => "0000000101001001111001",
			5258 => "0010011111000000000100",
			5259 => "0000001101001001111001",
			5260 => "0000000101001001111001",
			5261 => "0011000100011000000100",
			5262 => "0000000101001001111001",
			5263 => "1111111101001001111001",
			5264 => "0010110101110100000100",
			5265 => "0000001101001001111001",
			5266 => "0000000101001001111001",
			5267 => "0010110101110100000100",
			5268 => "1111111101001001111001",
			5269 => "0011001001110100001000",
			5270 => "0000010101011100000100",
			5271 => "0000001101001001111001",
			5272 => "0000000101001001111001",
			5273 => "0011010011000000000100",
			5274 => "1111111101001001111001",
			5275 => "0011011111101000000100",
			5276 => "0000000101001001111001",
			5277 => "0000000101001001111001",
			5278 => "0000000010111101001100",
			5279 => "0000111010000100110000",
			5280 => "0000000101000100011100",
			5281 => "0000101101000100010100",
			5282 => "0010010000111100001100",
			5283 => "0011100100001000000100",
			5284 => "0000000101001100010101",
			5285 => "0001111101100000000100",
			5286 => "0000000101001100010101",
			5287 => "0000000101001100010101",
			5288 => "0010011110010100000100",
			5289 => "0000000101001100010101",
			5290 => "0000000101001100010101",
			5291 => "0001101101111100000100",
			5292 => "0000000101001100010101",
			5293 => "0000000101001100010101",
			5294 => "0010001000100100000100",
			5295 => "0000000101001100010101",
			5296 => "0010100000001000000100",
			5297 => "0000000101001100010101",
			5298 => "0011111111010100001000",
			5299 => "0011001001110100000100",
			5300 => "0000000101001100010101",
			5301 => "0000000101001100010101",
			5302 => "0000000101001100010101",
			5303 => "0001111111011100001100",
			5304 => "0010011000010000001000",
			5305 => "0001100100110100000100",
			5306 => "0000000101001100010101",
			5307 => "0000000101001100010101",
			5308 => "0000000101001100010101",
			5309 => "0001011110010000000100",
			5310 => "0000000101001100010101",
			5311 => "0010011010100000001000",
			5312 => "0001101000010000000100",
			5313 => "0000000101001100010101",
			5314 => "0000000101001100010101",
			5315 => "0000000101001100010101",
			5316 => "1111111101001100010101",
			5317 => "0010100010101101001100",
			5318 => "0000010000111101000000",
			5319 => "0011101110101000100000",
			5320 => "0000000110011000011100",
			5321 => "0011001100110000010000",
			5322 => "0011111011000000001000",
			5323 => "0001101111001100000100",
			5324 => "0000001101001111011001",
			5325 => "1111111101001111011001",
			5326 => "0010010101011100000100",
			5327 => "0000010101001111011001",
			5328 => "0000001101001111011001",
			5329 => "0001111110001100001000",
			5330 => "0010011011111100000100",
			5331 => "0000000101001111011001",
			5332 => "0000001101001111011001",
			5333 => "1111111101001111011001",
			5334 => "1111111101001111011001",
			5335 => "0000111000001100011000",
			5336 => "0000000001010100001100",
			5337 => "0010010100111100001000",
			5338 => "0011100010000100000100",
			5339 => "0000001101001111011001",
			5340 => "0000001101001111011001",
			5341 => "1111111101001111011001",
			5342 => "0011001011000000000100",
			5343 => "0000001101001111011001",
			5344 => "0000110111010100000100",
			5345 => "1111111101001111011001",
			5346 => "0000000101001111011001",
			5347 => "0001111000011000000100",
			5348 => "0000010101001111011001",
			5349 => "0000001101001111011001",
			5350 => "0010010100111100001000",
			5351 => "0001011001010000000100",
			5352 => "1111111101001111011001",
			5353 => "0000001101001111011001",
			5354 => "1111111101001111011001",
			5355 => "0010100011101000001100",
			5356 => "0001001111101000000100",
			5357 => "1111111101001111011001",
			5358 => "0000001000101100000100",
			5359 => "0000011101001111011001",
			5360 => "0000000101001111011001",
			5361 => "0001011111100100000100",
			5362 => "1111111101001111011001",
			5363 => "0001011000100000000100",
			5364 => "0000000101001111011001",
			5365 => "1111111101001111011001",
			5366 => "0010101010100101010000",
			5367 => "0011101110101000101100",
			5368 => "0001101001011000011000",
			5369 => "0011000110000100010100",
			5370 => "0011100100001000000100",
			5371 => "1111111101010010100101",
			5372 => "0000010110101000001000",
			5373 => "0011001000111000000100",
			5374 => "0000010101010010100101",
			5375 => "0000000101010010100101",
			5376 => "0010010101011100000100",
			5377 => "0000000101010010100101",
			5378 => "0000000101010010100101",
			5379 => "0000101101010010100101",
			5380 => "0010110100001000000100",
			5381 => "1111111101010010100101",
			5382 => "0011000110000100001100",
			5383 => "0001000111010000000100",
			5384 => "0000000101010010100101",
			5385 => "0000010111100100000100",
			5386 => "0000001101010010100101",
			5387 => "0000000101010010100101",
			5388 => "1111111101010010100101",
			5389 => "0010010100111100100000",
			5390 => "0001111111011100010100",
			5391 => "0000110111010100010000",
			5392 => "0001101101111100001000",
			5393 => "0011010111111100000100",
			5394 => "0000001101010010100101",
			5395 => "0000000101010010100101",
			5396 => "0000111100010000000100",
			5397 => "1111110101010010100101",
			5398 => "0000000101010010100101",
			5399 => "0000010101010010100101",
			5400 => "0001111111011100001000",
			5401 => "0011101100010000000100",
			5402 => "0000001101010010100101",
			5403 => "1111111101010010100101",
			5404 => "1111111101010010100101",
			5405 => "1111111101010010100101",
			5406 => "0010100111110100001100",
			5407 => "0000100110101100000100",
			5408 => "1111111101010010100101",
			5409 => "0000111000100000000100",
			5410 => "0000011101010010100101",
			5411 => "0000001101010010100101",
			5412 => "0001011111100100000100",
			5413 => "1111111101010010100101",
			5414 => "0000101101000000000100",
			5415 => "0000001101010010100101",
			5416 => "1111111101010010100101",
			5417 => "0001111101100000000100",
			5418 => "1111111101010100110001",
			5419 => "0010100111101100001100",
			5420 => "0011100100001000000100",
			5421 => "0000000101010100110001",
			5422 => "0011000100011000000100",
			5423 => "0000000101010100110001",
			5424 => "0000000101010100110001",
			5425 => "0001010101001000011000",
			5426 => "0011011010001000010100",
			5427 => "0011010111111100010000",
			5428 => "0000111100010000001000",
			5429 => "0010000111110100000100",
			5430 => "0000000101010100110001",
			5431 => "0000000101010100110001",
			5432 => "0000011001011000000100",
			5433 => "0000000101010100110001",
			5434 => "0000000101010100110001",
			5435 => "1111111101010100110001",
			5436 => "0000000101010100110001",
			5437 => "0010110100010000001100",
			5438 => "0011010111111100000100",
			5439 => "0000000101010100110001",
			5440 => "0011011010001000000100",
			5441 => "0000000101010100110001",
			5442 => "0000000101010100110001",
			5443 => "0001110111010000001100",
			5444 => "0000010000111100001000",
			5445 => "0011010111111100000100",
			5446 => "0000000101010100110001",
			5447 => "0000000101010100110001",
			5448 => "0000000101010100110001",
			5449 => "0011011111101000000100",
			5450 => "0000000101010100110001",
			5451 => "0000000101010100110001",
			5452 => "0011011010011100001000",
			5453 => "0010101100011000000100",
			5454 => "0000000101010110110101",
			5455 => "1111111101010110110101",
			5456 => "0000010101011100111000",
			5457 => "0000110111010100101000",
			5458 => "0010110010001000100000",
			5459 => "0000111100010000010000",
			5460 => "0010100111101100001000",
			5461 => "0011111010011100000100",
			5462 => "0000000101010110110101",
			5463 => "0000000101010110110101",
			5464 => "0010000111110100000100",
			5465 => "0000000101010110110101",
			5466 => "1111111101010110110101",
			5467 => "0000011001011000001000",
			5468 => "0001111111011100000100",
			5469 => "0000001101010110110101",
			5470 => "0000000101010110110101",
			5471 => "0000000001010100000100",
			5472 => "0000000101010110110101",
			5473 => "0000000101010110110101",
			5474 => "0000101110110100000100",
			5475 => "0000000101010110110101",
			5476 => "1111111101010110110101",
			5477 => "0001110111010000001100",
			5478 => "0010110010001000000100",
			5479 => "0000000101010110110101",
			5480 => "0001111111011100000100",
			5481 => "0000001101010110110101",
			5482 => "0000000101010110110101",
			5483 => "0000000101010110110101",
			5484 => "0000000101010110110101",
			5485 => "0000001100000101010100",
			5486 => "0011001000000000110100",
			5487 => "0011101110101000010100",
			5488 => "0001100001000100010000",
			5489 => "0011000110000100001100",
			5490 => "0011100100001000000100",
			5491 => "0000000101011010001001",
			5492 => "0010010000111100000100",
			5493 => "0000001101011010001001",
			5494 => "0000000101011010001001",
			5495 => "0000000101011010001001",
			5496 => "1111111101011010001001",
			5497 => "0010100000001000001000",
			5498 => "0000010000111100000100",
			5499 => "0000001101011010001001",
			5500 => "0000000101011010001001",
			5501 => "0000111010000100001100",
			5502 => "0010110000011100000100",
			5503 => "0000000101011010001001",
			5504 => "0000001100000100000100",
			5505 => "1111111101011010001001",
			5506 => "0000000101011010001001",
			5507 => "0000000001110000000100",
			5508 => "0000001101011010001001",
			5509 => "0001010101001000000100",
			5510 => "0000000101011010001001",
			5511 => "0000000101011010001001",
			5512 => "0000111001100000000100",
			5513 => "1111111101011010001001",
			5514 => "0001000111011000001000",
			5515 => "0010100000001000000100",
			5516 => "0000001101011010001001",
			5517 => "0000000101011010001001",
			5518 => "0011001000000000001000",
			5519 => "0000000001010100000100",
			5520 => "0000001101011010001001",
			5521 => "0000000101011010001001",
			5522 => "0010001000010100000100",
			5523 => "1111111101011010001001",
			5524 => "0010110100010000000100",
			5525 => "0000001101011010001001",
			5526 => "0000000101011010001001",
			5527 => "0011011111010000000100",
			5528 => "1111111101011010001001",
			5529 => "0001101011001100001000",
			5530 => "0010011000010000000100",
			5531 => "0000001101011010001001",
			5532 => "0000000101011010001001",
			5533 => "0011010011000000000100",
			5534 => "1111111101011010001001",
			5535 => "0011001011011100000100",
			5536 => "0000001101011010001001",
			5537 => "0000000101011010001001",
			5538 => "0000001100000101100000",
			5539 => "0010001000100100100000",
			5540 => "0011100100001000000100",
			5541 => "0000000101011101110101",
			5542 => "0000010110101000001100",
			5543 => "0010111101111000001000",
			5544 => "0011001000111000000100",
			5545 => "0000001101011101110101",
			5546 => "0000000101011101110101",
			5547 => "0000011101011101110101",
			5548 => "0010110100001000000100",
			5549 => "1111111101011101110101",
			5550 => "0000010000111100001000",
			5551 => "0001101101111100000100",
			5552 => "0000001101011101110101",
			5553 => "0000000101011101110101",
			5554 => "0000000101011101110101",
			5555 => "0001111000011000100000",
			5556 => "0001110001101000010000",
			5557 => "0011010101110000001000",
			5558 => "0000101001100000000100",
			5559 => "1111111101011101110101",
			5560 => "0000000101011101110101",
			5561 => "0000010000111100000100",
			5562 => "0000001101011101110101",
			5563 => "0000000101011101110101",
			5564 => "0000100010000100001000",
			5565 => "0001010111100000000100",
			5566 => "0000000101011101110101",
			5567 => "1111111101011101110101",
			5568 => "0001011001010000000100",
			5569 => "1111110101011101110101",
			5570 => "0000000101011101110101",
			5571 => "0001111000011000010000",
			5572 => "0011101100010000001000",
			5573 => "0010011111000000000100",
			5574 => "0000001101011101110101",
			5575 => "0000000101011101110101",
			5576 => "0011011001011100000100",
			5577 => "0000100101011101110101",
			5578 => "0000001101011101110101",
			5579 => "0001100100110100000100",
			5580 => "0000001101011101110101",
			5581 => "0001000000010000001000",
			5582 => "0001010101001000000100",
			5583 => "0000000101011101110101",
			5584 => "1111111101011101110101",
			5585 => "0000000101011101110101",
			5586 => "0000011111001100000100",
			5587 => "1111111101011101110101",
			5588 => "0010011101011000001000",
			5589 => "0001101011001100000100",
			5590 => "0000010101011101110101",
			5591 => "0000000101011101110101",
			5592 => "0001010000010000001000",
			5593 => "0001101010011000000100",
			5594 => "0000000101011101110101",
			5595 => "1111111101011101110101",
			5596 => "0000001101011101110101",
			5597 => "0000001011010101001100",
			5598 => "0011000001101001001000",
			5599 => "0010000111110100011100",
			5600 => "0011101110101000010100",
			5601 => "0000010111100100001100",
			5602 => "0011101011000000001000",
			5603 => "0011000110000100000100",
			5604 => "0000000101100000110001",
			5605 => "0000000101100000110001",
			5606 => "0000001101100000110001",
			5607 => "0011001100110000000100",
			5608 => "0000000101100000110001",
			5609 => "1111111101100000110001",
			5610 => "0010011001100100000100",
			5611 => "0000001101100000110001",
			5612 => "0000000101100000110001",
			5613 => "0000111100010000010100",
			5614 => "0011000100011000001100",
			5615 => "0011011110000100001000",
			5616 => "0001110110100100000100",
			5617 => "0000000101100000110001",
			5618 => "0000000101100000110001",
			5619 => "0000000101100000110001",
			5620 => "0010110101100100000100",
			5621 => "0000000101100000110001",
			5622 => "1111111101100000110001",
			5623 => "0010001000100100001000",
			5624 => "0010110101100100000100",
			5625 => "0000000101100000110001",
			5626 => "0000001101100000110001",
			5627 => "0000111010000100001000",
			5628 => "0010110010001000000100",
			5629 => "0000000101100000110001",
			5630 => "1111111101100000110001",
			5631 => "0000000001010100000100",
			5632 => "0000001101100000110001",
			5633 => "0000000101100000110001",
			5634 => "0000010101100000110001",
			5635 => "0010110101100100000100",
			5636 => "1111111101100000110001",
			5637 => "0010111011011100001000",
			5638 => "0011100110111100000100",
			5639 => "0000001101100000110001",
			5640 => "0000000101100000110001",
			5641 => "0001011111100100000100",
			5642 => "1111111101100000110001",
			5643 => "0000000101100000110001",
			5644 => "0000001001101001011000",
			5645 => "0011101110101000100000",
			5646 => "0000100000110100011100",
			5647 => "0001111100101000011000",
			5648 => "0011100001101000010000",
			5649 => "0011000110000100001000",
			5650 => "0011000100000000000100",
			5651 => "0000000101100100100101",
			5652 => "1111111101100100100101",
			5653 => "0001010110100100000100",
			5654 => "0000001101100100100101",
			5655 => "0000000101100100100101",
			5656 => "0011000110000100000100",
			5657 => "0000001101100100100101",
			5658 => "0000000101100100100101",
			5659 => "1111111101100100100101",
			5660 => "1111111101100100100101",
			5661 => "0011001000000000011000",
			5662 => "0010010100111100010100",
			5663 => "0001111111011100010000",
			5664 => "0001111000011000001000",
			5665 => "0010011111000000000100",
			5666 => "0000001101100100100101",
			5667 => "0000000101100100100101",
			5668 => "0000100110010000000100",
			5669 => "0000000101100100100101",
			5670 => "0000001101100100100101",
			5671 => "0000000101100100100101",
			5672 => "1111111101100100100101",
			5673 => "0011011010001000010100",
			5674 => "0000000101000100001000",
			5675 => "0000111100000000000100",
			5676 => "0000000101100100100101",
			5677 => "0000001101100100100101",
			5678 => "0000101111010100001000",
			5679 => "0010111011011100000100",
			5680 => "0000000101100100100101",
			5681 => "1111111101100100100101",
			5682 => "0000000101100100100101",
			5683 => "0010110100010000000100",
			5684 => "0000001101100100100101",
			5685 => "0011100111010100000100",
			5686 => "0000000101100100100101",
			5687 => "0000000101100100100101",
			5688 => "0000100010110000010100",
			5689 => "0010000110011100010000",
			5690 => "0011011111010000000100",
			5691 => "1111111101100100100101",
			5692 => "0010111011011100001000",
			5693 => "0011100110111100000100",
			5694 => "0000001101100100100101",
			5695 => "0000000101100100100101",
			5696 => "1111111101100100100101",
			5697 => "1111111101100100100101",
			5698 => "0010100001010000001100",
			5699 => "0001010010000000000100",
			5700 => "0000011101100100100101",
			5701 => "0000111101001000000100",
			5702 => "0000000101100100100101",
			5703 => "0000001101100100100101",
			5704 => "1111111101100100100101",
			5705 => "0010001001000101100000",
			5706 => "0010001000100100100000",
			5707 => "0011100100001000000100",
			5708 => "0000000101101000011001",
			5709 => "0000010110101000000100",
			5710 => "0000001101101000011001",
			5711 => "0011110010001000001100",
			5712 => "0000010111100100001000",
			5713 => "0001110110000100000100",
			5714 => "0000000101101000011001",
			5715 => "0000001101101000011001",
			5716 => "1111111101101000011001",
			5717 => "0010011111000000000100",
			5718 => "0000001101101000011001",
			5719 => "0001101101111100000100",
			5720 => "0000001101101000011001",
			5721 => "0000000101101000011001",
			5722 => "0001111000011000100000",
			5723 => "0001110001101000010000",
			5724 => "0011010101110000001000",
			5725 => "0000101001100000000100",
			5726 => "1111111101101000011001",
			5727 => "0000000101101000011001",
			5728 => "0010010100111100000100",
			5729 => "0000001101101000011001",
			5730 => "0000000101101000011001",
			5731 => "0000100010000100001000",
			5732 => "0001010111100000000100",
			5733 => "0000000101101000011001",
			5734 => "1111111101101000011001",
			5735 => "0011110110111100000100",
			5736 => "1111110101101000011001",
			5737 => "0000000101101000011001",
			5738 => "0001111000011000010000",
			5739 => "0000111010000100001000",
			5740 => "0010011111000000000100",
			5741 => "0000001101101000011001",
			5742 => "0000000101101000011001",
			5743 => "0000010000111100000100",
			5744 => "0000001101101000011001",
			5745 => "0000000101101000011001",
			5746 => "0001100100110100000100",
			5747 => "0000001101101000011001",
			5748 => "0011010011001000001000",
			5749 => "0001010101001000000100",
			5750 => "0000000101101000011001",
			5751 => "1111111101101000011001",
			5752 => "0000000101101000011001",
			5753 => "0000011111001100000100",
			5754 => "1111111101101000011001",
			5755 => "0010011101011000001000",
			5756 => "0010001001101000000100",
			5757 => "0000001101101000011001",
			5758 => "0000000101101000011001",
			5759 => "0001010000010000001100",
			5760 => "0010000001010000001000",
			5761 => "0010010101010000000100",
			5762 => "0000000101101000011001",
			5763 => "0000000101101000011001",
			5764 => "1111111101101000011001",
			5765 => "0000001101101000011001",
			5766 => "0001111101100000000100",
			5767 => "1111111101101011011101",
			5768 => "0001111000011000111100",
			5769 => "0010000111110100011000",
			5770 => "0000101101000100010000",
			5771 => "0001101101011100000100",
			5772 => "0000001101101011011101",
			5773 => "0011001100110000001000",
			5774 => "0011111010011100000100",
			5775 => "0000000101101011011101",
			5776 => "0000000101101011011101",
			5777 => "0000000101101011011101",
			5778 => "0010011001100100000100",
			5779 => "0000001101101011011101",
			5780 => "0000000101101011011101",
			5781 => "0011010010011100010100",
			5782 => "0000000110011100000100",
			5783 => "0000000101101011011101",
			5784 => "0011110111011000001000",
			5785 => "0001110001101000000100",
			5786 => "1111111101101011011101",
			5787 => "0000000101101011011101",
			5788 => "0001011100100100000100",
			5789 => "0000000101101011011101",
			5790 => "0000000101101011011101",
			5791 => "0010100000001000000100",
			5792 => "0000001101101011011101",
			5793 => "0001101101111100000100",
			5794 => "1111111101101011011101",
			5795 => "0001101100011000000100",
			5796 => "0000000101101011011101",
			5797 => "0000000101101011011101",
			5798 => "0001111111011100010000",
			5799 => "0010011000010000001100",
			5800 => "0000100110010000000100",
			5801 => "0000000101101011011101",
			5802 => "0011010101110000000100",
			5803 => "0000000101101011011101",
			5804 => "0000001101101011011101",
			5805 => "0000000101101011011101",
			5806 => "0011101011111000000100",
			5807 => "0000000101101011011101",
			5808 => "0010011010100000001100",
			5809 => "0010001001101000001000",
			5810 => "0001100101010000000100",
			5811 => "0000000101101011011101",
			5812 => "0000000101101011011101",
			5813 => "0000000101101011011101",
			5814 => "0000000101101011011101",
			5815 => "0001111101100000000100",
			5816 => "1111111101101110010011",
			5817 => "0010100001010001010100",
			5818 => "0011011010001000111100",
			5819 => "0010100000001000100000",
			5820 => "0011000100011000010000",
			5821 => "0000101101000100001000",
			5822 => "0001111100101000000100",
			5823 => "0000000101101110010011",
			5824 => "0000000101101110010011",
			5825 => "0000010000111100000100",
			5826 => "0000001101101110010011",
			5827 => "0000000101101110010011",
			5828 => "0001011100100100001000",
			5829 => "0001101101111100000100",
			5830 => "0000000101101110010011",
			5831 => "1111111101101110010011",
			5832 => "0000101110110100000100",
			5833 => "0000001101101110010011",
			5834 => "0000000101101110010011",
			5835 => "0000111010000100001100",
			5836 => "0011111111010100001000",
			5837 => "0001101101111100000100",
			5838 => "0000000101101110010011",
			5839 => "1111111101101110010011",
			5840 => "0000000101101110010011",
			5841 => "0000100111011000001000",
			5842 => "0001111000011000000100",
			5843 => "0000000101101110010011",
			5844 => "0000000101101110010011",
			5845 => "0000100110101100000100",
			5846 => "1111111101101110010011",
			5847 => "0000000101101110010011",
			5848 => "0001111111011100001000",
			5849 => "0000010000111100000100",
			5850 => "0000001101101110010011",
			5851 => "0000000101101110010011",
			5852 => "0000111000101000000100",
			5853 => "0000000101101110010011",
			5854 => "0000011101111100001000",
			5855 => "0011010110010000000100",
			5856 => "0000000101101110010011",
			5857 => "0000001101101110010011",
			5858 => "0000000101101110010011",
			5859 => "1111111101101110010011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1940, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3878, initial_addr_3'length));
	end generate gen_rom_4;

	gen_rom_5: if SELECT_ROM = 5 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000000000000001110101",
			29 => "0000000000000001111001",
			30 => "0000000000000001111101",
			31 => "0000000000000010000001",
			32 => "0000000000000010000101",
			33 => "0001001011001000000100",
			34 => "0000000000000010010001",
			35 => "0000000000000010010001",
			36 => "0001001011001000000100",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0001001011001000000100",
			40 => "0000000000000010101001",
			41 => "0000000000000010101001",
			42 => "0001110111010000000100",
			43 => "0000000000000010110101",
			44 => "0000000000000010110101",
			45 => "0000101110000000000100",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0001001011100100000100",
			49 => "0000000000000011001101",
			50 => "0000000000000011001101",
			51 => "0011000100011000000100",
			52 => "0000000000000011011001",
			53 => "0000000000000011011001",
			54 => "0001001011100100000100",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0001000001100100000100",
			58 => "0000000000000011110001",
			59 => "0000000000000011110001",
			60 => "0001001011100100000100",
			61 => "0000000000000011111101",
			62 => "0000000000000011111101",
			63 => "0011000100011000000100",
			64 => "0000000000000100001001",
			65 => "0000000000000100001001",
			66 => "0011001001110100000100",
			67 => "0000000000000100011101",
			68 => "0000011101011100000100",
			69 => "0000000000000100011101",
			70 => "0000000000000100011101",
			71 => "0001111111011100000100",
			72 => "0000000000000100110001",
			73 => "0000011101011100000100",
			74 => "0000000000000100110001",
			75 => "0000000000000100110001",
			76 => "0011000100011000000100",
			77 => "0000000000000101000101",
			78 => "0011110100101000000100",
			79 => "0000000000000101000101",
			80 => "0000000000000101000101",
			81 => "0001110111010000001000",
			82 => "0001001111101100000100",
			83 => "0000000000000101100001",
			84 => "0000000000000101100001",
			85 => "0010010100111100000100",
			86 => "0000000000000101100001",
			87 => "0000000000000101100001",
			88 => "0001111111011100001000",
			89 => "0001001010101000000100",
			90 => "0000000000000101111101",
			91 => "0000000000000101111101",
			92 => "0000010000111100000100",
			93 => "0000000000000101111101",
			94 => "0000000000000101111101",
			95 => "0000100101010100000100",
			96 => "1111111000000110011001",
			97 => "0010011000010000001000",
			98 => "0001100101010000000100",
			99 => "0000010000000110011001",
			100 => "0000001000000110011001",
			101 => "1111111000000110011001",
			102 => "0011000100011000000100",
			103 => "1111111000000110110101",
			104 => "0000011111001100001000",
			105 => "0011110100101000000100",
			106 => "0000000000000110110101",
			107 => "0000000000000110110101",
			108 => "0000000000000110110101",
			109 => "0011001001110100000100",
			110 => "0000000000000111010001",
			111 => "0000011101011100001000",
			112 => "0010001101100000000100",
			113 => "0000000000000111010001",
			114 => "0000000000000111010001",
			115 => "0000000000000111010001",
			116 => "0011000100011000000100",
			117 => "0000000000000111101101",
			118 => "0000101111010100000100",
			119 => "0000000000000111101101",
			120 => "0000110100000100000100",
			121 => "0000000000000111101101",
			122 => "0000000000000111101101",
			123 => "0011000100011000000100",
			124 => "0000000000001000001001",
			125 => "0000101111010100000100",
			126 => "0000000000001000001001",
			127 => "0011110100101000000100",
			128 => "0000000000001000001001",
			129 => "0000000000001000001001",
			130 => "0011000100011000000100",
			131 => "0000000000001000100101",
			132 => "0011110100101000000100",
			133 => "0000000000001000100101",
			134 => "0000101111010100000100",
			135 => "0000000000001000100101",
			136 => "0000000000001000100101",
			137 => "0011000100011000000100",
			138 => "0000000000001001000001",
			139 => "0000101111010100000100",
			140 => "0000000000001001000001",
			141 => "0000110100000100000100",
			142 => "0000000000001001000001",
			143 => "0000000000001001000001",
			144 => "0000100101010100001100",
			145 => "0001000000000100000100",
			146 => "1111111000001001100101",
			147 => "0000110100000100000100",
			148 => "1111111000001001100101",
			149 => "0000001000001001100101",
			150 => "0000010000111100000100",
			151 => "0000001000001001100101",
			152 => "1111111000001001100101",
			153 => "0000100101010100001100",
			154 => "0001111111011100000100",
			155 => "1111111000001010001001",
			156 => "0010110010001000000100",
			157 => "0000001000001010001001",
			158 => "1111111000001010001001",
			159 => "0000010000111100000100",
			160 => "0000001000001010001001",
			161 => "0000000000001010001001",
			162 => "0001111111011100001100",
			163 => "0000101110000000000100",
			164 => "1111111000001010101101",
			165 => "0000001100001000000100",
			166 => "0000000000001010101101",
			167 => "0000000000001010101101",
			168 => "0000011111001100000100",
			169 => "0000001000001010101101",
			170 => "0000000000001010101101",
			171 => "0011001001110100001000",
			172 => "0001000100110000000100",
			173 => "1111111000001011010001",
			174 => "0000000000001011010001",
			175 => "0000011101011100001000",
			176 => "0000000101100100000100",
			177 => "0000001000001011010001",
			178 => "0000000000001011010001",
			179 => "0000000000001011010001",
			180 => "0011001001110100001000",
			181 => "0001000100110000000100",
			182 => "1111111000001011110101",
			183 => "0000000000001011110101",
			184 => "0000010000111100001000",
			185 => "0001111000011000000100",
			186 => "0000000000001011110101",
			187 => "0000000000001011110101",
			188 => "0000000000001011110101",
			189 => "0011000100011000000100",
			190 => "1111111000001100011001",
			191 => "0000011111001100001000",
			192 => "0001111111011100000100",
			193 => "0000000000001100011001",
			194 => "0000001000001100011001",
			195 => "0011001011011100000100",
			196 => "0000000000001100011001",
			197 => "0000000000001100011001",
			198 => "0011000100011000000100",
			199 => "1111111000001100111101",
			200 => "0000011111001100001000",
			201 => "0011110100101000000100",
			202 => "0000000000001100111101",
			203 => "0000000000001100111101",
			204 => "0000001101111000000100",
			205 => "0000000000001100111101",
			206 => "0000000000001100111101",
			207 => "0000100011110100010000",
			208 => "0000101110111000001000",
			209 => "0000100101010100000100",
			210 => "1101010000001101101001",
			211 => "1101011000001101101001",
			212 => "0000010111101000000100",
			213 => "1110101000001101101001",
			214 => "1101010000001101101001",
			215 => "0000011101111100000100",
			216 => "1110110000001101101001",
			217 => "1101010000001101101001",
			218 => "0001001011001000000100",
			219 => "1111111000001110001101",
			220 => "0011000100011000000100",
			221 => "0000000000001110001101",
			222 => "0000010000111100001000",
			223 => "0000010010001100000100",
			224 => "0000000000001110001101",
			225 => "0000000000001110001101",
			226 => "0000000000001110001101",
			227 => "0011000100011000000100",
			228 => "1111111000001110110001",
			229 => "0000011111001100001100",
			230 => "0001101010011000000100",
			231 => "0000000000001110110001",
			232 => "0000000101110100000100",
			233 => "0000000000001110110001",
			234 => "0000000000001110110001",
			235 => "0000000000001110110001",
			236 => "0001001011001000000100",
			237 => "0000000000001111010101",
			238 => "0011000100011000000100",
			239 => "0000000000001111010101",
			240 => "0000010000111100001000",
			241 => "0000010010001100000100",
			242 => "0000000000001111010101",
			243 => "0000000000001111010101",
			244 => "0000000000001111010101",
			245 => "0011000100011000000100",
			246 => "0000000000001111111001",
			247 => "0000010000111100001100",
			248 => "0000101111010100000100",
			249 => "0000000000001111111001",
			250 => "0000000101110100000100",
			251 => "0000000000001111111001",
			252 => "0000000000001111111001",
			253 => "0000000000001111111001",
			254 => "0011000100011000000100",
			255 => "0000000000010000011101",
			256 => "0000010000111100001100",
			257 => "0011110100101000000100",
			258 => "0000000000010000011101",
			259 => "0000101111010100000100",
			260 => "0000000000010000011101",
			261 => "0000000000010000011101",
			262 => "0000000000010000011101",
			263 => "0000100101010100010000",
			264 => "0011000100011000000100",
			265 => "1111111000010001001001",
			266 => "0001000000000100000100",
			267 => "1111111000010001001001",
			268 => "0001000111001100000100",
			269 => "0000011000010001001001",
			270 => "0000000000010001001001",
			271 => "0000010000111100000100",
			272 => "0000001000010001001001",
			273 => "1111111000010001001001",
			274 => "0000100101010100010000",
			275 => "0011000100011000000100",
			276 => "1111111000010001110101",
			277 => "0000011111001100001000",
			278 => "0011111011110100000100",
			279 => "0000000000010001110101",
			280 => "0000001000010001110101",
			281 => "1111111000010001110101",
			282 => "0000011110010100000100",
			283 => "0000001000010001110101",
			284 => "0000000000010001110101",
			285 => "0000100101010100010000",
			286 => "0001001111101100000100",
			287 => "1111111000010010100001",
			288 => "0000001010111100001000",
			289 => "0011000011011100000100",
			290 => "0000000000010010100001",
			291 => "0000001000010010100001",
			292 => "1111111000010010100001",
			293 => "0000011110010100000100",
			294 => "0000001000010010100001",
			295 => "0000000000010010100001",
			296 => "0000100101010100010000",
			297 => "0010101010100100001100",
			298 => "0001110111010000000100",
			299 => "1111111000010011001101",
			300 => "0001001000001100000100",
			301 => "0000000000010011001101",
			302 => "0000001000010011001101",
			303 => "1111111000010011001101",
			304 => "0000010000111100000100",
			305 => "0000001000010011001101",
			306 => "0000000000010011001101",
			307 => "0001000000101100001000",
			308 => "0011000100000100000100",
			309 => "1111111000010011111001",
			310 => "0000000000010011111001",
			311 => "0011000100011000000100",
			312 => "1111111000010011111001",
			313 => "0000011111001100001000",
			314 => "0000010010001100000100",
			315 => "0000000000010011111001",
			316 => "0000001000010011111001",
			317 => "0000000000010011111001",
			318 => "0011001001110100010000",
			319 => "0000101000101000000100",
			320 => "1111111000010100101101",
			321 => "0000000000001100000100",
			322 => "1111111000010100101101",
			323 => "0010101001101000000100",
			324 => "0000001000010100101101",
			325 => "0000000000010100101101",
			326 => "0000010000111100001000",
			327 => "0000001011010100000100",
			328 => "0000000000010100101101",
			329 => "0000001000010100101101",
			330 => "1111111000010100101101",
			331 => "0000101110111000010100",
			332 => "0000100101010100000100",
			333 => "1111111000010101100001",
			334 => "0011001111011100000100",
			335 => "0000011000010101100001",
			336 => "0011000100000100000100",
			337 => "1111111000010101100001",
			338 => "0011000001011000000100",
			339 => "0000001000010101100001",
			340 => "0000000000010101100001",
			341 => "0000010111101000000100",
			342 => "0000011000010101100001",
			343 => "1111111000010101100001",
			344 => "0011000100011000000100",
			345 => "0000000000010110001101",
			346 => "0001100010101100010000",
			347 => "0001101010011000000100",
			348 => "0000000000010110001101",
			349 => "0000110100000100000100",
			350 => "0000000000010110001101",
			351 => "0000101111010100000100",
			352 => "0000000000010110001101",
			353 => "0000000000010110001101",
			354 => "0000000000010110001101",
			355 => "0011000100011000000100",
			356 => "1111111000010111000001",
			357 => "0000011111001100010000",
			358 => "0001101010011000000100",
			359 => "0000000000010111000001",
			360 => "0000010010001100000100",
			361 => "0000000000010111000001",
			362 => "0000011111001100000100",
			363 => "0000001000010111000001",
			364 => "0000000000010111000001",
			365 => "0011001011011100000100",
			366 => "0000000000010111000001",
			367 => "0000000000010111000001",
			368 => "0000100101010100011000",
			369 => "0011000100011000000100",
			370 => "1111111000010111111101",
			371 => "0011101001100000010000",
			372 => "0001101010011000000100",
			373 => "1111111000010111111101",
			374 => "0001101011001100001000",
			375 => "0000101111010100000100",
			376 => "0000000000010111111101",
			377 => "0000001000010111111101",
			378 => "0000000000010111111101",
			379 => "1111111000010111111101",
			380 => "0010010100101100000100",
			381 => "0000001000010111111101",
			382 => "0000000000010111111101",
			383 => "0000100101010100011100",
			384 => "0011000100011000000100",
			385 => "1111111000011001001011",
			386 => "0011000100011000000100",
			387 => "0000000000011001001011",
			388 => "0011001001110100010000",
			389 => "0011001001110100000100",
			390 => "1111111000011001001011",
			391 => "0011001001110100000100",
			392 => "0000000000011001001011",
			393 => "0011001001110100000100",
			394 => "1111111000011001001011",
			395 => "0000000000011001001011",
			396 => "1111111000011001001011",
			397 => "0000010000111100001000",
			398 => "0011111001001100000100",
			399 => "0000001000011001001011",
			400 => "0000001000011001001011",
			401 => "1111111000011001001011",
			402 => "0000000000011001001101",
			403 => "0000000000011001010001",
			404 => "0000000000011001010101",
			405 => "0000000000011001011001",
			406 => "0000000000011001011101",
			407 => "0000000000011001100001",
			408 => "0000000000011001100101",
			409 => "0000000000011001101001",
			410 => "0000000000011001101101",
			411 => "0000000000011001110001",
			412 => "0000000000011001110101",
			413 => "0000000000011001111001",
			414 => "0000000000011001111101",
			415 => "0000000000011010000001",
			416 => "0000000000011010000101",
			417 => "0000000000011010001001",
			418 => "0000000000011010001101",
			419 => "0000000000011010010001",
			420 => "0000000000011010010101",
			421 => "0000000000011010011001",
			422 => "0000000000011010011101",
			423 => "0000000000011010100001",
			424 => "0000000000011010100101",
			425 => "0000000000011010101001",
			426 => "0000000000011010101101",
			427 => "0000000000011010110001",
			428 => "0000000000011010110101",
			429 => "0000000000011010111001",
			430 => "0000000000011010111101",
			431 => "0000000000011011000001",
			432 => "0000000000011011000101",
			433 => "0000000000011011001001",
			434 => "0000000000011011001101",
			435 => "0001001011001000000100",
			436 => "0000000000011011011001",
			437 => "0000000000011011011001",
			438 => "0001001011001000000100",
			439 => "0000000000011011100101",
			440 => "0000000000011011100101",
			441 => "0001110111010000000100",
			442 => "0000000000011011110001",
			443 => "0000000000011011110001",
			444 => "0000101110000000000100",
			445 => "0000000000011011111101",
			446 => "0000000000011011111101",
			447 => "0001111111011100000100",
			448 => "0000000000011100001001",
			449 => "0000000000011100001001",
			450 => "0001001011100100000100",
			451 => "0000000000011100010101",
			452 => "0000000000011100010101",
			453 => "0001110011100000000100",
			454 => "0000000000011100100001",
			455 => "0000000000011100100001",
			456 => "0001001011100100000100",
			457 => "0000000000011100101101",
			458 => "0000000000011100101101",
			459 => "0001000001100100000100",
			460 => "0000000000011100111001",
			461 => "0000000000011100111001",
			462 => "0001001011100100000100",
			463 => "0000000000011101000101",
			464 => "0000000000011101000101",
			465 => "0000100101010100000100",
			466 => "1111111000011101011001",
			467 => "0000010000111100000100",
			468 => "0000001000011101011001",
			469 => "1111111000011101011001",
			470 => "0011001001110100000100",
			471 => "0000000000011101101101",
			472 => "0000011101011100000100",
			473 => "0000000000011101101101",
			474 => "0000000000011101101101",
			475 => "0001111111011100000100",
			476 => "0000000000011110000001",
			477 => "0000011101011100000100",
			478 => "0000000000011110000001",
			479 => "0000000000011110000001",
			480 => "0011000100011000000100",
			481 => "0000000000011110010101",
			482 => "0000101111010100000100",
			483 => "0000000000011110010101",
			484 => "0000000000011110010101",
			485 => "0001110111010000001000",
			486 => "0001001111101100000100",
			487 => "0000000000011110110001",
			488 => "0000000000011110110001",
			489 => "0000010000111100000100",
			490 => "0000000000011110110001",
			491 => "0000000000011110110001",
			492 => "0000100101010100000100",
			493 => "1111111000011111001101",
			494 => "0000011110010100001000",
			495 => "0011111010110100000100",
			496 => "0000011000011111001101",
			497 => "0000010000011111001101",
			498 => "1111111000011111001101",
			499 => "0000100101010100000100",
			500 => "1111111000011111101001",
			501 => "0000010000111100001000",
			502 => "0011111001001100000100",
			503 => "0000010000011111101001",
			504 => "0000001000011111101001",
			505 => "1111111000011111101001",
			506 => "0010111010001100000100",
			507 => "1111111000100000000101",
			508 => "0000011111001100001000",
			509 => "0001010111100000000100",
			510 => "0000000000100000000101",
			511 => "0000000000100000000101",
			512 => "0000000000100000000101",
			513 => "0011000100011000000100",
			514 => "0000000000100000100001",
			515 => "0000101111010100000100",
			516 => "0000000000100000100001",
			517 => "0000110100000100000100",
			518 => "0000000000100000100001",
			519 => "0000000000100000100001",
			520 => "0001110011100000000100",
			521 => "0000000000100000111101",
			522 => "0000101111010100000100",
			523 => "0000000000100000111101",
			524 => "0000110100000100000100",
			525 => "0000000000100000111101",
			526 => "0000000000100000111101",
			527 => "0011000100011000000100",
			528 => "0000000000100001011001",
			529 => "0000101111010100000100",
			530 => "0000000000100001011001",
			531 => "0011010010001000000100",
			532 => "0000000000100001011001",
			533 => "0000000000100001011001",
			534 => "0010111001110100000100",
			535 => "0000000000100001110101",
			536 => "0000101111010100000100",
			537 => "0000000000100001110101",
			538 => "0011110100101000000100",
			539 => "0000000000100001110101",
			540 => "0000000000100001110101",
			541 => "0010111001110100000100",
			542 => "0000000000100010010001",
			543 => "0000101111010100000100",
			544 => "0000000000100010010001",
			545 => "0000110100000100000100",
			546 => "0000000000100010010001",
			547 => "0000000000100010010001",
			548 => "0000100101010100001100",
			549 => "0001111111011100000100",
			550 => "1111111000100010110101",
			551 => "0010110010001000000100",
			552 => "0000001000100010110101",
			553 => "1111111000100010110101",
			554 => "0000010000111100000100",
			555 => "0000001000100010110101",
			556 => "0000000000100010110101",
			557 => "0000100101010100001100",
			558 => "0010101010100100001000",
			559 => "0010000001010000000100",
			560 => "1111111000100011011001",
			561 => "0000001000100011011001",
			562 => "1111111000100011011001",
			563 => "0000010000111100000100",
			564 => "0000001000100011011001",
			565 => "0000000000100011011001",
			566 => "0011001001110100001100",
			567 => "0000101110000000000100",
			568 => "1111111000100011111101",
			569 => "0000101110000000000100",
			570 => "0000000000100011111101",
			571 => "0000000000100011111101",
			572 => "0000011101011100000100",
			573 => "0000001000100011111101",
			574 => "0000000000100011111101",
			575 => "0011001001110100001000",
			576 => "0001000100110000000100",
			577 => "1111111000100100100001",
			578 => "0000000000100100100001",
			579 => "0000011101011100001000",
			580 => "0000000101100100000100",
			581 => "0000001000100100100001",
			582 => "0000000000100100100001",
			583 => "0000000000100100100001",
			584 => "0001001011100100001000",
			585 => "0011111101001000000100",
			586 => "1111111000100101000101",
			587 => "0000000000100101000101",
			588 => "0010111001110100000100",
			589 => "0000000000100101000101",
			590 => "0000010010001100000100",
			591 => "0000000000100101000101",
			592 => "0000000000100101000101",
			593 => "0011000100011000000100",
			594 => "1111111000100101101001",
			595 => "0000011111001100001000",
			596 => "0001111111011100000100",
			597 => "0000000000100101101001",
			598 => "0000001000100101101001",
			599 => "0011001011011100000100",
			600 => "0000000000100101101001",
			601 => "0000000000100101101001",
			602 => "0011000100011000000100",
			603 => "1111111000100110001101",
			604 => "0000011111001100001000",
			605 => "0011110100101000000100",
			606 => "0000000000100110001101",
			607 => "0000000000100110001101",
			608 => "0000001101111000000100",
			609 => "0000000000100110001101",
			610 => "0000000000100110001101",
			611 => "0001001011001000000100",
			612 => "1111111000100110110001",
			613 => "0011000100011000000100",
			614 => "0000000000100110110001",
			615 => "0000010000111100001000",
			616 => "0000010010001100000100",
			617 => "0000000000100110110001",
			618 => "0000001000100110110001",
			619 => "0000000000100110110001",
			620 => "0001001011001000000100",
			621 => "1111111000100111010101",
			622 => "0010111001110100000100",
			623 => "0000000000100111010101",
			624 => "0000010000111100001000",
			625 => "0000010010001100000100",
			626 => "0000000000100111010101",
			627 => "0000000000100111010101",
			628 => "0000000000100111010101",
			629 => "0001001011001000000100",
			630 => "0000000000100111111001",
			631 => "0011000100011000000100",
			632 => "0000000000100111111001",
			633 => "0010011000010000001000",
			634 => "0000110100000100000100",
			635 => "0000000000100111111001",
			636 => "0000000000100111111001",
			637 => "0000000000100111111001",
			638 => "0001110011100000000100",
			639 => "0000000000101000011101",
			640 => "0000010000111100001100",
			641 => "0000101111010100000100",
			642 => "0000000000101000011101",
			643 => "0000010010001100000100",
			644 => "0000000000101000011101",
			645 => "0000000000101000011101",
			646 => "0000000000101000011101",
			647 => "0011000100011000000100",
			648 => "0000000000101001000001",
			649 => "0000010000111100001100",
			650 => "0001101010011000000100",
			651 => "0000000000101001000001",
			652 => "0000000101100100000100",
			653 => "0000000000101001000001",
			654 => "0000000000101001000001",
			655 => "0000000000101001000001",
			656 => "0011000100011000000100",
			657 => "0000000000101001100101",
			658 => "0000010000111100001100",
			659 => "0011110100101000000100",
			660 => "0000000000101001100101",
			661 => "0001101010011000000100",
			662 => "0000000000101001100101",
			663 => "0000000000101001100101",
			664 => "0000000000101001100101",
			665 => "0000100101010100010000",
			666 => "0011000100011000000100",
			667 => "1111111000101010010001",
			668 => "0000011111001100001000",
			669 => "0000111100101100000100",
			670 => "0000000000101010010001",
			671 => "0000010000101010010001",
			672 => "1111111000101010010001",
			673 => "0000010000111100000100",
			674 => "0000001000101010010001",
			675 => "1111111000101010010001",
			676 => "0011110010111000010000",
			677 => "0011000100011000000100",
			678 => "1111111000101010111101",
			679 => "0000011111001100001000",
			680 => "0000010010001100000100",
			681 => "0000000000101010111101",
			682 => "0000001000101010111101",
			683 => "1111111000101010111101",
			684 => "0000011011111100000100",
			685 => "0000001000101010111101",
			686 => "0000000000101010111101",
			687 => "0000100101010100010000",
			688 => "0000000000001100000100",
			689 => "1111111000101011101001",
			690 => "0010000010011000001000",
			691 => "0011001010000000000100",
			692 => "0000000000101011101001",
			693 => "0000001000101011101001",
			694 => "1111111000101011101001",
			695 => "0000011110010100000100",
			696 => "0000001000101011101001",
			697 => "0000000000101011101001",
			698 => "0001000000101100001000",
			699 => "0000100101010100000100",
			700 => "1111111000101100010101",
			701 => "0000000000101100010101",
			702 => "0011000100011000000100",
			703 => "1111111000101100010101",
			704 => "0000011111001100001000",
			705 => "0000010010001100000100",
			706 => "0000000000101100010101",
			707 => "0000001000101100010101",
			708 => "0000000000101100010101",
			709 => "0000100101010100010000",
			710 => "0001000000000100000100",
			711 => "1111111000101101000001",
			712 => "0010000010011000001000",
			713 => "0000101100111000000100",
			714 => "0000000000101101000001",
			715 => "0000000000101101000001",
			716 => "0000000000101101000001",
			717 => "0010011000010000000100",
			718 => "0000001000101101000001",
			719 => "0000000000101101000001",
			720 => "0011001001110100010000",
			721 => "0000101000101000000100",
			722 => "1111111000101101110101",
			723 => "0000000000001100000100",
			724 => "0000000000101101110101",
			725 => "0010101001101000000100",
			726 => "0000000000101101110101",
			727 => "0000000000101101110101",
			728 => "0000010000111100001000",
			729 => "0000001011010100000100",
			730 => "0000000000101101110101",
			731 => "0000001000101101110101",
			732 => "1111111000101101110101",
			733 => "0001001011001000000100",
			734 => "1111111000101110100001",
			735 => "0011000100011000000100",
			736 => "0000000000101110100001",
			737 => "0000010000111100001100",
			738 => "0000101000101000000100",
			739 => "0000000000101110100001",
			740 => "0001001111110100000100",
			741 => "0000000000101110100001",
			742 => "0000000000101110100001",
			743 => "0000000000101110100001",
			744 => "0011000100011000000100",
			745 => "1111111000101111010101",
			746 => "0000011111001100010000",
			747 => "0001101010011000000100",
			748 => "0000000000101111010101",
			749 => "0000010010001100000100",
			750 => "0000000000101111010101",
			751 => "0000011111001100000100",
			752 => "0000001000101111010101",
			753 => "0000000000101111010101",
			754 => "0011001011011100000100",
			755 => "1111111000101111010101",
			756 => "0000000000101111010101",
			757 => "0000100101010100011000",
			758 => "0011000100011000000100",
			759 => "1111111000110000010001",
			760 => "0000000000001100001100",
			761 => "0011101001100000001000",
			762 => "0011110110111100000100",
			763 => "1111111000110000010001",
			764 => "0000010000110000010001",
			765 => "1111111000110000010001",
			766 => "0011111011011100000100",
			767 => "0000000000110000010001",
			768 => "0000001000110000010001",
			769 => "0000010000111100000100",
			770 => "0000001000110000010001",
			771 => "1111111000110000010001",
			772 => "0000100101010100011100",
			773 => "0011000100011000000100",
			774 => "1111111000110001010101",
			775 => "0000000000001100010000",
			776 => "0011101001100000001100",
			777 => "0000110110111100000100",
			778 => "1111111000110001010101",
			779 => "0011100110010000000100",
			780 => "0000000000110001010101",
			781 => "0000100000110001010101",
			782 => "1111111000110001010101",
			783 => "0011111011011100000100",
			784 => "0000000000110001010101",
			785 => "0000010000110001010101",
			786 => "0000010000111100000100",
			787 => "0000001000110001010101",
			788 => "1111111000110001010101",
			789 => "0000100101010100100000",
			790 => "0011000100011000000100",
			791 => "1111111000110010100011",
			792 => "0000000000001100010100",
			793 => "0010111011011100010000",
			794 => "0010111011011100000100",
			795 => "1111111000110010100011",
			796 => "0010101010100100001000",
			797 => "0001001110110100000100",
			798 => "0000000000110010100011",
			799 => "0000011000110010100011",
			800 => "0000000000110010100011",
			801 => "1111111000110010100011",
			802 => "0011111011011100000100",
			803 => "0000000000110010100011",
			804 => "0000010000110010100011",
			805 => "0000010000111100000100",
			806 => "0000001000110010100011",
			807 => "1111111000110010100011",
			808 => "0000000000110010100101",
			809 => "0000000000110010101001",
			810 => "0000000000110010101101",
			811 => "0000000000110010110001",
			812 => "0000000000110010110101",
			813 => "0000000000110010111001",
			814 => "0000000000110010111101",
			815 => "0000000000110011000001",
			816 => "0000000000110011000101",
			817 => "0000000000110011001001",
			818 => "0000000000110011001101",
			819 => "0000000000110011010001",
			820 => "0000000000110011010101",
			821 => "0000000000110011011001",
			822 => "0000000000110011011101",
			823 => "0000000000110011100001",
			824 => "0000000000110011100101",
			825 => "0000000000110011101001",
			826 => "0000000000110011101101",
			827 => "0000000000110011110001",
			828 => "0000000000110011110101",
			829 => "0000000000110011111001",
			830 => "0000000000110011111101",
			831 => "0000000000110100000001",
			832 => "0000000000110100000101",
			833 => "0000000000110100001001",
			834 => "0000000000110100001101",
			835 => "0000000000110100010001",
			836 => "0000000000110100010101",
			837 => "0000000000110100011001",
			838 => "0000000000110100011101",
			839 => "0000000000110100100001",
			840 => "0001001011001000000100",
			841 => "0000000000110100101101",
			842 => "0000000000110100101101",
			843 => "0001001011001000000100",
			844 => "0000000000110100111001",
			845 => "0000000000110100111001",
			846 => "0001001011001000000100",
			847 => "0000000000110101000101",
			848 => "0000000000110101000101",
			849 => "0001110111010000000100",
			850 => "0000000000110101010001",
			851 => "0000000000110101010001",
			852 => "0001001011001000000100",
			853 => "0000000000110101011101",
			854 => "0000000000110101011101",
			855 => "0001111111011100000100",
			856 => "0000000000110101101001",
			857 => "0000000000110101101001",
			858 => "0001001011100100000100",
			859 => "0000000000110101110101",
			860 => "0000000000110101110101",
			861 => "0001001011100100000100",
			862 => "0000000000110110000001",
			863 => "0000000000110110000001",
			864 => "0001000001100100000100",
			865 => "0000000000110110001101",
			866 => "0000000000110110001101",
			867 => "0001001011100100000100",
			868 => "0000000000110110011001",
			869 => "0000000000110110011001",
			870 => "0011000100011000000100",
			871 => "0000000000110110100101",
			872 => "0000000000110110100101",
			873 => "0000100101010100000100",
			874 => "1111111000110110111001",
			875 => "0010011000010000000100",
			876 => "0000001000110110111001",
			877 => "1111111000110110111001",
			878 => "0001111111011100000100",
			879 => "0000000000110111001101",
			880 => "0000011101011100000100",
			881 => "0000000000110111001101",
			882 => "0000000000110111001101",
			883 => "0011000100011000000100",
			884 => "0000000000110111100001",
			885 => "0011110100101000000100",
			886 => "0000000000110111100001",
			887 => "0000000000110111100001",
			888 => "0000100101010100001000",
			889 => "0000000001111100000100",
			890 => "1111111000110111111101",
			891 => "0000000000110111111101",
			892 => "0000011110010100000100",
			893 => "0000000000110111111101",
			894 => "0000000000110111111101",
			895 => "0001110111010000001000",
			896 => "0001001111101100000100",
			897 => "0000000000111000011001",
			898 => "0000000000111000011001",
			899 => "0000010000111100000100",
			900 => "0000000000111000011001",
			901 => "0000000000111000011001",
			902 => "0000100101010100000100",
			903 => "1111111000111000110101",
			904 => "0000010000111100001000",
			905 => "0001100101010000000100",
			906 => "0000010000111000110101",
			907 => "0000001000111000110101",
			908 => "1111111000111000110101",
			909 => "0011000100011000000100",
			910 => "1111111000111001010001",
			911 => "0000011111001100001000",
			912 => "0001001111110100000100",
			913 => "0000000000111001010001",
			914 => "0000000000111001010001",
			915 => "0000000000111001010001",
			916 => "0000001001110000001100",
			917 => "0011000111010000001000",
			918 => "0000100011110100000100",
			919 => "0000000000111001101101",
			920 => "0000000000111001101101",
			921 => "0000000000111001101101",
			922 => "0000000000111001101101",
			923 => "0011000100011000000100",
			924 => "0000000000111010001001",
			925 => "0000101111010100000100",
			926 => "0000000000111010001001",
			927 => "0000110100000100000100",
			928 => "0000000000111010001001",
			929 => "0000000000111010001001",
			930 => "0011000100011000000100",
			931 => "0000000000111010100101",
			932 => "0000101111010100000100",
			933 => "0000000000111010100101",
			934 => "0000110100000100000100",
			935 => "0000000000111010100101",
			936 => "0000000000111010100101",
			937 => "0011000100011000000100",
			938 => "0000000000111011000001",
			939 => "0011110100101000000100",
			940 => "0000000000111011000001",
			941 => "0000101111010100000100",
			942 => "0000000000111011000001",
			943 => "0000000000111011000001",
			944 => "0011000100011000000100",
			945 => "0000000000111011011101",
			946 => "0011110100101000000100",
			947 => "0000000000111011011101",
			948 => "0000101111010100000100",
			949 => "0000000000111011011101",
			950 => "0000000000111011011101",
			951 => "0000100101010100001100",
			952 => "0011000100011000000100",
			953 => "1111111000111100000001",
			954 => "0011000100011000000100",
			955 => "0000000000111100000001",
			956 => "1111111000111100000001",
			957 => "0000010000111100000100",
			958 => "0000001000111100000001",
			959 => "1111111000111100000001",
			960 => "0000100101010100001100",
			961 => "0001111111011100000100",
			962 => "1111111000111100100101",
			963 => "0010110010001000000100",
			964 => "0000001000111100100101",
			965 => "1111111000111100100101",
			966 => "0000010000111100000100",
			967 => "0000001000111100100101",
			968 => "0000000000111100100101",
			969 => "0011001001110100001100",
			970 => "0000101110000000000100",
			971 => "1111111000111101001001",
			972 => "0000101110000000000100",
			973 => "0000000000111101001001",
			974 => "0000000000111101001001",
			975 => "0000011101011100000100",
			976 => "0000001000111101001001",
			977 => "1111111000111101001001",
			978 => "0011001001110100001000",
			979 => "0001000100110000000100",
			980 => "1111111000111101101101",
			981 => "0000000000111101101101",
			982 => "0000011101011100001000",
			983 => "0000000101100100000100",
			984 => "0000001000111101101101",
			985 => "0000000000111101101101",
			986 => "0000000000111101101101",
			987 => "0001111111011100001000",
			988 => "0001001111101100000100",
			989 => "1111111000111110010001",
			990 => "0000000000111110010001",
			991 => "0000010000111100001000",
			992 => "0000001011010100000100",
			993 => "0000000000111110010001",
			994 => "0000001000111110010001",
			995 => "0000000000111110010001",
			996 => "0001111111011100001000",
			997 => "0001001111101100000100",
			998 => "1111111000111110110101",
			999 => "0000000000111110110101",
			1000 => "0010010100111100001000",
			1001 => "0000001011010100000100",
			1002 => "0000000000111110110101",
			1003 => "0000000000111110110101",
			1004 => "0000000000111110110101",
			1005 => "0011000100011000000100",
			1006 => "1111111000111111011001",
			1007 => "0000011111001100001000",
			1008 => "0011110100101000000100",
			1009 => "0000000000111111011001",
			1010 => "0000000000111111011001",
			1011 => "0000100001001100000100",
			1012 => "0000000000111111011001",
			1013 => "0000000000111111011001",
			1014 => "0011000100011000000100",
			1015 => "1111111000111111111101",
			1016 => "0010011010011000001000",
			1017 => "0001001111110100000100",
			1018 => "0000000000111111111101",
			1019 => "0000000000111111111101",
			1020 => "0010010100111100000100",
			1021 => "0000000000111111111101",
			1022 => "0000000000111111111101",
			1023 => "0001001011001000000100",
			1024 => "1111111001000000100001",
			1025 => "0011000100011000000100",
			1026 => "0000000001000000100001",
			1027 => "0000010000111100001000",
			1028 => "0000010010001100000100",
			1029 => "0000000001000000100001",
			1030 => "0000001001000000100001",
			1031 => "0000000001000000100001",
			1032 => "0011000100011000000100",
			1033 => "1111111001000001000101",
			1034 => "0000011111001100001100",
			1035 => "0001101010011000000100",
			1036 => "0000000001000001000101",
			1037 => "0000000101110100000100",
			1038 => "0000000001000001000101",
			1039 => "0000000001000001000101",
			1040 => "0000000001000001000101",
			1041 => "0001001011001000000100",
			1042 => "0000000001000001101001",
			1043 => "0001110011100000000100",
			1044 => "0000000001000001101001",
			1045 => "0000010000111100001000",
			1046 => "0000010010001100000100",
			1047 => "0000000001000001101001",
			1048 => "0000000001000001101001",
			1049 => "0000000001000001101001",
			1050 => "0011000100011000000100",
			1051 => "0000000001000010001101",
			1052 => "0000010000111100001100",
			1053 => "0000101111010100000100",
			1054 => "0000000001000010001101",
			1055 => "0000000101110100000100",
			1056 => "0000000001000010001101",
			1057 => "0000000001000010001101",
			1058 => "0000000001000010001101",
			1059 => "0011000100011000000100",
			1060 => "0000000001000010110001",
			1061 => "0000010000111100001100",
			1062 => "0000001011010100000100",
			1063 => "0000000001000010110001",
			1064 => "0000010010001100000100",
			1065 => "0000000001000010110001",
			1066 => "0000000001000010110001",
			1067 => "0000000001000010110001",
			1068 => "0000100101010100010000",
			1069 => "0011000100011000000100",
			1070 => "1111111001000011011101",
			1071 => "0000000110000100000100",
			1072 => "1111111001000011011101",
			1073 => "0010001001110000000100",
			1074 => "0000111001000011011101",
			1075 => "0000000001000011011101",
			1076 => "0000010000111100000100",
			1077 => "0000001001000011011101",
			1078 => "1111111001000011011101",
			1079 => "0000100101010100010000",
			1080 => "0011000100011000000100",
			1081 => "1111111001000100001001",
			1082 => "0000011111001100001000",
			1083 => "0001101010011000000100",
			1084 => "0000000001000100001001",
			1085 => "0000001001000100001001",
			1086 => "1111111001000100001001",
			1087 => "0000010000111100000100",
			1088 => "0000001001000100001001",
			1089 => "1111111001000100001001",
			1090 => "0000100101010100010000",
			1091 => "0001001111101100000100",
			1092 => "1111111001000100110101",
			1093 => "0010000010111100001000",
			1094 => "0000100110100000000100",
			1095 => "0000000001000100110101",
			1096 => "0000001001000100110101",
			1097 => "1111111001000100110101",
			1098 => "0000011110010100000100",
			1099 => "0000001001000100110101",
			1100 => "0000000001000100110101",
			1101 => "0000100101010100010000",
			1102 => "0010101010100100001100",
			1103 => "0001110111010000000100",
			1104 => "1111111001000101100001",
			1105 => "0001001000001100000100",
			1106 => "0000000001000101100001",
			1107 => "0000001001000101100001",
			1108 => "1111111001000101100001",
			1109 => "0000010000111100000100",
			1110 => "0000001001000101100001",
			1111 => "0000000001000101100001",
			1112 => "0000100101010100010000",
			1113 => "0010001000110000000100",
			1114 => "1111111001000110001101",
			1115 => "0011000100011000000100",
			1116 => "1111111001000110001101",
			1117 => "0000100001011100000100",
			1118 => "0000000001000110001101",
			1119 => "0000001001000110001101",
			1120 => "0000010000111100000100",
			1121 => "0000001001000110001101",
			1122 => "0000000001000110001101",
			1123 => "0001111111011100001000",
			1124 => "0001001111101100000100",
			1125 => "1111111001000110111001",
			1126 => "0000000001000110111001",
			1127 => "0011001001110100000100",
			1128 => "0000000001000110111001",
			1129 => "0001100010101100001000",
			1130 => "0000001011010100000100",
			1131 => "0000000001000110111001",
			1132 => "0000000001000110111001",
			1133 => "0000000001000110111001",
			1134 => "0011001001110100010000",
			1135 => "0000101000101000000100",
			1136 => "1111111001000111101101",
			1137 => "0001000100110000000100",
			1138 => "0000000001000111101101",
			1139 => "0010101011010100000100",
			1140 => "0000000001000111101101",
			1141 => "0000000001000111101101",
			1142 => "0000011101011100000100",
			1143 => "0000001001000111101101",
			1144 => "0000010000111100000100",
			1145 => "0000000001000111101101",
			1146 => "1111111001000111101101",
			1147 => "0001001011001000000100",
			1148 => "1111111001001000011001",
			1149 => "0011000100011000000100",
			1150 => "0000000001001000011001",
			1151 => "0000010000111100001100",
			1152 => "0000101000101000000100",
			1153 => "0000000001001000011001",
			1154 => "0001001111110100000100",
			1155 => "0000000001001000011001",
			1156 => "0000000001001000011001",
			1157 => "0000000001001000011001",
			1158 => "0011000100011000000100",
			1159 => "1111111001001001001101",
			1160 => "0000011111001100010000",
			1161 => "0001101010011000000100",
			1162 => "0000000001001001001101",
			1163 => "0000010010001100000100",
			1164 => "0000000001001001001101",
			1165 => "0000011111001100000100",
			1166 => "0000001001001001001101",
			1167 => "0000000001001001001101",
			1168 => "0011001011011100000100",
			1169 => "1111111001001001001101",
			1170 => "0000000001001001001101",
			1171 => "0011110010111000011000",
			1172 => "0001001011100100000100",
			1173 => "1111111001001010001001",
			1174 => "0011110100101000000100",
			1175 => "1111111001001010001001",
			1176 => "0001101001100100000100",
			1177 => "0000011001001010001001",
			1178 => "0000010111100100000100",
			1179 => "0000001001001010001001",
			1180 => "0000000011011100000100",
			1181 => "0000000001001010001001",
			1182 => "0000000001001010001001",
			1183 => "0000010000111100000100",
			1184 => "0000001001001010001001",
			1185 => "1111111001001010001001",
			1186 => "0000100101010100011100",
			1187 => "0011000100011000000100",
			1188 => "1111111001001011010101",
			1189 => "0011000100011000000100",
			1190 => "0000000001001011010101",
			1191 => "0011001001110100010000",
			1192 => "0011001001110100000100",
			1193 => "1111111001001011010101",
			1194 => "0011001001110100000100",
			1195 => "0000001001001011010101",
			1196 => "0011001001110100000100",
			1197 => "1111111001001011010101",
			1198 => "0000000001001011010101",
			1199 => "1111111001001011010101",
			1200 => "0010011000010000001000",
			1201 => "0011111001001100000100",
			1202 => "0000010001001011010101",
			1203 => "0000001001001011010101",
			1204 => "1111111001001011010101",
			1205 => "0000110010111000101000",
			1206 => "0000110011110000100000",
			1207 => "0001101000010000010100",
			1208 => "0011011010000100010000",
			1209 => "0000110101000000000100",
			1210 => "1111111001001100110011",
			1211 => "0000111100001100001000",
			1212 => "0000111100001100000100",
			1213 => "0000000001001100110011",
			1214 => "0000000001001100110011",
			1215 => "1111111001001100110011",
			1216 => "0000000001001100110011",
			1217 => "0000011111001100001000",
			1218 => "0000111101101100000100",
			1219 => "1111111001001100110011",
			1220 => "0000010001001100110011",
			1221 => "1111111001001100110011",
			1222 => "0000000111111000000100",
			1223 => "1111111001001100110011",
			1224 => "0000010001001100110011",
			1225 => "0000011110010100000100",
			1226 => "0000010001001100110011",
			1227 => "1111111001001100110011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(402, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(808, initial_addr_3'length));
	end generate gen_rom_5;

	gen_rom_6: if SELECT_ROM = 6 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000000000000001110101",
			29 => "0000000000000001111001",
			30 => "0000100111100000000100",
			31 => "0000000000000010000101",
			32 => "0000000000000010000101",
			33 => "0000111010101100000100",
			34 => "0000000000000010010001",
			35 => "0000000000000010010001",
			36 => "0000101100100100000100",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0000101100100100000100",
			40 => "0000000000000010101001",
			41 => "0000000000000010101001",
			42 => "0001101101111100001000",
			43 => "0001101011111100000100",
			44 => "0000000000000010111101",
			45 => "0000000000000010111101",
			46 => "0000000000000010111101",
			47 => "0001101101111100001000",
			48 => "0001101011111100000100",
			49 => "0000000000000011010001",
			50 => "0000000000000011010001",
			51 => "0000000000000011010001",
			52 => "0001001011100100001000",
			53 => "0011011001110100000100",
			54 => "0000000000000011100101",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0001101101111100001000",
			58 => "0001101011111100000100",
			59 => "0000000000000011111001",
			60 => "0000000000000011111001",
			61 => "0000000000000011111001",
			62 => "0001101101111100001000",
			63 => "0001101011111100000100",
			64 => "0000000000000100001101",
			65 => "0000000000000100001101",
			66 => "0000000000000100001101",
			67 => "0000101100100100000100",
			68 => "0000000000000100100001",
			69 => "0000110111000000000100",
			70 => "0000000000000100100001",
			71 => "0000000000000100100001",
			72 => "0001101101111100001000",
			73 => "0001101011111100000100",
			74 => "0000000000000100110101",
			75 => "0000000000000100110101",
			76 => "0000000000000100110101",
			77 => "0001101101111100001000",
			78 => "0001101011111100000100",
			79 => "0000000000000101001001",
			80 => "0000000000000101001001",
			81 => "0000000000000101001001",
			82 => "0001101101111100001000",
			83 => "0001101011111100000100",
			84 => "0000000000000101011101",
			85 => "0000000000000101011101",
			86 => "0000000000000101011101",
			87 => "0001101101111100001000",
			88 => "0001101011111100000100",
			89 => "0000000000000101110001",
			90 => "0000000000000101110001",
			91 => "0000000000000101110001",
			92 => "0001101101111100001000",
			93 => "0001101011111100000100",
			94 => "0000000000000110001101",
			95 => "0000000000000110001101",
			96 => "0000100111100000000100",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0001101101111100001100",
			100 => "0000100111100000001000",
			101 => "0001101011111100000100",
			102 => "0000000000000110101001",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0000100111100000001100",
			107 => "0001101101111100001000",
			108 => "0001101011111100000100",
			109 => "0000000000000111001101",
			110 => "0000000000000111001101",
			111 => "0000000000000111001101",
			112 => "0000101000001100000100",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0011011001110100001000",
			116 => "0000110001110100000100",
			117 => "0000000000000111110001",
			118 => "0000000000000111110001",
			119 => "0011101100101100000100",
			120 => "0000000000000111110001",
			121 => "0011100111011000000100",
			122 => "0000000000000111110001",
			123 => "0000000000000111110001",
			124 => "0001000011011000000100",
			125 => "0000000000001000010101",
			126 => "0011000011011100001100",
			127 => "0001101101111100001000",
			128 => "0001100111101000000100",
			129 => "0000000000001000010101",
			130 => "0000000000001000010101",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0001101101111100010000",
			134 => "0000110100011000000100",
			135 => "0000000000001000111001",
			136 => "0001101011111100000100",
			137 => "0000000000001000111001",
			138 => "0011011001110100000100",
			139 => "0000000000001000111001",
			140 => "0000000000001000111001",
			141 => "0000000000001000111001",
			142 => "0001101101111100010000",
			143 => "0001101011111100000100",
			144 => "0000000000001001100101",
			145 => "0010000100010100001000",
			146 => "0010001001000100000100",
			147 => "0000000000001001100101",
			148 => "0000000000001001100101",
			149 => "0000000000001001100101",
			150 => "0000110111000100000100",
			151 => "0000000000001001100101",
			152 => "0000000000001001100101",
			153 => "0001101101111100010000",
			154 => "0000110100011000001000",
			155 => "0001000100111000000100",
			156 => "0000000000001010011001",
			157 => "0000000000001010011001",
			158 => "0001001111101000000100",
			159 => "0000000000001010011001",
			160 => "0000000000001010011001",
			161 => "0001001010010000001000",
			162 => "0001010001101000000100",
			163 => "0000000000001010011001",
			164 => "0000000000001010011001",
			165 => "0000000000001010011001",
			166 => "0011100001010100010000",
			167 => "0010000100000000001100",
			168 => "0011110001111100001000",
			169 => "0001001110001000000100",
			170 => "0000001000001011010101",
			171 => "0000010000001011010101",
			172 => "1111111000001011010101",
			173 => "1111111000001011010101",
			174 => "0011110001111100001100",
			175 => "0001110000101000001000",
			176 => "0000011100100000000100",
			177 => "0000010000001011010101",
			178 => "1111111000001011010101",
			179 => "1111111000001011010101",
			180 => "1111111000001011010101",
			181 => "0000100111100000010100",
			182 => "0000011100110100010000",
			183 => "0001101101111100001100",
			184 => "0001101011111100000100",
			185 => "0000000000001100001001",
			186 => "0000000001001000000100",
			187 => "0000000000001100001001",
			188 => "0000000000001100001001",
			189 => "0000000000001100001001",
			190 => "0000000000001100001001",
			191 => "0000110111000000000100",
			192 => "0000000000001100001001",
			193 => "0000000000001100001001",
			194 => "0001000011011000000100",
			195 => "1111111000001100110101",
			196 => "0001101101111100010000",
			197 => "0001111110001100001100",
			198 => "0001101110010100000100",
			199 => "0000000000001100110101",
			200 => "0000101110110100000100",
			201 => "0000001000001100110101",
			202 => "0000000000001100110101",
			203 => "0000000000001100110101",
			204 => "0000000000001100110101",
			205 => "0001101101111100010100",
			206 => "0011011010111100000100",
			207 => "0000000000001101100001",
			208 => "0000101110101000000100",
			209 => "0000000000001101100001",
			210 => "0000111100001000000100",
			211 => "0000000000001101100001",
			212 => "0010110101100100000100",
			213 => "0000000000001101100001",
			214 => "0000000000001101100001",
			215 => "0000000000001101100001",
			216 => "0000010000011000010100",
			217 => "0001011010111000010000",
			218 => "0001101101111100001100",
			219 => "0001100111101000000100",
			220 => "0000000000001110100101",
			221 => "0000101100010100000100",
			222 => "0000001000001110100101",
			223 => "0000000000001110100101",
			224 => "0000000000001110100101",
			225 => "0000000000001110100101",
			226 => "0011011010011100000100",
			227 => "1111111000001110100101",
			228 => "0011001000111000001000",
			229 => "0011100010001000000100",
			230 => "0000001000001110100101",
			231 => "0000000000001110100101",
			232 => "1111111000001110100101",
			233 => "0001000011011000000100",
			234 => "1111111000001111011001",
			235 => "0011000011011100010100",
			236 => "0010111100001000001100",
			237 => "0010010000011000001000",
			238 => "0011111010111000000100",
			239 => "0000000000001111011001",
			240 => "0000000000001111011001",
			241 => "0000000000001111011001",
			242 => "0001101100011000000100",
			243 => "0000000000001111011001",
			244 => "0000000000001111011001",
			245 => "0000000000001111011001",
			246 => "0001001011100100011000",
			247 => "0010000110011000001000",
			248 => "0000100111010100000100",
			249 => "1111111000010000100101",
			250 => "0000001000010000100101",
			251 => "0001001101110100000100",
			252 => "1111111000010000100101",
			253 => "0011011001110100000100",
			254 => "1111111000010000100101",
			255 => "0011010001011000000100",
			256 => "0000000000010000100101",
			257 => "0000000000010000100101",
			258 => "0010111001110000001100",
			259 => "0000100011001000001000",
			260 => "0001101110010100000100",
			261 => "0000000000010000100101",
			262 => "0000001000010000100101",
			263 => "0000000000010000100101",
			264 => "1111111000010000100101",
			265 => "0011011001110100011000",
			266 => "0001001011100100001000",
			267 => "0011110011011100000100",
			268 => "0000000000010001110001",
			269 => "0000000000010001110001",
			270 => "0000100011001000001100",
			271 => "0010100010101000001000",
			272 => "0010100101000100000100",
			273 => "0000000000010001110001",
			274 => "0000000000010001110001",
			275 => "0000000000010001110001",
			276 => "0000000000010001110001",
			277 => "0010100110011000001100",
			278 => "0001001111101000000100",
			279 => "0000000000010001110001",
			280 => "0000011101101000000100",
			281 => "0000000000010001110001",
			282 => "0000000000010001110001",
			283 => "0000000000010001110001",
			284 => "0001101101111100011100",
			285 => "0011011010111100010000",
			286 => "0011111010111000001100",
			287 => "0001000000101100000100",
			288 => "0000000000010010101101",
			289 => "0001101110010100000100",
			290 => "0000000000010010101101",
			291 => "0000000000010010101101",
			292 => "0000000000010010101101",
			293 => "0010011110100000000100",
			294 => "0000000000010010101101",
			295 => "0001001111101000000100",
			296 => "0000000000010010101101",
			297 => "0000001000010010101101",
			298 => "0000000000010010101101",
			299 => "0001101101111100011100",
			300 => "0011011010111100001100",
			301 => "0011111010111000001000",
			302 => "0010100110011100000100",
			303 => "0000000000010011101001",
			304 => "0000000000010011101001",
			305 => "0000000000010011101001",
			306 => "0001001011110000000100",
			307 => "0000000000010011101001",
			308 => "0010011110100000000100",
			309 => "0000000000010011101001",
			310 => "0001100001111000000100",
			311 => "0000000000010011101001",
			312 => "0000000000010011101001",
			313 => "0000000000010011101001",
			314 => "0001100001111000011100",
			315 => "0000110111000000001000",
			316 => "0001100111101000000100",
			317 => "0000000000010100111101",
			318 => "0000000000010100111101",
			319 => "0000110100011000001100",
			320 => "0011110101101100000100",
			321 => "0000000000010100111101",
			322 => "0000011110011100000100",
			323 => "0000000000010100111101",
			324 => "0000000000010100111101",
			325 => "0010101010100100000100",
			326 => "0000000000010100111101",
			327 => "0000000000010100111101",
			328 => "0001010100000100001000",
			329 => "0000110111000100000100",
			330 => "0000000000010100111101",
			331 => "1111111000010100111101",
			332 => "0010110111001000000100",
			333 => "0000000000010100111101",
			334 => "0000000000010100111101",
			335 => "0001000011011000001100",
			336 => "0010000110011000001000",
			337 => "0000001001101000000100",
			338 => "0000000000010110000001",
			339 => "0000001000010110000001",
			340 => "1111111000010110000001",
			341 => "0001101101111100010100",
			342 => "0001111110001100010000",
			343 => "0001100111101000000100",
			344 => "0000000000010110000001",
			345 => "0000010000011000000100",
			346 => "0000001000010110000001",
			347 => "0001000000100000000100",
			348 => "0000000000010110000001",
			349 => "0000000000010110000001",
			350 => "0000000000010110000001",
			351 => "1111111000010110000001",
			352 => "0001000011011000000100",
			353 => "0000000000010110110101",
			354 => "0011000011011100010100",
			355 => "0001101101111100010000",
			356 => "0001101110010100000100",
			357 => "0000000000010110110101",
			358 => "0000101100000000001000",
			359 => "0010000100010100000100",
			360 => "0000000000010110110101",
			361 => "0000000000010110110101",
			362 => "0000000000010110110101",
			363 => "0000000000010110110101",
			364 => "0000000000010110110101",
			365 => "0001101101111100011100",
			366 => "0000110100011000010100",
			367 => "0000010000011000010000",
			368 => "0001010011100000001100",
			369 => "0001101110010100000100",
			370 => "0000000000010111110001",
			371 => "0000100011001000000100",
			372 => "0000000000010111110001",
			373 => "0000000000010111110001",
			374 => "0000000000010111110001",
			375 => "1111111000010111110001",
			376 => "0001001111101000000100",
			377 => "0000000000010111110001",
			378 => "0000001000010111110001",
			379 => "1111111000010111110001",
			380 => "0010110110000100010100",
			381 => "0001000101100000001000",
			382 => "0000011100100000000100",
			383 => "0000000000011001000101",
			384 => "1111111000011001000101",
			385 => "0000100011001000001000",
			386 => "0010001011000100000100",
			387 => "0000001000011001000101",
			388 => "0000000000011001000101",
			389 => "0000000000011001000101",
			390 => "0011000100001000010100",
			391 => "0010100001010000010000",
			392 => "0001001111101000000100",
			393 => "0000000000011001000101",
			394 => "0000011101101000001000",
			395 => "0011000100000000000100",
			396 => "0000000000011001000101",
			397 => "0000001000011001000101",
			398 => "0000000000011001000101",
			399 => "0000000000011001000101",
			400 => "0000000000011001000101",
			401 => "0001101101111100100000",
			402 => "0000110100011000010100",
			403 => "0010100110011100000100",
			404 => "0000000000011010001001",
			405 => "0000010000011000001100",
			406 => "0001010100011000001000",
			407 => "0011111010011100000100",
			408 => "0000000000011010001001",
			409 => "0000000000011010001001",
			410 => "0000000000011010001001",
			411 => "0000000000011010001001",
			412 => "0001001111101000000100",
			413 => "0000000000011010001001",
			414 => "0001010111001000000100",
			415 => "0000000000011010001001",
			416 => "0000000000011010001001",
			417 => "0000000000011010001001",
			418 => "0001101101111100100000",
			419 => "0000110100011000010100",
			420 => "0000010000011000010000",
			421 => "0001010100011000001100",
			422 => "0000100011001000001000",
			423 => "0010100110011100000100",
			424 => "0000000000011011001101",
			425 => "0000000000011011001101",
			426 => "0000000000011011001101",
			427 => "0000000000011011001101",
			428 => "0000000000011011001101",
			429 => "0001001111101000000100",
			430 => "0000000000011011001101",
			431 => "0001010111001000000100",
			432 => "0000000000011011001101",
			433 => "0000000000011011001101",
			434 => "0000000000011011001101",
			435 => "0011100001010100011000",
			436 => "0001101101111100010000",
			437 => "0000100011001000001100",
			438 => "0001101110010100000100",
			439 => "0000000000011100101001",
			440 => "0010001011000100000100",
			441 => "0000001000011100101001",
			442 => "0000000000011100101001",
			443 => "0000000000011100101001",
			444 => "0001101101111100000100",
			445 => "0000000000011100101001",
			446 => "0000000000011100101001",
			447 => "0001000011011000000100",
			448 => "1111111000011100101001",
			449 => "0001101101111100010000",
			450 => "0011101100001000001100",
			451 => "0000101100100100001000",
			452 => "0001001011100100000100",
			453 => "0000000000011100101001",
			454 => "0000001000011100101001",
			455 => "1111111000011100101001",
			456 => "0000001000011100101001",
			457 => "1111111000011100101001",
			458 => "0000010000011000010100",
			459 => "0001011010111000010000",
			460 => "0001101101111100001100",
			461 => "0001101110010100000100",
			462 => "0000000000011110000101",
			463 => "0000100011001000000100",
			464 => "0000001000011110000101",
			465 => "0000000000011110000101",
			466 => "0000000000011110000101",
			467 => "1111111000011110000101",
			468 => "0010000110011000001000",
			469 => "0001001000100000000100",
			470 => "1111111000011110000101",
			471 => "0000001000011110000101",
			472 => "0001000011011000000100",
			473 => "1111111000011110000101",
			474 => "0001000001101100001100",
			475 => "0011011011011100000100",
			476 => "0000000000011110000101",
			477 => "0001010001011000000100",
			478 => "0000000000011110000101",
			479 => "0000000000011110000101",
			480 => "1111111000011110000101",
			481 => "0001000011011000001100",
			482 => "0010000110011000001000",
			483 => "0000001011010100000100",
			484 => "1111111000011111010001",
			485 => "0000001000011111010001",
			486 => "1111111000011111010001",
			487 => "0001101101111100011000",
			488 => "0001111110001100010100",
			489 => "0001101110010100000100",
			490 => "0000000000011111010001",
			491 => "0000010000011000001000",
			492 => "0000100011001000000100",
			493 => "0000001000011111010001",
			494 => "0000000000011111010001",
			495 => "0000010110000000000100",
			496 => "0000000000011111010001",
			497 => "0000000000011111010001",
			498 => "0000000000011111010001",
			499 => "1111111000011111010001",
			500 => "0000110111000000010000",
			501 => "0001101101111100001100",
			502 => "0011110001111100001000",
			503 => "0010000000101000000100",
			504 => "0000001000100000110101",
			505 => "0000001000100000110101",
			506 => "0000000000100000110101",
			507 => "1111111000100000110101",
			508 => "0011111101010100010000",
			509 => "0001011010111100001100",
			510 => "0000011100100000001000",
			511 => "0001010011011100000100",
			512 => "0000001000100000110101",
			513 => "0000010000100000110101",
			514 => "1111111000100000110101",
			515 => "1111111000100000110101",
			516 => "0001000011011000000100",
			517 => "1111111000100000110101",
			518 => "0001101101111100001100",
			519 => "0001100001111000000100",
			520 => "1111111000100000110101",
			521 => "0001001111011000000100",
			522 => "0000101000100000110101",
			523 => "1111111000100000110101",
			524 => "1111111000100000110101",
			525 => "0001000011011000001100",
			526 => "0010000110011000001000",
			527 => "0001001111100100000100",
			528 => "0000000000100010001001",
			529 => "0000001000100010001001",
			530 => "1111111000100010001001",
			531 => "0001101101111100011100",
			532 => "0001111110001100011000",
			533 => "0000010000011000001100",
			534 => "0001100111101000000100",
			535 => "0000000000100010001001",
			536 => "0000100011001000000100",
			537 => "0000001000100010001001",
			538 => "0000000000100010001001",
			539 => "0010001111001000001000",
			540 => "0001100101011100000100",
			541 => "0000000000100010001001",
			542 => "0000001000100010001001",
			543 => "0000000000100010001001",
			544 => "0000000000100010001001",
			545 => "0000000000100010001001",
			546 => "0000110111000000001100",
			547 => "0001101101111100001000",
			548 => "0011111010111000000100",
			549 => "0000001000100011111101",
			550 => "0000000000100011111101",
			551 => "1111111000100011111101",
			552 => "0011111010111000010100",
			553 => "0001011010111100010000",
			554 => "0001001011100100000100",
			555 => "1111111000100011111101",
			556 => "0001110100010100001000",
			557 => "0001011000111000000100",
			558 => "0000000000100011111101",
			559 => "0000001000100011111101",
			560 => "0000010000100011111101",
			561 => "1111111000100011111101",
			562 => "0001000011011000001100",
			563 => "0001101110010100001000",
			564 => "0001101011111100000100",
			565 => "1111111000100011111101",
			566 => "0000001000100011111101",
			567 => "1111111000100011111101",
			568 => "0001101101111100001100",
			569 => "0001011100101000000100",
			570 => "1111111000100011111101",
			571 => "0010110111001000000100",
			572 => "0000011000100011111101",
			573 => "1111111000100011111101",
			574 => "1111111000100011111101",
			575 => "0000111000101100010100",
			576 => "0001101101111100010000",
			577 => "0001101110010100000100",
			578 => "1111111000100110000001",
			579 => "0000101110010000001000",
			580 => "0000000101001000000100",
			581 => "0000001000100110000001",
			582 => "0000000000100110000001",
			583 => "0000011000100110000001",
			584 => "1111111000100110000001",
			585 => "0000010000011000100000",
			586 => "0000100111100000001100",
			587 => "0000110011111100001000",
			588 => "0001101101111100000100",
			589 => "0000001000100110000001",
			590 => "0000000000100110000001",
			591 => "0000010000100110000001",
			592 => "0010011110100000001100",
			593 => "0000100101001000001000",
			594 => "0000100101001000000100",
			595 => "0000000000100110000001",
			596 => "0000000000100110000001",
			597 => "1111111000100110000001",
			598 => "0011001010000000000100",
			599 => "0000000000100110000001",
			600 => "0000001000100110000001",
			601 => "0001001101110100000100",
			602 => "1111111000100110000001",
			603 => "0001101101111100001000",
			604 => "0001100111101000000100",
			605 => "0000000000100110000001",
			606 => "0000001000100110000001",
			607 => "1111111000100110000001",
			608 => "0001000011011000010000",
			609 => "0001101110010100001100",
			610 => "0000101110101000000100",
			611 => "0000000000100111100101",
			612 => "0000110001111100000100",
			613 => "0000000000100111100101",
			614 => "0000000000100111100101",
			615 => "1111111000100111100101",
			616 => "0001101101111100100000",
			617 => "0001111110001100011100",
			618 => "0001000000101100001100",
			619 => "0010001001101000001000",
			620 => "0010101000100100000100",
			621 => "0000000000100111100101",
			622 => "0000000000100111100101",
			623 => "0000000000100111100101",
			624 => "0001101110010100000100",
			625 => "0000000000100111100101",
			626 => "0000101110110100001000",
			627 => "0010001011000100000100",
			628 => "0000001000100111100101",
			629 => "0000000000100111100101",
			630 => "0000000000100111100101",
			631 => "0000000000100111100101",
			632 => "0000000000100111100101",
			633 => "0000110111000000001100",
			634 => "0001101101111100001000",
			635 => "0001100111101000000100",
			636 => "0000000000101001100001",
			637 => "0000001000101001100001",
			638 => "0000000000101001100001",
			639 => "0001000011011000001100",
			640 => "0010000110011000001000",
			641 => "0000001001101000000100",
			642 => "1111111000101001100001",
			643 => "0000011000101001100001",
			644 => "1111111000101001100001",
			645 => "0000101110000100011000",
			646 => "0001101101111100010100",
			647 => "0011000000101000001100",
			648 => "0000010000011000001000",
			649 => "0001100111101000000100",
			650 => "0000000000101001100001",
			651 => "0000001000101001100001",
			652 => "1111111000101001100001",
			653 => "0000011110011100000100",
			654 => "0000000000101001100001",
			655 => "0000001000101001100001",
			656 => "0000000000101001100001",
			657 => "0001101101111100001100",
			658 => "0001100001111000000100",
			659 => "1111111000101001100001",
			660 => "0001001111110100000100",
			661 => "0000001000101001100001",
			662 => "0000000000101001100001",
			663 => "1111111000101001100001",
			664 => "0011100001110000010100",
			665 => "0001101101111100010000",
			666 => "0011111010111000001100",
			667 => "0000000111100000001000",
			668 => "0001000000000100000100",
			669 => "0000000000101011101101",
			670 => "0000001000101011101101",
			671 => "0000000000101011101101",
			672 => "0000000000101011101101",
			673 => "1111111000101011101101",
			674 => "0001000011011000001100",
			675 => "0001101110010100001000",
			676 => "0001101011111100000100",
			677 => "1111111000101011101101",
			678 => "0000000000101011101101",
			679 => "1111111000101011101101",
			680 => "0010001111001000001100",
			681 => "0000110100011000000100",
			682 => "0000000000101011101101",
			683 => "0011001100110000000100",
			684 => "0000001000101011101101",
			685 => "0000000000101011101101",
			686 => "0000101110101000001100",
			687 => "0000011100100000001000",
			688 => "0000000101001000000100",
			689 => "0000001000101011101101",
			690 => "0000000000101011101101",
			691 => "0000000000101011101101",
			692 => "0001101101111100001100",
			693 => "0001101101111100000100",
			694 => "1111111000101011101101",
			695 => "0001010001101000000100",
			696 => "0000000000101011101101",
			697 => "0000000000101011101101",
			698 => "1111111000101011101101",
			699 => "0000111000101100010100",
			700 => "0001101101111100010000",
			701 => "0001101110010100000100",
			702 => "1111111000101110000011",
			703 => "0000000101001000001000",
			704 => "0000101110010000000100",
			705 => "0000001000101110000011",
			706 => "0000000000101110000011",
			707 => "0000000000101110000011",
			708 => "1111111000101110000011",
			709 => "0011111010111000010000",
			710 => "0011011100101100001100",
			711 => "0000011100100000001000",
			712 => "0001011001110000000100",
			713 => "0000000000101110000011",
			714 => "0000001000101110000011",
			715 => "1111111000101110000011",
			716 => "1111111000101110000011",
			717 => "0001000011011000001100",
			718 => "0001101110010100001000",
			719 => "0001101011111100000100",
			720 => "1111111000101110000011",
			721 => "0000001000101110000011",
			722 => "1111111000101110000011",
			723 => "0000100111100000001000",
			724 => "0001101101111100000100",
			725 => "0000001000101110000011",
			726 => "0000000000101110000011",
			727 => "0000101110110100010000",
			728 => "0000101110110100001000",
			729 => "0001001010010000000100",
			730 => "1111111000101110000011",
			731 => "0000000000101110000011",
			732 => "0001000001001100000100",
			733 => "0000010000101110000011",
			734 => "1111111000101110000011",
			735 => "1111111000101110000011",
			736 => "0000000000101110000101",
			737 => "0000000000101110001001",
			738 => "0000000000101110001101",
			739 => "0000000000101110010001",
			740 => "0000000000101110010101",
			741 => "0000000000101110011001",
			742 => "0000000000101110011101",
			743 => "0000000000101110100001",
			744 => "0000000000101110100101",
			745 => "0000000000101110101001",
			746 => "0000000000101110101101",
			747 => "0000000000101110110001",
			748 => "0000000000101110110101",
			749 => "0000000000101110111001",
			750 => "0000000000101110111101",
			751 => "0000000000101111000001",
			752 => "0000000000101111000101",
			753 => "0000000000101111001001",
			754 => "0000000000101111001101",
			755 => "0000000000101111010001",
			756 => "0000000000101111010101",
			757 => "0000000000101111011001",
			758 => "0000000000101111011101",
			759 => "0000000000101111100001",
			760 => "0000000000101111100101",
			761 => "0000000000101111101001",
			762 => "0000000000101111101101",
			763 => "0000000000101111110001",
			764 => "0000000000101111110101",
			765 => "0001000011011000000100",
			766 => "0000000000110000000001",
			767 => "0000000000110000000001",
			768 => "0000100111100000000100",
			769 => "0000000000110000001101",
			770 => "0000000000110000001101",
			771 => "0000111010101100000100",
			772 => "0000000000110000011001",
			773 => "0000000000110000011001",
			774 => "0000101100100100000100",
			775 => "0000000000110000100101",
			776 => "0000000000110000100101",
			777 => "0001101101111100001000",
			778 => "0001100111101000000100",
			779 => "0000000000110000111001",
			780 => "0000000000110000111001",
			781 => "0000000000110000111001",
			782 => "0001101101111100001000",
			783 => "0001101011111100000100",
			784 => "0000000000110001001101",
			785 => "0000000000110001001101",
			786 => "0000000000110001001101",
			787 => "0001101101111100001000",
			788 => "0001101011111100000100",
			789 => "0000000000110001100001",
			790 => "0000000000110001100001",
			791 => "0000000000110001100001",
			792 => "0001001011100100001000",
			793 => "0000110100011000000100",
			794 => "0000000000110001110101",
			795 => "0000000000110001110101",
			796 => "0000000000110001110101",
			797 => "0001101101111100001000",
			798 => "0001101011111100000100",
			799 => "0000000000110010001001",
			800 => "0000000000110010001001",
			801 => "0000000000110010001001",
			802 => "0001101101111100001000",
			803 => "0001101011111100000100",
			804 => "0000000000110010011101",
			805 => "0000000000110010011101",
			806 => "0000000000110010011101",
			807 => "0000101100100100000100",
			808 => "0000000000110010110001",
			809 => "0000110111000000000100",
			810 => "0000000000110010110001",
			811 => "0000000000110010110001",
			812 => "0001101101111100001000",
			813 => "0001101011111100000100",
			814 => "0000000000110011000101",
			815 => "0000000000110011000101",
			816 => "0000000000110011000101",
			817 => "0001101101111100001000",
			818 => "0001101011111100000100",
			819 => "0000000000110011011001",
			820 => "0000000000110011011001",
			821 => "0000000000110011011001",
			822 => "0001101101111100001000",
			823 => "0001101011111100000100",
			824 => "0000000000110011101101",
			825 => "0000000000110011101101",
			826 => "0000000000110011101101",
			827 => "0001101101111100001000",
			828 => "0001101011111100000100",
			829 => "0000000000110100000001",
			830 => "0000000000110100000001",
			831 => "0000000000110100000001",
			832 => "0001000101100000001100",
			833 => "0011110011011100000100",
			834 => "0000000000110100011101",
			835 => "0001010110100100000100",
			836 => "0000000000110100011101",
			837 => "0000000000110100011101",
			838 => "0000000000110100011101",
			839 => "0001101101111100001100",
			840 => "0001101011111100000100",
			841 => "0000000000110100111001",
			842 => "0001101101111100000100",
			843 => "0000000000110100111001",
			844 => "0000000000110100111001",
			845 => "0000000000110100111001",
			846 => "0000100111100000001100",
			847 => "0001101101111100001000",
			848 => "0001101011111100000100",
			849 => "0000000000110101011101",
			850 => "0000000000110101011101",
			851 => "0000000000110101011101",
			852 => "0000101000001100000100",
			853 => "0000000000110101011101",
			854 => "0000000000110101011101",
			855 => "0001101101111100010000",
			856 => "0000110100011000000100",
			857 => "0000000000110110000001",
			858 => "0000001011010100000100",
			859 => "0000000000110110000001",
			860 => "0011011011000000000100",
			861 => "0000000000110110000001",
			862 => "0000000000110110000001",
			863 => "0000000000110110000001",
			864 => "0001000011011000000100",
			865 => "0000000000110110100101",
			866 => "0011000011011100001100",
			867 => "0000101110110100001000",
			868 => "0010000100010100000100",
			869 => "0000000000110110100101",
			870 => "0000000000110110100101",
			871 => "0000000000110110100101",
			872 => "0000000000110110100101",
			873 => "0000100111100000010000",
			874 => "0000011100110100001100",
			875 => "0001001111101000000100",
			876 => "0000000000110111010001",
			877 => "0001001101110000000100",
			878 => "0000000000110111010001",
			879 => "0000000000110111010001",
			880 => "0000000000110111010001",
			881 => "0000110111000000000100",
			882 => "0000000000110111010001",
			883 => "0000000000110111010001",
			884 => "0001101101111100010000",
			885 => "0001101011111100000100",
			886 => "0000000000110111111101",
			887 => "0000001011010100000100",
			888 => "0000000000110111111101",
			889 => "0010000100010100000100",
			890 => "0000000000110111111101",
			891 => "0000000000110111111101",
			892 => "0000110111000100000100",
			893 => "0000000000110111111101",
			894 => "0000000000110111111101",
			895 => "0000110111000000001100",
			896 => "0001101101111100001000",
			897 => "0011110111001000000100",
			898 => "0000010000111000110001",
			899 => "1111111000111000110001",
			900 => "1111111000111000110001",
			901 => "0011110001111100001100",
			902 => "0001011010111100001000",
			903 => "0000011100100000000100",
			904 => "0000010000111000110001",
			905 => "1111111000111000110001",
			906 => "1111111000111000110001",
			907 => "1111111000111000110001",
			908 => "0000110111000000010000",
			909 => "0001101101111100001100",
			910 => "0011110111001000001000",
			911 => "0010100001110100000100",
			912 => "0000001000111001101101",
			913 => "0000000000111001101101",
			914 => "1111111000111001101101",
			915 => "1111111000111001101101",
			916 => "0011110001111100001100",
			917 => "0010110000101000001000",
			918 => "0000011100100000000100",
			919 => "0000001000111001101101",
			920 => "1111111000111001101101",
			921 => "1111111000111001101101",
			922 => "1111111000111001101101",
			923 => "0000100111100000010100",
			924 => "0000011100110100010000",
			925 => "0001101101111100001100",
			926 => "0001101011111100000100",
			927 => "0000000000111010100001",
			928 => "0001001101110000000100",
			929 => "0000000000111010100001",
			930 => "0000000000111010100001",
			931 => "0000000000111010100001",
			932 => "0000000000111010100001",
			933 => "0000110111000000000100",
			934 => "0000000000111010100001",
			935 => "0000000000111010100001",
			936 => "0001000011011000000100",
			937 => "1111111000111011001101",
			938 => "0001110110000100010000",
			939 => "0001101101111100001100",
			940 => "0001100111101000000100",
			941 => "0000000000111011001101",
			942 => "0010001011000100000100",
			943 => "0000000000111011001101",
			944 => "0000000000111011001101",
			945 => "0000000000111011001101",
			946 => "0000000000111011001101",
			947 => "0000110111000000010000",
			948 => "0001101101111100001100",
			949 => "0011110111001000001000",
			950 => "0011011101100000000100",
			951 => "0000001000111100010001",
			952 => "0000000000111100010001",
			953 => "1111111000111100010001",
			954 => "1111111000111100010001",
			955 => "0011110001111100001100",
			956 => "0010110000101000001000",
			957 => "0000011100100000000100",
			958 => "0000001000111100010001",
			959 => "1111111000111100010001",
			960 => "1111111000111100010001",
			961 => "0001101101111100000100",
			962 => "1111111000111100010001",
			963 => "1111111000111100010001",
			964 => "0001000011011000001000",
			965 => "0001101110010100000100",
			966 => "0000000000111101010101",
			967 => "1111111000111101010101",
			968 => "0000100111100000010000",
			969 => "0001101101111100001100",
			970 => "0001001101110000001000",
			971 => "0001100111101000000100",
			972 => "0000000000111101010101",
			973 => "0000000000111101010101",
			974 => "0000000000111101010101",
			975 => "0000000000111101010101",
			976 => "0010000110001000000100",
			977 => "0000000000111101010101",
			978 => "0000110111000000000100",
			979 => "0000000000111101010101",
			980 => "0000000000111101010101",
			981 => "0000111010101100001100",
			982 => "0010100010101000001000",
			983 => "0010010000011000000100",
			984 => "0000011000111110100001",
			985 => "0000010000111110100001",
			986 => "1111111000111110100001",
			987 => "0000111000101100001100",
			988 => "0000001001001000001000",
			989 => "0001011000111000000100",
			990 => "1111111000111110100001",
			991 => "0000100000111110100001",
			992 => "1111111000111110100001",
			993 => "0011110001111100001100",
			994 => "0010110000101000001000",
			995 => "0010010110000000000100",
			996 => "0000011000111110100001",
			997 => "1111111000111110100001",
			998 => "1111111000111110100001",
			999 => "1111111000111110100001",
			1000 => "0000010000011000010100",
			1001 => "0001011010111000010000",
			1002 => "0001101101111100001100",
			1003 => "0001100111101000000100",
			1004 => "0000000000111111101101",
			1005 => "0000100011001000000100",
			1006 => "0000001000111111101101",
			1007 => "0000000000111111101101",
			1008 => "0000000000111111101101",
			1009 => "0000000000111111101101",
			1010 => "0010000110011000001000",
			1011 => "0000100111010100000100",
			1012 => "1111111000111111101101",
			1013 => "0000001000111111101101",
			1014 => "0011011001110100000100",
			1015 => "1111111000111111101101",
			1016 => "0011011001110100000100",
			1017 => "0000000000111111101101",
			1018 => "1111111000111111101101",
			1019 => "0001101101111100011100",
			1020 => "0000110100011000010000",
			1021 => "0000001001110000000100",
			1022 => "1111111001000000101001",
			1023 => "0000100111100000001000",
			1024 => "0000001100100100000100",
			1025 => "0000000001000000101001",
			1026 => "0000000001000000101001",
			1027 => "0000000001000000101001",
			1028 => "0000001011010100000100",
			1029 => "0000000001000000101001",
			1030 => "0011011001001000000100",
			1031 => "0000000001000000101001",
			1032 => "0000001001000000101001",
			1033 => "1111111001000000101001",
			1034 => "0001101101111100011100",
			1035 => "0011011010111100010000",
			1036 => "0010010110000000001100",
			1037 => "0011111010111000001000",
			1038 => "0001101110010100000100",
			1039 => "0000000001000001100101",
			1040 => "0000000001000001100101",
			1041 => "0000000001000001100101",
			1042 => "0000000001000001100101",
			1043 => "0010011110100000000100",
			1044 => "0000000001000001100101",
			1045 => "0001001111101000000100",
			1046 => "0000000001000001100101",
			1047 => "0000001001000001100101",
			1048 => "0000000001000001100101",
			1049 => "0001101101111100011100",
			1050 => "0011011010111100001100",
			1051 => "0010010110000000001000",
			1052 => "0010100110011100000100",
			1053 => "0000000001000010100001",
			1054 => "0000000001000010100001",
			1055 => "0000000001000010100001",
			1056 => "0001001011110000000100",
			1057 => "0000000001000010100001",
			1058 => "0010011110100000000100",
			1059 => "0000000001000010100001",
			1060 => "0001100001111000000100",
			1061 => "0000000001000010100001",
			1062 => "0000000001000010100001",
			1063 => "0000000001000010100001",
			1064 => "0010011100110100011100",
			1065 => "0000110001110100001000",
			1066 => "0011111101111000000100",
			1067 => "0000001001000011110101",
			1068 => "0000000001000011110101",
			1069 => "0001010011011100001000",
			1070 => "0010010000011000000100",
			1071 => "0000000001000011110101",
			1072 => "0000000001000011110101",
			1073 => "0001011010111000001000",
			1074 => "0010100110011100000100",
			1075 => "0000000001000011110101",
			1076 => "0000001001000011110101",
			1077 => "0000000001000011110101",
			1078 => "0011011010011100000100",
			1079 => "1111111001000011110101",
			1080 => "0001101101111100001000",
			1081 => "0000001001101000000100",
			1082 => "0000000001000011110101",
			1083 => "0000001001000011110101",
			1084 => "1111111001000011110101",
			1085 => "0011011001110100001100",
			1086 => "0001000100111000001000",
			1087 => "0010010000011000000100",
			1088 => "0000000001000100111001",
			1089 => "0000000001000100111001",
			1090 => "0000000001000100111001",
			1091 => "0011000100001000010100",
			1092 => "0010100001010000010000",
			1093 => "0001001111101000000100",
			1094 => "0000000001000100111001",
			1095 => "0000011101101000001000",
			1096 => "0011000100000000000100",
			1097 => "0000000001000100111001",
			1098 => "0000000001000100111001",
			1099 => "0000000001000100111001",
			1100 => "0000000001000100111001",
			1101 => "0000000001000100111001",
			1102 => "0001000011011000000100",
			1103 => "1111111001000101110101",
			1104 => "0011000011011100011000",
			1105 => "0011011010111100010000",
			1106 => "0001000101100000001000",
			1107 => "0000011100100000000100",
			1108 => "0000000001000101110101",
			1109 => "1111111001000101110101",
			1110 => "0011111010111000000100",
			1111 => "0000001001000101110101",
			1112 => "0000000001000101110101",
			1113 => "0000101110110100000100",
			1114 => "0000001001000101110101",
			1115 => "0000000001000101110101",
			1116 => "0000000001000101110101",
			1117 => "0001101101111100100000",
			1118 => "0001011100101000010000",
			1119 => "0011111010111000001100",
			1120 => "0010100110011100000100",
			1121 => "0000000001000110111001",
			1122 => "0001100111101000000100",
			1123 => "0000000001000110111001",
			1124 => "0000000001000110111001",
			1125 => "1111111001000110111001",
			1126 => "0001001111101000000100",
			1127 => "0000000001000110111001",
			1128 => "0000010000011000000100",
			1129 => "0000000001000110111001",
			1130 => "0010111000111000000100",
			1131 => "0000000001000110111001",
			1132 => "0000001001000110111001",
			1133 => "1111111001000110111001",
			1134 => "0011100101000100010000",
			1135 => "0011111010111000001100",
			1136 => "0001000101001100000100",
			1137 => "0000000001001000001101",
			1138 => "0010100010101000000100",
			1139 => "0000000001001000001101",
			1140 => "0000000001001000001101",
			1141 => "0000000001001000001101",
			1142 => "0011011010011100001000",
			1143 => "0000011100100000000100",
			1144 => "0000000001001000001101",
			1145 => "1111111001001000001101",
			1146 => "0011000100001000010000",
			1147 => "0010101001000100001100",
			1148 => "0001001011110000000100",
			1149 => "0000000001001000001101",
			1150 => "0000011101011100000100",
			1151 => "0000000001001000001101",
			1152 => "0000000001001000001101",
			1153 => "0000000001001000001101",
			1154 => "0000000001001000001101",
			1155 => "0001101101111100100000",
			1156 => "0000110100011000010100",
			1157 => "0010100110011100000100",
			1158 => "0000000001001001010001",
			1159 => "0000100111100000001100",
			1160 => "0001001011100100000100",
			1161 => "0000000001001001010001",
			1162 => "0000000001001000000100",
			1163 => "0000000001001001010001",
			1164 => "0000000001001001010001",
			1165 => "0000000001001001010001",
			1166 => "0001001111101000000100",
			1167 => "0000000001001001010001",
			1168 => "0001010111001000000100",
			1169 => "0000000001001001010001",
			1170 => "0000000001001001010001",
			1171 => "0000000001001001010001",
			1172 => "0000110111000000001100",
			1173 => "0010000100000000001000",
			1174 => "0001100111101000000100",
			1175 => "0000000001001010101101",
			1176 => "0000001001001010101101",
			1177 => "1111111001001010101101",
			1178 => "0011111101010100010000",
			1179 => "0011001100001000001100",
			1180 => "0001001101000000000100",
			1181 => "1111111001001010101101",
			1182 => "0001100001111000000100",
			1183 => "0000001001001010101101",
			1184 => "0000010001001010101101",
			1185 => "1111111001001010101101",
			1186 => "0001000011011000000100",
			1187 => "1111111001001010101101",
			1188 => "0001101101111100001100",
			1189 => "0001100001111000000100",
			1190 => "1111111001001010101101",
			1191 => "0001001111011000000100",
			1192 => "0000011001001010101101",
			1193 => "1111111001001010101101",
			1194 => "1111111001001010101101",
			1195 => "0011100001010100011000",
			1196 => "0001101101111100010000",
			1197 => "0011111010111000001100",
			1198 => "0001000101001100000100",
			1199 => "0000000001001100001001",
			1200 => "0010001011000100000100",
			1201 => "0000001001001100001001",
			1202 => "0000000001001100001001",
			1203 => "0000000001001100001001",
			1204 => "0001101101111100000100",
			1205 => "0000000001001100001001",
			1206 => "0000000001001100001001",
			1207 => "0001000011011000000100",
			1208 => "1111111001001100001001",
			1209 => "0001101101111100010000",
			1210 => "0000111100101100001100",
			1211 => "0011111101010100001000",
			1212 => "0001001101100100000100",
			1213 => "0000000001001100001001",
			1214 => "0000000001001100001001",
			1215 => "1111111001001100001001",
			1216 => "0000001001001100001001",
			1217 => "1111111001001100001001",
			1218 => "0011011001110100011000",
			1219 => "0001000100111000001000",
			1220 => "0000011100100000000100",
			1221 => "0000000001001101100101",
			1222 => "1111111001001101100101",
			1223 => "0000100011001000001100",
			1224 => "0001000101100000000100",
			1225 => "0000000001001101100101",
			1226 => "0001011110110000000100",
			1227 => "0000000001001101100101",
			1228 => "0000000001001101100101",
			1229 => "0000000001001101100101",
			1230 => "0011000100001000010100",
			1231 => "0010100001010000010000",
			1232 => "0001001111101000000100",
			1233 => "0000000001001101100101",
			1234 => "0000011101101000001000",
			1235 => "0011000100000000000100",
			1236 => "0000000001001101100101",
			1237 => "0000001001001101100101",
			1238 => "0000000001001101100101",
			1239 => "0000000001001101100101",
			1240 => "0000000001001101100101",
			1241 => "0001000011011000001100",
			1242 => "0010000110011000001000",
			1243 => "0000001001101000000100",
			1244 => "0000000001001110110001",
			1245 => "0000001001001110110001",
			1246 => "1111111001001110110001",
			1247 => "0001101101111100011000",
			1248 => "0001111110001100010100",
			1249 => "0001101110010100000100",
			1250 => "0000000001001110110001",
			1251 => "0000010000011000001000",
			1252 => "0000100011001000000100",
			1253 => "0000001001001110110001",
			1254 => "0000000001001110110001",
			1255 => "0000010110000000000100",
			1256 => "0000000001001110110001",
			1257 => "0000000001001110110001",
			1258 => "0000000001001110110001",
			1259 => "1111111001001110110001",
			1260 => "0000010000011000010100",
			1261 => "0001011010111000010000",
			1262 => "0001001011100100000100",
			1263 => "0000000001010000010101",
			1264 => "0010100110011100000100",
			1265 => "0000000001010000010101",
			1266 => "0011111010011100000100",
			1267 => "0000001001010000010101",
			1268 => "0000000001010000010101",
			1269 => "0000000001010000010101",
			1270 => "0010000110011000001100",
			1271 => "0011110111010100000100",
			1272 => "1111111001010000010101",
			1273 => "0011011110010000000100",
			1274 => "0000001001010000010101",
			1275 => "0000000001010000010101",
			1276 => "0001001101110100000100",
			1277 => "1111111001010000010101",
			1278 => "0001000000100000000100",
			1279 => "0000000001010000010101",
			1280 => "0001000001100100001000",
			1281 => "0001000000101100000100",
			1282 => "0000000001010000010101",
			1283 => "0000000001010000010101",
			1284 => "1111111001010000010101",
			1285 => "0000110111000000001100",
			1286 => "0001101101111100001000",
			1287 => "0001100111101000000100",
			1288 => "0000000001010010000001",
			1289 => "0000001001010010000001",
			1290 => "1111111001010010000001",
			1291 => "0001000011011000001100",
			1292 => "0010000110011000001000",
			1293 => "0001001000100000000100",
			1294 => "1111111001010010000001",
			1295 => "0000100001010010000001",
			1296 => "1111111001010010000001",
			1297 => "0000101110000100010000",
			1298 => "0010111100001000001000",
			1299 => "0011111010111100000100",
			1300 => "0000001001010010000001",
			1301 => "1111111001010010000001",
			1302 => "0010011100100000000100",
			1303 => "0000000001010010000001",
			1304 => "0000001001010010000001",
			1305 => "0001101101111100001100",
			1306 => "0001100001111000000100",
			1307 => "1111111001010010000001",
			1308 => "0001001111110100000100",
			1309 => "0000001001010010000001",
			1310 => "0000000001010010000001",
			1311 => "1111111001010010000001",
			1312 => "0000110111000000010000",
			1313 => "0001101101111100001000",
			1314 => "0001100111101000000100",
			1315 => "0000000001010011110101",
			1316 => "0000001001010011110101",
			1317 => "0000111010101100000100",
			1318 => "0000000001010011110101",
			1319 => "0000000001010011110101",
			1320 => "0001000011011000001100",
			1321 => "0000001011010100001000",
			1322 => "0001001101101100000100",
			1323 => "1111111001010011110101",
			1324 => "0000010001010011110101",
			1325 => "1111111001010011110101",
			1326 => "0000000011010000001000",
			1327 => "0011001100110000000100",
			1328 => "0000010001010011110101",
			1329 => "0000000001010011110101",
			1330 => "0001101101111100010100",
			1331 => "0001100001111000001000",
			1332 => "0011111010111100000100",
			1333 => "0000000001010011110101",
			1334 => "1111111001010011110101",
			1335 => "0001111101111000001000",
			1336 => "0001111011000100000100",
			1337 => "0000000001010011110101",
			1338 => "0000001001010011110101",
			1339 => "0000000001010011110101",
			1340 => "1111111001010011110101",
			1341 => "0000110111000000010100",
			1342 => "0001101101111100001100",
			1343 => "0001100111101000000100",
			1344 => "0000000001010101101001",
			1345 => "0010100111000100000100",
			1346 => "0000001001010101101001",
			1347 => "0000000001010101101001",
			1348 => "0000111010101100000100",
			1349 => "0000000001010101101001",
			1350 => "0000000001010101101001",
			1351 => "0001101101111100100100",
			1352 => "0011011010011100011000",
			1353 => "0010100001010100001000",
			1354 => "0011110110000100000100",
			1355 => "0000000001010101101001",
			1356 => "1111111001010101101001",
			1357 => "0000001110110000001100",
			1358 => "0011111110110000000100",
			1359 => "0000001001010101101001",
			1360 => "0011111000011000000100",
			1361 => "0000000001010101101001",
			1362 => "0000000001010101101001",
			1363 => "0000000001010101101001",
			1364 => "0000001011010100000100",
			1365 => "1111111001010101101001",
			1366 => "0011111011011100000100",
			1367 => "0000000001010101101001",
			1368 => "0000010001010101101001",
			1369 => "1111111001010101101001",
			1370 => "0000111000101100011000",
			1371 => "0001101110010100000100",
			1372 => "1111111001010111100101",
			1373 => "0001101101111100010000",
			1374 => "0001001111111000001100",
			1375 => "0011111110110000001000",
			1376 => "0011010011011100000100",
			1377 => "0000001001010111100101",
			1378 => "0000001001010111100101",
			1379 => "0000000001010111100101",
			1380 => "0000000001010111100101",
			1381 => "1111111001010111100101",
			1382 => "0011111010111000010000",
			1383 => "0011001100001000001100",
			1384 => "0000011100100000001000",
			1385 => "0001100111101000000100",
			1386 => "0000000001010111100101",
			1387 => "0000001001010111100101",
			1388 => "1111111001010111100101",
			1389 => "1111111001010111100101",
			1390 => "0001001101110100000100",
			1391 => "1111111001010111100101",
			1392 => "0001101101111100010000",
			1393 => "0010011110100000000100",
			1394 => "1111111001010111100101",
			1395 => "0011110001101000000100",
			1396 => "1111111001010111100101",
			1397 => "0001101110010100000100",
			1398 => "0000000001010111100101",
			1399 => "0000001001010111100101",
			1400 => "1111111001010111100101",
			1401 => "0000111000101100010100",
			1402 => "0010000100000000010000",
			1403 => "0001000101100000000100",
			1404 => "0000000001011001101001",
			1405 => "0011111010111000001000",
			1406 => "0010111011000100000100",
			1407 => "0000001001011001101001",
			1408 => "0000010001011001101001",
			1409 => "0000000001011001101001",
			1410 => "1111111001011001101001",
			1411 => "0011111010111000010000",
			1412 => "0011001100001000001100",
			1413 => "0000011100100000001000",
			1414 => "0011001010000000000100",
			1415 => "0000000001011001101001",
			1416 => "0000001001011001101001",
			1417 => "1111111001011001101001",
			1418 => "1111111001011001101001",
			1419 => "0001001101110100000100",
			1420 => "1111111001011001101001",
			1421 => "0001000000100000001100",
			1422 => "0010010110101000000100",
			1423 => "0000000001011001101001",
			1424 => "0000010110101000000100",
			1425 => "0000010001011001101001",
			1426 => "0000000001011001101001",
			1427 => "0001000001100100001100",
			1428 => "0010011011101000000100",
			1429 => "1111111001011001101001",
			1430 => "0010011101011000000100",
			1431 => "0000001001011001101001",
			1432 => "0000000001011001101001",
			1433 => "1111111001011001101001",
			1434 => "0011100001010100010100",
			1435 => "0001101101111100010000",
			1436 => "0001101110010100000100",
			1437 => "0000000001011011100101",
			1438 => "0000101100010100001000",
			1439 => "0000000111100000000100",
			1440 => "0000001001011011100101",
			1441 => "0000000001011011100101",
			1442 => "0000000001011011100101",
			1443 => "0000000001011011100101",
			1444 => "0001000011011000001100",
			1445 => "0001101110010100001000",
			1446 => "0001101011111100000100",
			1447 => "1111111001011011100101",
			1448 => "0000000001011011100101",
			1449 => "1111111001011011100101",
			1450 => "0001101101111100011100",
			1451 => "0011101100001000011000",
			1452 => "0001000100111000001100",
			1453 => "0000110011111100001000",
			1454 => "0011101001101000000100",
			1455 => "0000000001011011100101",
			1456 => "0000000001011011100101",
			1457 => "1111111001011011100101",
			1458 => "0001011000000000001000",
			1459 => "0001110111111000000100",
			1460 => "0000000001011011100101",
			1461 => "0000001001011011100101",
			1462 => "0000000001011011100101",
			1463 => "0000001001011011100101",
			1464 => "1111111001011011100101",
			1465 => "0000110111000000010000",
			1466 => "0001101101111100001100",
			1467 => "0011111010111000001000",
			1468 => "0011000100000000000100",
			1469 => "0000001001011101111011",
			1470 => "0000000001011101111011",
			1471 => "0000000001011101111011",
			1472 => "1111111001011101111011",
			1473 => "0011111010111000010100",
			1474 => "0001011010111100010000",
			1475 => "0001001011100100000100",
			1476 => "1111111001011101111011",
			1477 => "0001011000111000000100",
			1478 => "0000000001011101111011",
			1479 => "0011110000001100000100",
			1480 => "0000001001011101111011",
			1481 => "0000010001011101111011",
			1482 => "1111111001011101111011",
			1483 => "0001000011011000001100",
			1484 => "0001101110010100001000",
			1485 => "0001101011111100000100",
			1486 => "1111111001011101111011",
			1487 => "0000001001011101111011",
			1488 => "1111111001011101111011",
			1489 => "0010001111001000001100",
			1490 => "0000011110100000000100",
			1491 => "1111111001011101111011",
			1492 => "0010110111001000000100",
			1493 => "0000010001011101111011",
			1494 => "0000000001011101111011",
			1495 => "0001101101111100001100",
			1496 => "0001011100101000000100",
			1497 => "1111111001011101111011",
			1498 => "0001011010011100000100",
			1499 => "0000001001011101111011",
			1500 => "1111111001011101111011",
			1501 => "1111111001011101111011",
			1502 => "0000000001011101111101",
			1503 => "0000000001011110000001",
			1504 => "0000000001011110000101",
			1505 => "0000000001011110001001",
			1506 => "0000000001011110001101",
			1507 => "0000000001011110010001",
			1508 => "0000000001011110010101",
			1509 => "0000000001011110011001",
			1510 => "0000000001011110011101",
			1511 => "0000000001011110100001",
			1512 => "0000000001011110100101",
			1513 => "0000000001011110101001",
			1514 => "0000000001011110101101",
			1515 => "0000000001011110110001",
			1516 => "0000000001011110110101",
			1517 => "0000000001011110111001",
			1518 => "0000000001011110111101",
			1519 => "0000000001011111000001",
			1520 => "0000000001011111000101",
			1521 => "0000000001011111001001",
			1522 => "0000000001011111001101",
			1523 => "0000000001011111010001",
			1524 => "0000000001011111010101",
			1525 => "0000000001011111011001",
			1526 => "0000000001011111011101",
			1527 => "0000000001011111100001",
			1528 => "0000000001011111100101",
			1529 => "0000000001011111101001",
			1530 => "0000000001011111101101",
			1531 => "0000100111100000000100",
			1532 => "0000000001011111111001",
			1533 => "0000000001011111111001",
			1534 => "0011101010110000000100",
			1535 => "0000000001100000000101",
			1536 => "0000000001100000000101",
			1537 => "0000101100100100000100",
			1538 => "0000000001100000010001",
			1539 => "0000000001100000010001",
			1540 => "0000101100100100000100",
			1541 => "0000000001100000011101",
			1542 => "0000000001100000011101",
			1543 => "0001101101111100001000",
			1544 => "0001100111101000000100",
			1545 => "0000000001100000110001",
			1546 => "0000000001100000110001",
			1547 => "0000000001100000110001",
			1548 => "0000010000011000000100",
			1549 => "0000000001100001000101",
			1550 => "0011011001110100000100",
			1551 => "0000000001100001000101",
			1552 => "0000000001100001000101",
			1553 => "0001101101111100001000",
			1554 => "0001101011111100000100",
			1555 => "0000000001100001011001",
			1556 => "0000000001100001011001",
			1557 => "0000000001100001011001",
			1558 => "0001001011100100001000",
			1559 => "0000110100011000000100",
			1560 => "0000000001100001101101",
			1561 => "0000000001100001101101",
			1562 => "0000000001100001101101",
			1563 => "0001101101111100001000",
			1564 => "0001101011111100000100",
			1565 => "0000000001100010000001",
			1566 => "0000000001100010000001",
			1567 => "0000000001100010000001",
			1568 => "0000101100100100000100",
			1569 => "0000000001100010010101",
			1570 => "0000110111000000000100",
			1571 => "0000000001100010010101",
			1572 => "0000000001100010010101",
			1573 => "0001101101111100001000",
			1574 => "0001101011111100000100",
			1575 => "0000000001100010101001",
			1576 => "0000000001100010101001",
			1577 => "0000000001100010101001",
			1578 => "0001101101111100001000",
			1579 => "0001101011111100000100",
			1580 => "0000000001100010111101",
			1581 => "0000000001100010111101",
			1582 => "0000000001100010111101",
			1583 => "0001101101111100001000",
			1584 => "0001101011111100000100",
			1585 => "0000000001100011010001",
			1586 => "0000000001100011010001",
			1587 => "0000000001100011010001",
			1588 => "0001101101111100001000",
			1589 => "0001101011111100000100",
			1590 => "0000000001100011100101",
			1591 => "0000000001100011100101",
			1592 => "0000000001100011100101",
			1593 => "0000100111100000001000",
			1594 => "0000100000110100000100",
			1595 => "0000000001100100000001",
			1596 => "0000000001100100000001",
			1597 => "0000101000001100000100",
			1598 => "0000000001100100000001",
			1599 => "0000000001100100000001",
			1600 => "0001000101100000001100",
			1601 => "0011110011011100000100",
			1602 => "0000000001100100011101",
			1603 => "0001010110100100000100",
			1604 => "0000000001100100011101",
			1605 => "0000000001100100011101",
			1606 => "0000000001100100011101",
			1607 => "0001101101111100001100",
			1608 => "0001101011111100000100",
			1609 => "0000000001100100111001",
			1610 => "0001101101111100000100",
			1611 => "0000000001100100111001",
			1612 => "0000000001100100111001",
			1613 => "0000000001100100111001",
			1614 => "0000100111100000001100",
			1615 => "0001101011111100000100",
			1616 => "0000000001100101011101",
			1617 => "0001101101111100000100",
			1618 => "0000000001100101011101",
			1619 => "0000000001100101011101",
			1620 => "0000101000001100000100",
			1621 => "0000000001100101011101",
			1622 => "0000000001100101011101",
			1623 => "0001000101100000010000",
			1624 => "0000100111010000000100",
			1625 => "0000000001100110000001",
			1626 => "0010110000001100001000",
			1627 => "0000011110011100000100",
			1628 => "0000000001100110000001",
			1629 => "0000000001100110000001",
			1630 => "0000000001100110000001",
			1631 => "0000000001100110000001",
			1632 => "0001000011011000000100",
			1633 => "0000000001100110100101",
			1634 => "0001110110000100001100",
			1635 => "0001101101111100001000",
			1636 => "0001101110010100000100",
			1637 => "0000000001100110100101",
			1638 => "0000000001100110100101",
			1639 => "0000000001100110100101",
			1640 => "0000000001100110100101",
			1641 => "0001101101111100010000",
			1642 => "0001001111101000000100",
			1643 => "0000000001100111010001",
			1644 => "0001101011111100000100",
			1645 => "0000000001100111010001",
			1646 => "0010000100010100000100",
			1647 => "0000000001100111010001",
			1648 => "0000000001100111010001",
			1649 => "0001001010010000000100",
			1650 => "0000000001100111010001",
			1651 => "0000000001100111010001",
			1652 => "0011011001110100001000",
			1653 => "0000110001110100000100",
			1654 => "0000000001100111111101",
			1655 => "0000000001100111111101",
			1656 => "0001101101111100001100",
			1657 => "0000110100011000000100",
			1658 => "0000000001100111111101",
			1659 => "0001101011111100000100",
			1660 => "0000000001100111111101",
			1661 => "0000000001100111111101",
			1662 => "0000000001100111111101",
			1663 => "0001000011011000001100",
			1664 => "0010000110011000001000",
			1665 => "0001001000100000000100",
			1666 => "1111111001101000110001",
			1667 => "0000001001101000110001",
			1668 => "1111111001101000110001",
			1669 => "0001101101111100001100",
			1670 => "0001111110001100001000",
			1671 => "0001101110010100000100",
			1672 => "0000000001101000110001",
			1673 => "0000001001101000110001",
			1674 => "0000000001101000110001",
			1675 => "1111111001101000110001",
			1676 => "0001000011011000001000",
			1677 => "0001101110010100000100",
			1678 => "0000000001101001100101",
			1679 => "1111111001101001100101",
			1680 => "0001101101111100010000",
			1681 => "0011001100110000001100",
			1682 => "0001100111101000000100",
			1683 => "0000000001101001100101",
			1684 => "0010001011000100000100",
			1685 => "0000000001101001100101",
			1686 => "0000000001101001100101",
			1687 => "0000000001101001100101",
			1688 => "0000000001101001100101",
			1689 => "0001000011011000000100",
			1690 => "1111111001101010010001",
			1691 => "0001101101111100010000",
			1692 => "0001111110001100001100",
			1693 => "0001101110010100000100",
			1694 => "0000000001101010010001",
			1695 => "0000101110110100000100",
			1696 => "0000001001101010010001",
			1697 => "0000000001101010010001",
			1698 => "0000000001101010010001",
			1699 => "0000000001101010010001",
			1700 => "0001000011011000000100",
			1701 => "1111111001101010111101",
			1702 => "0011000011011100010000",
			1703 => "0001101101111100001100",
			1704 => "0001100111101000000100",
			1705 => "0000000001101010111101",
			1706 => "0010001011000100000100",
			1707 => "0000000001101010111101",
			1708 => "0000000001101010111101",
			1709 => "0000000001101010111101",
			1710 => "0000000001101010111101",
			1711 => "0000111010101100001000",
			1712 => "0001101101111100000100",
			1713 => "1110110001101011111001",
			1714 => "1101010001101011111001",
			1715 => "0000110111000000001000",
			1716 => "0000000011100000000100",
			1717 => "1110011001101011111001",
			1718 => "1101001001101011111001",
			1719 => "0011110001111100001100",
			1720 => "0010110000101000001000",
			1721 => "0000011100100000000100",
			1722 => "1110110001101011111001",
			1723 => "1101010001101011111001",
			1724 => "1101001001101011111001",
			1725 => "1101001001101011111001",
			1726 => "0001000011011000001000",
			1727 => "0001101110010100000100",
			1728 => "0000000001101100111101",
			1729 => "1111111001101100111101",
			1730 => "0000100111100000010000",
			1731 => "0001101101111100001100",
			1732 => "0000000001001000001000",
			1733 => "0001100111101000000100",
			1734 => "0000000001101100111101",
			1735 => "0000000001101100111101",
			1736 => "0000000001101100111101",
			1737 => "0000000001101100111101",
			1738 => "0010000110001000000100",
			1739 => "0000000001101100111101",
			1740 => "0000110111000000000100",
			1741 => "0000000001101100111101",
			1742 => "0000000001101100111101",
			1743 => "0000010000011000010100",
			1744 => "0001011010111000010000",
			1745 => "0001101101111100001100",
			1746 => "0001101110010100000100",
			1747 => "0000000001101110001001",
			1748 => "0000100011001000000100",
			1749 => "0000001001101110001001",
			1750 => "0000000001101110001001",
			1751 => "0000000001101110001001",
			1752 => "1111111001101110001001",
			1753 => "0010000110011000001000",
			1754 => "0001001000100000000100",
			1755 => "1111111001101110001001",
			1756 => "0000010001101110001001",
			1757 => "0001000011011000000100",
			1758 => "1111111001101110001001",
			1759 => "0001000001101100000100",
			1760 => "0000000001101110001001",
			1761 => "1111111001101110001001",
			1762 => "0001000011011000001100",
			1763 => "0010000110011000001000",
			1764 => "0001001111100100000100",
			1765 => "0000000001101111010101",
			1766 => "0000000001101111010101",
			1767 => "1111111001101111010101",
			1768 => "0011100111111000010000",
			1769 => "0011111010111000001100",
			1770 => "0001011110110000001000",
			1771 => "0000011100100000000100",
			1772 => "0000000001101111010101",
			1773 => "0000000001101111010101",
			1774 => "0000000001101111010101",
			1775 => "0000000001101111010101",
			1776 => "0000101110110100001000",
			1777 => "0010001000101100000100",
			1778 => "0000001001101111010101",
			1779 => "0000000001101111010101",
			1780 => "0000000001101111010101",
			1781 => "0001101101111100011100",
			1782 => "0011011010111100010000",
			1783 => "0011111010111000001100",
			1784 => "0010100110011100000100",
			1785 => "0000000001110000010001",
			1786 => "0001100111101000000100",
			1787 => "0000000001110000010001",
			1788 => "0000000001110000010001",
			1789 => "0000000001110000010001",
			1790 => "0001001111101000000100",
			1791 => "0000000001110000010001",
			1792 => "0001000101001100000100",
			1793 => "0000001001110000010001",
			1794 => "0000000001110000010001",
			1795 => "1111111001110000010001",
			1796 => "0001101101111100011100",
			1797 => "0011011010111100010000",
			1798 => "0011111010111000001100",
			1799 => "0010010110000000001000",
			1800 => "0001101110010100000100",
			1801 => "0000000001110001001101",
			1802 => "0000000001110001001101",
			1803 => "0000000001110001001101",
			1804 => "0000000001110001001101",
			1805 => "0010011110100000000100",
			1806 => "0000000001110001001101",
			1807 => "0001001111101000000100",
			1808 => "0000000001110001001101",
			1809 => "0000000001110001001101",
			1810 => "0000000001110001001101",
			1811 => "0001000011011000001100",
			1812 => "0010000110011000001000",
			1813 => "0000001001101000000100",
			1814 => "0000000001110010100001",
			1815 => "0000001001110010100001",
			1816 => "1111111001110010100001",
			1817 => "0000100111100000010000",
			1818 => "0001001011100100001000",
			1819 => "0000000100000000000100",
			1820 => "0000000001110010100001",
			1821 => "0000000001110010100001",
			1822 => "0000000001001000000100",
			1823 => "0000001001110010100001",
			1824 => "0000000001110010100001",
			1825 => "0000000011010000001000",
			1826 => "0011011011011100000100",
			1827 => "0000000001110010100001",
			1828 => "0000000001110010100001",
			1829 => "0000110111000000000100",
			1830 => "0000000001110010100001",
			1831 => "0000000001110010100001",
			1832 => "0001100001111000100000",
			1833 => "0000110111000000001100",
			1834 => "0001100111101000000100",
			1835 => "0000000001110011111101",
			1836 => "0000000100000100000100",
			1837 => "0000000001110011111101",
			1838 => "0000000001110011111101",
			1839 => "0000110100011000001100",
			1840 => "0011110101101100000100",
			1841 => "0000000001110011111101",
			1842 => "0000011110011100000100",
			1843 => "0000000001110011111101",
			1844 => "0000000001110011111101",
			1845 => "0000001011010100000100",
			1846 => "0000000001110011111101",
			1847 => "0000000001110011111101",
			1848 => "0011011011011100001000",
			1849 => "0000110111000100000100",
			1850 => "0000000001110011111101",
			1851 => "1111111001110011111101",
			1852 => "0001010100000100000100",
			1853 => "0000000001110011111101",
			1854 => "0000000001110011111101",
			1855 => "0001000011011000001100",
			1856 => "0010000110011000001000",
			1857 => "0001001000100000000100",
			1858 => "0000000001110101001001",
			1859 => "0000001001110101001001",
			1860 => "1111111001110101001001",
			1861 => "0011000011011100011000",
			1862 => "0001001011100100001100",
			1863 => "0001111101100000001000",
			1864 => "0000011100100000000100",
			1865 => "0000000001110101001001",
			1866 => "0000000001110101001001",
			1867 => "0000001001110101001001",
			1868 => "0000100011001000001000",
			1869 => "0010100110011100000100",
			1870 => "0000000001110101001001",
			1871 => "0000001001110101001001",
			1872 => "0000000001110101001001",
			1873 => "0000000001110101001001",
			1874 => "0001101101111100011100",
			1875 => "0000110100011000010100",
			1876 => "0000010000011000010000",
			1877 => "0001010011100000001100",
			1878 => "0001101110010100000100",
			1879 => "0000000001110110000101",
			1880 => "0000100011001000000100",
			1881 => "0000001001110110000101",
			1882 => "0000000001110110000101",
			1883 => "0000000001110110000101",
			1884 => "1111111001110110000101",
			1885 => "0001001111101000000100",
			1886 => "0000000001110110000101",
			1887 => "0000001001110110000101",
			1888 => "1111111001110110000101",
			1889 => "0001101101111100100000",
			1890 => "0011011010111100010000",
			1891 => "0010010110000000001100",
			1892 => "0000100011001000001000",
			1893 => "0010100110011100000100",
			1894 => "0000000001110111001001",
			1895 => "0000000001110111001001",
			1896 => "0000000001110111001001",
			1897 => "0000000001110111001001",
			1898 => "0001001011110000000100",
			1899 => "0000000001110111001001",
			1900 => "0010011110100000000100",
			1901 => "0000000001110111001001",
			1902 => "0001100001111000000100",
			1903 => "0000000001110111001001",
			1904 => "0000000001110111001001",
			1905 => "0000000001110111001001",
			1906 => "0001101101111100100000",
			1907 => "0011011010111100010100",
			1908 => "0011111010111000010000",
			1909 => "0010100110011100000100",
			1910 => "0000000001111000001101",
			1911 => "0001101101111100001000",
			1912 => "0001100111101000000100",
			1913 => "0000000001111000001101",
			1914 => "0000000001111000001101",
			1915 => "0000000001111000001101",
			1916 => "0000000001111000001101",
			1917 => "0010011110100000000100",
			1918 => "0000000001111000001101",
			1919 => "0001001111101000000100",
			1920 => "0000000001111000001101",
			1921 => "0000001001111000001101",
			1922 => "0000000001111000001101",
			1923 => "0001101101111100100000",
			1924 => "0000110100011000010100",
			1925 => "0000010000011000010000",
			1926 => "0001010100011000001100",
			1927 => "0000100011001000001000",
			1928 => "0010100110011100000100",
			1929 => "0000000001111001010001",
			1930 => "0000000001111001010001",
			1931 => "0000000001111001010001",
			1932 => "0000000001111001010001",
			1933 => "0000000001111001010001",
			1934 => "0000001011010100000100",
			1935 => "0000000001111001010001",
			1936 => "0011011001001000000100",
			1937 => "0000000001111001010001",
			1938 => "0000000001111001010001",
			1939 => "0000000001111001010001",
			1940 => "0011100001010100001100",
			1941 => "0010101000101100001000",
			1942 => "0011111010111100000100",
			1943 => "0000001001111010101101",
			1944 => "1111111001111010101101",
			1945 => "1111111001111010101101",
			1946 => "0011111101010100010000",
			1947 => "0011001100001000001100",
			1948 => "0001001010101000000100",
			1949 => "1111111001111010101101",
			1950 => "0001110100010100000100",
			1951 => "0000001001111010101101",
			1952 => "0000010001111010101101",
			1953 => "1111111001111010101101",
			1954 => "0001000011011000000100",
			1955 => "1111111001111010101101",
			1956 => "0001101101111100001100",
			1957 => "0001100001111000000100",
			1958 => "1111111001111010101101",
			1959 => "0001001111011000000100",
			1960 => "0000010001111010101101",
			1961 => "1111111001111010101101",
			1962 => "1111111001111010101101",
			1963 => "0011100001010100011000",
			1964 => "0001101101111100010000",
			1965 => "0011111010111000001100",
			1966 => "0001100111101000000100",
			1967 => "0000000001111100001001",
			1968 => "0010001011000100000100",
			1969 => "0000001001111100001001",
			1970 => "0000000001111100001001",
			1971 => "0000000001111100001001",
			1972 => "0001101101111100000100",
			1973 => "0000000001111100001001",
			1974 => "0000000001111100001001",
			1975 => "0001000011011000000100",
			1976 => "1111111001111100001001",
			1977 => "0001101101111100010000",
			1978 => "0011101100001000001100",
			1979 => "0011111101010100001000",
			1980 => "0001001101100100000100",
			1981 => "0000000001111100001001",
			1982 => "0000000001111100001001",
			1983 => "1111111001111100001001",
			1984 => "0000001001111100001001",
			1985 => "1111111001111100001001",
			1986 => "0001000011011000001100",
			1987 => "0010000110011000001000",
			1988 => "0000001011010100000100",
			1989 => "1111111001111101010101",
			1990 => "0000001001111101010101",
			1991 => "1111111001111101010101",
			1992 => "0001101101111100011000",
			1993 => "0001111110001100010100",
			1994 => "0001101110010100000100",
			1995 => "0000000001111101010101",
			1996 => "0000010000011000001000",
			1997 => "0000100011001000000100",
			1998 => "0000001001111101010101",
			1999 => "0000000001111101010101",
			2000 => "0000010110000000000100",
			2001 => "0000000001111101010101",
			2002 => "0000000001111101010101",
			2003 => "0000000001111101010101",
			2004 => "1111111001111101010101",
			2005 => "0001101101111100100100",
			2006 => "0000110100011000011000",
			2007 => "0001001101000000001000",
			2008 => "0010010000011000000100",
			2009 => "0000000001111110100001",
			2010 => "1111111001111110100001",
			2011 => "0001010100011000001100",
			2012 => "0001100111101000000100",
			2013 => "0000000001111110100001",
			2014 => "0000000100000100000100",
			2015 => "0000001001111110100001",
			2016 => "0000000001111110100001",
			2017 => "0000000001111110100001",
			2018 => "0001001111101000000100",
			2019 => "0000000001111110100001",
			2020 => "0011011011000000000100",
			2021 => "0000000001111110100001",
			2022 => "0000001001111110100001",
			2023 => "1111111001111110100001",
			2024 => "0000110111000000010000",
			2025 => "0001001011011000000100",
			2026 => "0000000001111111111101",
			2027 => "0010100010101000001000",
			2028 => "0001100111101000000100",
			2029 => "0000000001111111111101",
			2030 => "0000001001111111111101",
			2031 => "0000000001111111111101",
			2032 => "0010101010100100001000",
			2033 => "0001001111101000000100",
			2034 => "1111111001111111111101",
			2035 => "0000010001111111111101",
			2036 => "0001000011011000000100",
			2037 => "1111111001111111111101",
			2038 => "0001101101111100010000",
			2039 => "0011100111111000001100",
			2040 => "0011110111001000001000",
			2041 => "0000101100100100000100",
			2042 => "0000000001111111111101",
			2043 => "0000000001111111111101",
			2044 => "1111111001111111111101",
			2045 => "0000001001111111111101",
			2046 => "1111111001111111111101",
			2047 => "0001000011011000010000",
			2048 => "0001101110010100001100",
			2049 => "0000101110101000000100",
			2050 => "0000000010000001011001",
			2051 => "0000110001111100000100",
			2052 => "0000000010000001011001",
			2053 => "0000000010000001011001",
			2054 => "1111111010000001011001",
			2055 => "0001101101111100011100",
			2056 => "0001111110001100011000",
			2057 => "0001000000101100001100",
			2058 => "0010101001000100001000",
			2059 => "0010101000010100000100",
			2060 => "0000000010000001011001",
			2061 => "0000000010000001011001",
			2062 => "0000000010000001011001",
			2063 => "0001101110010100000100",
			2064 => "0000000010000001011001",
			2065 => "0000101110110100000100",
			2066 => "0000001010000001011001",
			2067 => "0000000010000001011001",
			2068 => "0000000010000001011001",
			2069 => "0000000010000001011001",
			2070 => "0011100101000100010000",
			2071 => "0011111010111000001100",
			2072 => "0001101101111100001000",
			2073 => "0000110111000000000100",
			2074 => "0000001010000011000101",
			2075 => "0000000010000011000101",
			2076 => "0000000010000011000101",
			2077 => "0000000010000011000101",
			2078 => "0001000011011000001100",
			2079 => "0001101110010100001000",
			2080 => "0001101011111100000100",
			2081 => "1111111010000011000101",
			2082 => "0000000010000011000101",
			2083 => "1111111010000011000101",
			2084 => "0001101101111100011000",
			2085 => "0011101100001000010100",
			2086 => "0011110111001000001000",
			2087 => "0000001000011000000100",
			2088 => "0000001010000011000101",
			2089 => "0000000010000011000101",
			2090 => "0001001010010000000100",
			2091 => "1111111010000011000101",
			2092 => "0000101100010100000100",
			2093 => "0000000010000011000101",
			2094 => "0000000010000011000101",
			2095 => "0000001010000011000101",
			2096 => "1111111010000011000101",
			2097 => "0000110111000000010000",
			2098 => "0001101101111100001000",
			2099 => "0001100111101000000100",
			2100 => "0000000010000101000001",
			2101 => "0000001010000101000001",
			2102 => "0000111010101100000100",
			2103 => "0000000010000101000001",
			2104 => "0000000010000101000001",
			2105 => "0001000011011000001100",
			2106 => "0010000110011000001000",
			2107 => "0000001001101000000100",
			2108 => "1111111010000101000001",
			2109 => "0000010010000101000001",
			2110 => "1111111010000101000001",
			2111 => "0010001111001000010000",
			2112 => "0000101110110100001100",
			2113 => "0011111011011100000100",
			2114 => "0000000010000101000001",
			2115 => "0001011000111100000100",
			2116 => "0000000010000101000001",
			2117 => "0000001010000101000001",
			2118 => "0000000010000101000001",
			2119 => "0001101101111100010000",
			2120 => "0010001000110000000100",
			2121 => "1111111010000101000001",
			2122 => "0000101001011100001000",
			2123 => "0000001001001000000100",
			2124 => "0000001010000101000001",
			2125 => "0000000010000101000001",
			2126 => "0000000010000101000001",
			2127 => "1111111010000101000001",
			2128 => "0011100001110000010000",
			2129 => "0001101101111100001100",
			2130 => "0011111010111100001000",
			2131 => "0000000001000000000100",
			2132 => "0000001010000111000101",
			2133 => "0000000010000111000101",
			2134 => "1111111010000111000101",
			2135 => "1111111010000111000101",
			2136 => "0011111010111000001100",
			2137 => "0001011010111100001000",
			2138 => "0001001011100100000100",
			2139 => "1111111010000111000101",
			2140 => "0000001010000111000101",
			2141 => "1111111010000111000101",
			2142 => "0001000011011000001100",
			2143 => "0001101110010100001000",
			2144 => "0001101011111100000100",
			2145 => "1111111010000111000101",
			2146 => "0000001010000111000101",
			2147 => "1111111010000111000101",
			2148 => "0010001111001000001100",
			2149 => "0001010110100100000100",
			2150 => "1111111010000111000101",
			2151 => "0010110111001000000100",
			2152 => "0000011010000111000101",
			2153 => "0000000010000111000101",
			2154 => "0001101101111100001100",
			2155 => "0001011100101000000100",
			2156 => "1111111010000111000101",
			2157 => "0001011010011100000100",
			2158 => "0000010010000111000101",
			2159 => "1111111010000111000101",
			2160 => "1111111010000111000101",
			2161 => "0000110111000000010100",
			2162 => "0001001011011000000100",
			2163 => "0000000010001001010001",
			2164 => "0010100010101000001100",
			2165 => "0011000000101000001000",
			2166 => "0011110111001000000100",
			2167 => "0000001010001001010001",
			2168 => "0000000010001001010001",
			2169 => "0000001010001001010001",
			2170 => "0000000010001001010001",
			2171 => "0001000011011000001100",
			2172 => "0010101010100100001000",
			2173 => "0001001111101000000100",
			2174 => "1111111010001001010001",
			2175 => "0001000010001001010001",
			2176 => "1111111010001001010001",
			2177 => "0000101110000100010000",
			2178 => "0010111100001000001000",
			2179 => "0011111010111100000100",
			2180 => "0000001010001001010001",
			2181 => "1111111010001001010001",
			2182 => "0011000110000100000100",
			2183 => "0000010010001001010001",
			2184 => "0000000010001001010001",
			2185 => "0000101010001000010100",
			2186 => "0000101001011100001100",
			2187 => "0000100101001000001000",
			2188 => "0011000111111000000100",
			2189 => "0000000010001001010001",
			2190 => "0000000010001001010001",
			2191 => "1111111010001001010001",
			2192 => "0010101100000100000100",
			2193 => "0000001010001001010001",
			2194 => "0000000010001001010001",
			2195 => "1111111010001001010001",
			2196 => "0011100001010100010000",
			2197 => "0001101101111100001100",
			2198 => "0011111010111100001000",
			2199 => "0000000111100000000100",
			2200 => "0000001010001011011101",
			2201 => "1111111010001011011101",
			2202 => "1111111010001011011101",
			2203 => "1111111010001011011101",
			2204 => "0011111010111000010000",
			2205 => "0001110000101000001100",
			2206 => "0000011100100000001000",
			2207 => "0011110000001100000100",
			2208 => "0000001010001011011101",
			2209 => "0000010010001011011101",
			2210 => "1111111010001011011101",
			2211 => "1111111010001011011101",
			2212 => "0001000011011000001100",
			2213 => "0001101110010100001000",
			2214 => "0001101011111100000100",
			2215 => "1111111010001011011101",
			2216 => "0000001010001011011101",
			2217 => "1111111010001011011101",
			2218 => "0000100111100000001000",
			2219 => "0001101101111100000100",
			2220 => "0000001010001011011101",
			2221 => "0000000010001011011101",
			2222 => "0000101110110100010000",
			2223 => "0000101110110100001000",
			2224 => "0001001010010000000100",
			2225 => "1111111010001011011101",
			2226 => "0000000010001011011101",
			2227 => "0001000001001100000100",
			2228 => "0000011010001011011101",
			2229 => "1111111010001011011101",
			2230 => "1111111010001011011101",
			2231 => "0000111000101100010100",
			2232 => "0001101101111100010000",
			2233 => "0001101110010100000100",
			2234 => "1111111010001101111011",
			2235 => "0000000101001000001000",
			2236 => "0011110001111100000100",
			2237 => "0000001010001101111011",
			2238 => "0000000010001101111011",
			2239 => "0000000010001101111011",
			2240 => "1111111010001101111011",
			2241 => "0011111010111000010000",
			2242 => "0011011100101100001100",
			2243 => "0000011100100000001000",
			2244 => "0011110001111100000100",
			2245 => "0000001010001101111011",
			2246 => "0000100010001101111011",
			2247 => "1111111010001101111011",
			2248 => "1111111010001101111011",
			2249 => "0001000011011000001100",
			2250 => "0001101110010100001000",
			2251 => "0001101011111100000100",
			2252 => "1111111010001101111011",
			2253 => "0000001010001101111011",
			2254 => "1111111010001101111011",
			2255 => "0000100111100000001000",
			2256 => "0001101101111100000100",
			2257 => "0000001010001101111011",
			2258 => "0000000010001101111011",
			2259 => "0001000001101100001100",
			2260 => "0000101110110100000100",
			2261 => "1111111010001101111011",
			2262 => "0001101011001100000100",
			2263 => "0000010010001101111011",
			2264 => "0000000010001101111011",
			2265 => "0001101101111100001000",
			2266 => "0001101101111100000100",
			2267 => "1111111010001101111011",
			2268 => "0000001010001101111011",
			2269 => "1111111010001101111011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(736, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1502, initial_addr_3'length));
	end generate gen_rom_6;

	gen_rom_7: if SELECT_ROM = 7 generate
		bank <= (
			0 => "0001000110110001101000",
			1 => "0010011100011000111000",
			2 => "0011111110110100101000",
			3 => "0001001010000100001000",
			4 => "0001110100010100000100",
			5 => "0000000000000100010101",
			6 => "1111111000000100010101",
			7 => "0010010110101000010000",
			8 => "0011000100010100001000",
			9 => "0010010010001100000100",
			10 => "0000000000000100010101",
			11 => "0000000000000100010101",
			12 => "0011100100010100000100",
			13 => "0000000000000100010101",
			14 => "1111111000000100010101",
			15 => "0000011110100000001000",
			16 => "0011101100110000000100",
			17 => "0000001000000100010101",
			18 => "0000000000000100010101",
			19 => "0001100111101000000100",
			20 => "0000001000000100010101",
			21 => "0000000000000100010101",
			22 => "0001011000011000001000",
			23 => "0010011011111100000100",
			24 => "0000001000000100010101",
			25 => "1111111000000100010101",
			26 => "0000100101010100000100",
			27 => "0000001000000100010101",
			28 => "0000000000000100010101",
			29 => "0001101001111100011100",
			30 => "0010100001010000000100",
			31 => "1111111000000100010101",
			32 => "0011000100011000001100",
			33 => "0000100110001100001000",
			34 => "0001100100111100000100",
			35 => "0000000000000100010101",
			36 => "1111111000000100010101",
			37 => "0000000000000100010101",
			38 => "0011110101000000001000",
			39 => "0001001011100000000100",
			40 => "0000001000000100010101",
			41 => "0000000000000100010101",
			42 => "1111111000000100010101",
			43 => "0011100010110000001100",
			44 => "0001001110111000000100",
			45 => "0000000000000100010101",
			46 => "0011001000000000000100",
			47 => "0000000000000100010101",
			48 => "0000001000000100010101",
			49 => "0011000001011000000100",
			50 => "1111111000000100010101",
			51 => "0000000000000100010101",
			52 => "0001101011001100001100",
			53 => "0001000011111000000100",
			54 => "1111111000000100010101",
			55 => "0001001110011000000100",
			56 => "0000000000000100010101",
			57 => "1111111000000100010101",
			58 => "0000100010000100001000",
			59 => "0000011110011100000100",
			60 => "0000000000000100010101",
			61 => "0000001000000100010101",
			62 => "0010101100000100001100",
			63 => "0010001111000100000100",
			64 => "1111111000000100010101",
			65 => "0001000101100000000100",
			66 => "0000001000000100010101",
			67 => "0000000000000100010101",
			68 => "1111111000000100010101",
			69 => "0001111100101000111100",
			70 => "0000011100100000001000",
			71 => "0001101011001100000100",
			72 => "1111111000001000011001",
			73 => "0000000000001000011001",
			74 => "0001100001000100000100",
			75 => "1111111000001000011001",
			76 => "0001100100111100100000",
			77 => "0011100100010100010000",
			78 => "0001010101101100001000",
			79 => "0000111011000100000100",
			80 => "0000000000001000011001",
			81 => "0000000000001000011001",
			82 => "0001100001111000000100",
			83 => "0000001000001000011001",
			84 => "0000000000001000011001",
			85 => "0011111011011100001000",
			86 => "0001100111101000000100",
			87 => "0000001000001000011001",
			88 => "0000000000001000011001",
			89 => "0011000100000000000100",
			90 => "0000000000001000011001",
			91 => "0000000000001000011001",
			92 => "0011001100110000001100",
			93 => "0010101001101000001000",
			94 => "0010110111001000000100",
			95 => "1111111000001000011001",
			96 => "0000000000001000011001",
			97 => "0000001000001000011001",
			98 => "0000001000001000011001",
			99 => "0010001001101000010000",
			100 => "0000011011101000001100",
			101 => "0000011011101000000100",
			102 => "1111111000001000011001",
			103 => "0001010001011000000100",
			104 => "1111111000001000011001",
			105 => "0000001000001000011001",
			106 => "1111111000001000011001",
			107 => "0010000010011000101100",
			108 => "0011101101101100010100",
			109 => "0010010111101100010000",
			110 => "0011111100010000001000",
			111 => "0011010001011000000100",
			112 => "0000001000001000011001",
			113 => "1111111000001000011001",
			114 => "0001100100111100000100",
			115 => "0000010000001000011001",
			116 => "0000000000001000011001",
			117 => "1111111000001000011001",
			118 => "0001101001111100001000",
			119 => "0010001001101000000100",
			120 => "0000000000001000011001",
			121 => "1111111000001000011001",
			122 => "0011000111010000001000",
			123 => "0010100110011100000100",
			124 => "1111111000001000011001",
			125 => "0000000000001000011001",
			126 => "0011111010110100000100",
			127 => "0000010000001000011001",
			128 => "0000000000001000011001",
			129 => "0010000000110000001000",
			130 => "0010000000110000000100",
			131 => "1111111000001000011001",
			132 => "0000001000001000011001",
			133 => "1111111000001000011001",
			134 => "0011000000001101100000",
			135 => "0000010000011000010000",
			136 => "0000100001001000001000",
			137 => "0001100001111000000100",
			138 => "1111111000001100111101",
			139 => "0000001000001100111101",
			140 => "0001101011001100000100",
			141 => "1111111000001100111101",
			142 => "0000000000001100111101",
			143 => "0001000000010000010000",
			144 => "0011101000111000000100",
			145 => "0000000000001100111101",
			146 => "0010111110001100000100",
			147 => "1111111000001100111101",
			148 => "0010111101111000000100",
			149 => "0000000000001100111101",
			150 => "1111111000001100111101",
			151 => "0011000000101000100000",
			152 => "0011000100010100010000",
			153 => "0011000100010100001000",
			154 => "0000110100010100000100",
			155 => "0000000000001100111101",
			156 => "0000000000001100111101",
			157 => "0001000001101100000100",
			158 => "0000000000001100111101",
			159 => "1111111000001100111101",
			160 => "0001000100001100001000",
			161 => "0011000100010100000100",
			162 => "0000000000001100111101",
			163 => "0000000000001100111101",
			164 => "0011000100010100000100",
			165 => "0000000000001100111101",
			166 => "0000001000001100111101",
			167 => "0011000000101000010000",
			168 => "0010100001010000001000",
			169 => "0000100010000000000100",
			170 => "0000001000001100111101",
			171 => "0000010000001100111101",
			172 => "0001000010111000000100",
			173 => "1111111000001100111101",
			174 => "0000000000001100111101",
			175 => "0011000000101000001000",
			176 => "0011110101110100000100",
			177 => "0000000000001100111101",
			178 => "1111111000001100111101",
			179 => "0011101001110000000100",
			180 => "0000001000001100111101",
			181 => "0000000000001100111101",
			182 => "0010001001101000001000",
			183 => "0011100100000100000100",
			184 => "0000001000001100111101",
			185 => "1111111000001100111101",
			186 => "0001000110110000101000",
			187 => "0010000110001000010000",
			188 => "0000100101000000001100",
			189 => "0001001001001100001000",
			190 => "0001000010111000000100",
			191 => "0000000000001100111101",
			192 => "0000010000001100111101",
			193 => "1111111000001100111101",
			194 => "1111111000001100111101",
			195 => "0001000011101100001100",
			196 => "0001000101010100000100",
			197 => "0000000000001100111101",
			198 => "0011000111001000000100",
			199 => "0000000000001100111101",
			200 => "0000001000001100111101",
			201 => "0010000001110100000100",
			202 => "1111111000001100111101",
			203 => "0001100101010000000100",
			204 => "1111111000001100111101",
			205 => "0000001000001100111101",
			206 => "1111111000001100111101",
			207 => "0001111101111001100100",
			208 => "0001000001100101001000",
			209 => "0001100001000100001000",
			210 => "0001100001000100000100",
			211 => "1111111000010010000001",
			212 => "0000000000010010000001",
			213 => "0011101000111100100000",
			214 => "0010111100001000010000",
			215 => "0000110100000000001000",
			216 => "0001110111111000000100",
			217 => "0000000000010010000001",
			218 => "0000001000010010000001",
			219 => "0011110010001000000100",
			220 => "0000000000010010000001",
			221 => "0000001000010010000001",
			222 => "0001000101010100001000",
			223 => "0001100100110100000100",
			224 => "0000001000010010000001",
			225 => "0000000000010010000001",
			226 => "0010010111100100000100",
			227 => "0000001000010010000001",
			228 => "0000001000010010000001",
			229 => "0001000010111000010000",
			230 => "0001111000111000001000",
			231 => "0001101100011000000100",
			232 => "0000000000010010000001",
			233 => "1111111000010010000001",
			234 => "0010010001111000000100",
			235 => "0000001000010010000001",
			236 => "1111111000010010000001",
			237 => "0001101011001100001000",
			238 => "0010011101101000000100",
			239 => "0000000000010010000001",
			240 => "0000001000010010000001",
			241 => "0001111101100000000100",
			242 => "0000000000010010000001",
			243 => "0000001000010010000001",
			244 => "0001100100110100001000",
			245 => "0011011100101100000100",
			246 => "1111111000010010000001",
			247 => "0000000000010010000001",
			248 => "0001010100001000001100",
			249 => "0001101100011000000100",
			250 => "0000000000010010000001",
			251 => "0000001101111000000100",
			252 => "0000000000010010000001",
			253 => "0000001000010010000001",
			254 => "0011110110010000000100",
			255 => "1111111000010010000001",
			256 => "0000001000010010000001",
			257 => "0010001001101000001100",
			258 => "0001110001111100001000",
			259 => "0001110001111100000100",
			260 => "1111111000010010000001",
			261 => "0000001000010010000001",
			262 => "1111111000010010000001",
			263 => "0001000010010000110000",
			264 => "0010001111001000011000",
			265 => "0011111000000100001100",
			266 => "0001000100001100001000",
			267 => "0001000011001100000100",
			268 => "0000000000010010000001",
			269 => "0000010000010010000001",
			270 => "1111111000010010000001",
			271 => "0010001001101000000100",
			272 => "0000000000010010000001",
			273 => "0001110111110000000100",
			274 => "1111111000010010000001",
			275 => "0000000000010010000001",
			276 => "0011110000010100010000",
			277 => "0001001001001100001000",
			278 => "0010100110011100000100",
			279 => "0000000000010010000001",
			280 => "1111111000010010000001",
			281 => "0000000000111000000100",
			282 => "0000011000010010000001",
			283 => "0000001000010010000001",
			284 => "0001100100101100000100",
			285 => "1111111000010010000001",
			286 => "0000001000010010000001",
			287 => "1111111000010010000001",
			288 => "0001111110001101100100",
			289 => "0001000110110001000100",
			290 => "0001100001000100000100",
			291 => "1111111000010111001101",
			292 => "0001000100001100100000",
			293 => "0010101010110000010000",
			294 => "0000100010000000001000",
			295 => "0001100100110100000100",
			296 => "0000000000010111001101",
			297 => "0000000000010111001101",
			298 => "0001101010011000000100",
			299 => "0000001000010111001101",
			300 => "0000000000010111001101",
			301 => "0000101100010100001000",
			302 => "0010011101101000000100",
			303 => "0000000000010111001101",
			304 => "0000001000010111001101",
			305 => "0011000100000000000100",
			306 => "0000000000010111001101",
			307 => "0000000000010111001101",
			308 => "0010011001111000010000",
			309 => "0000111000111000001000",
			310 => "0000110000111000000100",
			311 => "0000001000010111001101",
			312 => "0000000000010111001101",
			313 => "0010110100010100000100",
			314 => "0000001000010111001101",
			315 => "1111111000010111001101",
			316 => "0001011101010100001000",
			317 => "0000111001110000000100",
			318 => "0000001000010111001101",
			319 => "0000000000010111001101",
			320 => "0011110010000000000100",
			321 => "0000000000010111001101",
			322 => "0000001000010111001101",
			323 => "0000011110100000011000",
			324 => "0010011110100000010100",
			325 => "0000011100100000000100",
			326 => "1111111000010111001101",
			327 => "0001011000111100001000",
			328 => "0001001110011000000100",
			329 => "1111111000010111001101",
			330 => "0000000000010111001101",
			331 => "0000101001011100000100",
			332 => "0000001000010111001101",
			333 => "1111111000010111001101",
			334 => "1111111000010111001101",
			335 => "0001000001001100000100",
			336 => "0000000000010111001101",
			337 => "1111111000010111001101",
			338 => "0010001001101000010000",
			339 => "0000011011101000001100",
			340 => "0000011011101000000100",
			341 => "1111111000010111001101",
			342 => "0010110100011000000100",
			343 => "1111111000010111001101",
			344 => "0000001000010111001101",
			345 => "1111111000010111001101",
			346 => "0001000010010000100100",
			347 => "0010100001010100011100",
			348 => "0001100100111100001100",
			349 => "0001100100111100001000",
			350 => "0000011101101000000100",
			351 => "0000001000010111001101",
			352 => "1111111000010111001101",
			353 => "0000001000010111001101",
			354 => "0001111111011100001000",
			355 => "0010001001101000000100",
			356 => "0000000000010111001101",
			357 => "1111111000010111001101",
			358 => "0001000000010100000100",
			359 => "0000001000010111001101",
			360 => "0000000000010111001101",
			361 => "0010100001110000000100",
			362 => "0000000000010111001101",
			363 => "0000001000010111001101",
			364 => "0001000000000000001100",
			365 => "0010000000110000000100",
			366 => "1111111000010111001101",
			367 => "0010100001110100000100",
			368 => "0000001000010111001101",
			369 => "1111111000010111001101",
			370 => "1111111000010111001101",
			371 => "0001111110001101111100",
			372 => "0000010000011000010000",
			373 => "0000100001001000001000",
			374 => "0001000101001100000100",
			375 => "0000001000011101011001",
			376 => "1111111000011101011001",
			377 => "0010100010101000000100",
			378 => "1111111000011101011001",
			379 => "0000000000011101011001",
			380 => "0001110100010100111100",
			381 => "0000110000101000100000",
			382 => "0001011000111100010000",
			383 => "0000111010000000001000",
			384 => "0000001100001000000100",
			385 => "0000000000011101011001",
			386 => "0000001000011101011001",
			387 => "0001011000111100000100",
			388 => "0000000000011101011001",
			389 => "1111111000011101011001",
			390 => "0010100101000100001000",
			391 => "0010011100110100000100",
			392 => "0000000000011101011001",
			393 => "0000001000011101011001",
			394 => "0011100111000000000100",
			395 => "0000000000011101011001",
			396 => "1111111000011101011001",
			397 => "0010010010001100001100",
			398 => "0011000100010100001000",
			399 => "0011100010111100000100",
			400 => "0000000000011101011001",
			401 => "1111111000011101011001",
			402 => "0000001000011101011001",
			403 => "0000111000111000001000",
			404 => "0010110111111000000100",
			405 => "1111111000011101011001",
			406 => "0000000000011101011001",
			407 => "0000101110010000000100",
			408 => "1111111000011101011001",
			409 => "0000000000011101011001",
			410 => "0001000000010000010000",
			411 => "0011101000111000000100",
			412 => "0000000000011101011001",
			413 => "0001110101101100000100",
			414 => "1111111000011101011001",
			415 => "0001110101101100000100",
			416 => "0000000000011101011001",
			417 => "1111111000011101011001",
			418 => "0010100111110100010000",
			419 => "0011010110000100001000",
			420 => "0011101010000000000100",
			421 => "0000000000011101011001",
			422 => "1111110000011101011001",
			423 => "0001001011101100000100",
			424 => "0000000000011101011001",
			425 => "0000001000011101011001",
			426 => "0011101000111000001000",
			427 => "0010010111100100000100",
			428 => "0000000000011101011001",
			429 => "0000001000011101011001",
			430 => "0000100100101000000100",
			431 => "0000000000011101011001",
			432 => "0000000000011101011001",
			433 => "0010100001010000011000",
			434 => "0011101010001100001100",
			435 => "0011010101100100001000",
			436 => "0011101011000000000100",
			437 => "0000000000011101011001",
			438 => "1111111000011101011001",
			439 => "0000001000011101011001",
			440 => "0010010001111000001000",
			441 => "0010010001111000000100",
			442 => "1111111000011101011001",
			443 => "0000000000011101011001",
			444 => "1111111000011101011001",
			445 => "0001000001001100101000",
			446 => "0010100001010100011100",
			447 => "0000101000101000001100",
			448 => "0001000011011000001000",
			449 => "0011111100010000000100",
			450 => "0000000000011101011001",
			451 => "0000001000011101011001",
			452 => "1111111000011101011001",
			453 => "0001111111011100001000",
			454 => "0010010101010000000100",
			455 => "0000000000011101011001",
			456 => "1111111000011101011001",
			457 => "0011110010111000000100",
			458 => "0000001000011101011001",
			459 => "0000000000011101011001",
			460 => "0010101100000100001000",
			461 => "0011110000010100000100",
			462 => "0000001000011101011001",
			463 => "1111111000011101011001",
			464 => "0000010000011101011001",
			465 => "0001000000000000001000",
			466 => "0001001010101000000100",
			467 => "1111111000011101011001",
			468 => "0000000000011101011001",
			469 => "1111111000011101011001",
			470 => "0001000000101110011000",
			471 => "0001010100011000111100",
			472 => "0001111101100000101000",
			473 => "0000010110101000100000",
			474 => "0011111011011100010000",
			475 => "0011100000111000001000",
			476 => "0010110100010100000100",
			477 => "0000000000100100000101",
			478 => "0000000000100100000101",
			479 => "0010100001010000000100",
			480 => "0000000000100100000101",
			481 => "0000000000100100000101",
			482 => "0001100100110100001000",
			483 => "0001010100001000000100",
			484 => "0000000000100100000101",
			485 => "0000001000100100000101",
			486 => "0011001010000000000100",
			487 => "0000001000100100000101",
			488 => "0000000000100100000101",
			489 => "0001001000000100000100",
			490 => "0000001000100100000101",
			491 => "0000000000100100000101",
			492 => "0011111110000100001100",
			493 => "0001101100011000001000",
			494 => "0011101101111000000100",
			495 => "0000001000100100000101",
			496 => "1111111000100100000101",
			497 => "0000001000100100000101",
			498 => "0011001000111000000100",
			499 => "1111111000100100000101",
			500 => "0000001000100100000101",
			501 => "0010100110011000101100",
			502 => "0000100101110000011100",
			503 => "0000101111010000001100",
			504 => "0011110101110100001000",
			505 => "0011110110110100000100",
			506 => "1111111000100100000101",
			507 => "0000000000100100000101",
			508 => "1111111000100100000101",
			509 => "0000100010011100001000",
			510 => "0001100111101000000100",
			511 => "0000000000100100000101",
			512 => "0000001000100100000101",
			513 => "0000100101110000000100",
			514 => "1111111000100100000101",
			515 => "0000001000100100000101",
			516 => "0001010011100000000100",
			517 => "1111111000100100000101",
			518 => "0001011000000000000100",
			519 => "0000001000100100000101",
			520 => "0010001011010100000100",
			521 => "1111111000100100000101",
			522 => "1111110000100100000101",
			523 => "0011001000111000010100",
			524 => "0011100001101000000100",
			525 => "1111111000100100000101",
			526 => "0001101001100100001000",
			527 => "0000010111100100000100",
			528 => "0000001000100100000101",
			529 => "1111111000100100000101",
			530 => "0011111100010000000100",
			531 => "1111111000100100000101",
			532 => "0000000000100100000101",
			533 => "0000000010111100010000",
			534 => "0011110101000000001000",
			535 => "0001000010111000000100",
			536 => "0000000000100100000101",
			537 => "0000001000100100000101",
			538 => "0010101100011100000100",
			539 => "1111111000100100000101",
			540 => "0000001000100100000101",
			541 => "0011001000111000000100",
			542 => "0000001000100100000101",
			543 => "0011001100110000000100",
			544 => "0000000000100100000101",
			545 => "0000000000100100000101",
			546 => "0010001101010000100000",
			547 => "0000010110000000001100",
			548 => "0001000110110000001000",
			549 => "0000010000011000000100",
			550 => "0000000000100100000101",
			551 => "0000001000100100000101",
			552 => "1111111000100100000101",
			553 => "0011000000101000000100",
			554 => "1111110000100100000101",
			555 => "0000001100001000000100",
			556 => "1111111000100100000101",
			557 => "0001101011001100000100",
			558 => "0000000000100100000101",
			559 => "0000011011101000000100",
			560 => "0000000000100100000101",
			561 => "0000000000100100000101",
			562 => "0001000101100000011000",
			563 => "0000000011011100001000",
			564 => "0000011011101000000100",
			565 => "1111111000100100000101",
			566 => "0000000000100100000101",
			567 => "0011011000111000000100",
			568 => "0000000000100100000101",
			569 => "0010110000101000000100",
			570 => "0000001000100100000101",
			571 => "0001111000111000000100",
			572 => "1111111000100100000101",
			573 => "0000000000100100000101",
			574 => "0011000000111000000100",
			575 => "0000000000100100000101",
			576 => "1111111000100100000101",
			577 => "0001000110110010011100",
			578 => "0010011100011001101000",
			579 => "0000101001010000111000",
			580 => "0011101000111000011000",
			581 => "0011011100101000001100",
			582 => "0001110100000000001000",
			583 => "0001100111101000000100",
			584 => "0000000000101010011001",
			585 => "0000000000101010011001",
			586 => "1111111000101010011001",
			587 => "0000010010001100001000",
			588 => "0000101111010000000100",
			589 => "0000001000101010011001",
			590 => "0000000000101010011001",
			591 => "1111111000101010011001",
			592 => "0010010111100100010000",
			593 => "0000111100101100001000",
			594 => "0010010110101000000100",
			595 => "1111111000101010011001",
			596 => "0000001000101010011001",
			597 => "0001010110000100000100",
			598 => "0000000000101010011001",
			599 => "1111111000101010011001",
			600 => "0001011101111000001000",
			601 => "0011100101101100000100",
			602 => "0000001000101010011001",
			603 => "0000000000101010011001",
			604 => "0000000010011000000100",
			605 => "0000000000101010011001",
			606 => "1111111000101010011001",
			607 => "0000100010011100010000",
			608 => "0001100001111000000100",
			609 => "0000000000101010011001",
			610 => "0000000010111100000100",
			611 => "0000010000101010011001",
			612 => "0001111100001000000100",
			613 => "0000001000101010011001",
			614 => "0000000000101010011001",
			615 => "0010000111000000010000",
			616 => "0000010110000000001000",
			617 => "0001011000111000000100",
			618 => "1111111000101010011001",
			619 => "0000000000101010011001",
			620 => "0010000110001000000100",
			621 => "0000000000101010011001",
			622 => "0000000000101010011001",
			623 => "0011110101100100001000",
			624 => "0010111011000100000100",
			625 => "0000001000101010011001",
			626 => "1111111000101010011001",
			627 => "0001101011001100000100",
			628 => "0000001000101010011001",
			629 => "0000000000101010011001",
			630 => "0001101001111100100000",
			631 => "0010001001101000000100",
			632 => "1111111000101010011001",
			633 => "0001110110100100001100",
			634 => "0000101100001100001000",
			635 => "0001100100111100000100",
			636 => "0000000000101010011001",
			637 => "1111111000101010011001",
			638 => "0000000000101010011001",
			639 => "0000101100001100001000",
			640 => "0010010100101100000100",
			641 => "0000001000101010011001",
			642 => "0000000000101010011001",
			643 => "0010010100101100000100",
			644 => "0000000000101010011001",
			645 => "1111111000101010011001",
			646 => "0011100010110000001100",
			647 => "0001001110111000000100",
			648 => "0000000000101010011001",
			649 => "0001111111011100000100",
			650 => "0000000000101010011001",
			651 => "0000001000101010011001",
			652 => "0001111001010100000100",
			653 => "1111111000101010011001",
			654 => "0000000000101010011001",
			655 => "0001101011001100010100",
			656 => "0001000011111000000100",
			657 => "1111111000101010011001",
			658 => "0001001101000000001000",
			659 => "0010010110000000000100",
			660 => "0000000000101010011001",
			661 => "0000000000101010011001",
			662 => "0000010000011000000100",
			663 => "1111111000101010011001",
			664 => "0000000000101010011001",
			665 => "0000100010000100001000",
			666 => "0000011110011100000100",
			667 => "0000000000101010011001",
			668 => "0000001000101010011001",
			669 => "0010000010011000010000",
			670 => "0010001111000100000100",
			671 => "1111111000101010011001",
			672 => "0000100010010100000100",
			673 => "0000000000101010011001",
			674 => "0000011011101000000100",
			675 => "0000001000101010011001",
			676 => "0000000000101010011001",
			677 => "1111111000101010011001",
			678 => "0001001011101100011000",
			679 => "0001100001111000010100",
			680 => "0010011101101000001000",
			681 => "0001011100101100000100",
			682 => "1111111000110000000101",
			683 => "0000000000110000000101",
			684 => "0000001011010100000100",
			685 => "1111111000110000000101",
			686 => "0001110100000000000100",
			687 => "0000000000110000000101",
			688 => "0000001000110000000101",
			689 => "1111111000110000000101",
			690 => "0001000011011001011000",
			691 => "0000001100001000110100",
			692 => "0001011000111100010100",
			693 => "0001011000111100010000",
			694 => "0000101110000100001000",
			695 => "0001100001111000000100",
			696 => "0000000000110000000101",
			697 => "0000001000110000000101",
			698 => "0000110100010100000100",
			699 => "1111111000110000000101",
			700 => "1111111000110000000101",
			701 => "1111110000110000000101",
			702 => "0010110111111000010000",
			703 => "0001000000010100001000",
			704 => "0000110100000000000100",
			705 => "0000001000110000000101",
			706 => "0000000000110000000101",
			707 => "0001110111111000000100",
			708 => "0000000000110000000101",
			709 => "0000001000110000000101",
			710 => "0010110111111000001000",
			711 => "0011000111111000000100",
			712 => "1111110000110000000101",
			713 => "0000000000110000000101",
			714 => "0010010110101000000100",
			715 => "0000000000110000000101",
			716 => "0000000000110000000101",
			717 => "0011100000101000011000",
			718 => "0010110111111000001100",
			719 => "0001011000111100001000",
			720 => "0001011000111100000100",
			721 => "0000001000110000000101",
			722 => "0000000000110000000101",
			723 => "1111111000110000000101",
			724 => "0010100001010100001000",
			725 => "0001110000101000000100",
			726 => "0000001000110000000101",
			727 => "0000001000110000000101",
			728 => "0000000000110000000101",
			729 => "0011100100000000000100",
			730 => "1111111000110000000101",
			731 => "0000010010001100000100",
			732 => "0000001000110000000101",
			733 => "0000000000110000000101",
			734 => "0011111001010100100100",
			735 => "0011101011000100100000",
			736 => "0001110111111000010000",
			737 => "0010101001101000001000",
			738 => "0010111110111100000100",
			739 => "1111111000110000000101",
			740 => "1111110000110000000101",
			741 => "0001010100000000000100",
			742 => "0000000000110000000101",
			743 => "0000000000110000000101",
			744 => "0011000111111000001000",
			745 => "0001000110110000000100",
			746 => "0000001000110000000101",
			747 => "0000000000110000000101",
			748 => "0000100011001000000100",
			749 => "1111111000110000000101",
			750 => "0000000000110000000101",
			751 => "1111110000110000000101",
			752 => "0001111101111000010100",
			753 => "0000101100010000001000",
			754 => "0000111101111000000100",
			755 => "0000001000110000000101",
			756 => "1111111000110000000101",
			757 => "0000001100001000000100",
			758 => "0000000000110000000101",
			759 => "0001000001001100000100",
			760 => "0000001000110000000101",
			761 => "0000000000110000000101",
			762 => "0000000100010100000100",
			763 => "1111111000110000000101",
			764 => "0000011001011000001000",
			765 => "0000111101000100000100",
			766 => "0000000000110000000101",
			767 => "1111111000110000000101",
			768 => "0000001000110000000101",
			769 => "0010000111000001110000",
			770 => "0000100010110100101100",
			771 => "0001101101111100101000",
			772 => "0010101000010100010100",
			773 => "0000101110101100001100",
			774 => "0001100001111000001000",
			775 => "0001001011110000000100",
			776 => "0000000000110110001001",
			777 => "0000000000110110001001",
			778 => "0000000000110110001001",
			779 => "0001100111101000000100",
			780 => "0000000000110110001001",
			781 => "1111111000110110001001",
			782 => "0011010110000100010000",
			783 => "0001100001111000001000",
			784 => "0011010011011100000100",
			785 => "0000000000110110001001",
			786 => "0000001000110110001001",
			787 => "0001101101111100000100",
			788 => "1111111000110110001001",
			789 => "0000000000110110001001",
			790 => "0000001000110110001001",
			791 => "1111111000110110001001",
			792 => "0000100010110100001000",
			793 => "0011111000011000000100",
			794 => "0000001000110110001001",
			795 => "0000000000110110001001",
			796 => "0001000010110000011100",
			797 => "0000111000111000001100",
			798 => "0011110100000100001000",
			799 => "0011100000110000000100",
			800 => "0000001000110110001001",
			801 => "0000000000110110001001",
			802 => "0000001000110110001001",
			803 => "0011010101101100001000",
			804 => "0001100111101000000100",
			805 => "1111111000110110001001",
			806 => "0000000000110110001001",
			807 => "0000110110000100000100",
			808 => "0000000000110110001001",
			809 => "0000000000110110001001",
			810 => "0001000010110000010000",
			811 => "0010010111100100001000",
			812 => "0001100111101000000100",
			813 => "0000001000110110001001",
			814 => "1111111000110110001001",
			815 => "0011011101111000000100",
			816 => "0000001000110110001001",
			817 => "0000000000110110001001",
			818 => "0001001000001000001000",
			819 => "0011000011011100000100",
			820 => "0000001000110110001001",
			821 => "1111111000110110001001",
			822 => "0001011010111100000100",
			823 => "0000000000110110001001",
			824 => "0000000000110110001001",
			825 => "0010100101000100010000",
			826 => "0001101010011000001000",
			827 => "0000010000011000000100",
			828 => "0000000000110110001001",
			829 => "0000001000110110001001",
			830 => "0000101100010100000100",
			831 => "0000000000110110001001",
			832 => "0000000000110110001001",
			833 => "0011000000110000001000",
			834 => "0010101011010100000100",
			835 => "1111111000110110001001",
			836 => "0000000000110110001001",
			837 => "0001101100011000100000",
			838 => "0001110100010100010000",
			839 => "0001110111111000001000",
			840 => "0011101100011100000100",
			841 => "0000000000110110001001",
			842 => "1111111000110110001001",
			843 => "0000010000011000000100",
			844 => "0000000000110110001001",
			845 => "0000001000110110001001",
			846 => "0000100111111100001000",
			847 => "0010000010111100000100",
			848 => "1111111000110110001001",
			849 => "0000000000110110001001",
			850 => "0011000110000100000100",
			851 => "0000000000110110001001",
			852 => "0000000000110110001001",
			853 => "0001001011100000001100",
			854 => "0001000011101100001000",
			855 => "0001101011001100000100",
			856 => "0000001000110110001001",
			857 => "0000000000110110001001",
			858 => "1111111000110110001001",
			859 => "0001000110110000001000",
			860 => "0010001000101100000100",
			861 => "0000000000110110001001",
			862 => "0000001000110110001001",
			863 => "0010000011010000000100",
			864 => "0000000000110110001001",
			865 => "0000000000110110001001",
			866 => "0001111101111010011000",
			867 => "0000010000011000100000",
			868 => "0000011100100000000100",
			869 => "1111111000111100111101",
			870 => "0000110000111000001100",
			871 => "0010111110111100000100",
			872 => "1111111000111100111101",
			873 => "0000101110101000000100",
			874 => "0000001000111100111101",
			875 => "0000000000111100111101",
			876 => "0010101100011100001100",
			877 => "0010000010101000001000",
			878 => "0000101101000100000100",
			879 => "0000000000111100111101",
			880 => "1111111000111100111101",
			881 => "0000000000111100111101",
			882 => "1111111000111100111101",
			883 => "0011100000001101000000",
			884 => "0001111100001000100000",
			885 => "0000111001110000010000",
			886 => "0001110111111000001000",
			887 => "0000100001000000000100",
			888 => "0000000000111100111101",
			889 => "1111111000111100111101",
			890 => "0000110111111000000100",
			891 => "0000001000111100111101",
			892 => "0000000000111100111101",
			893 => "0000100101110000001000",
			894 => "0011101100001000000100",
			895 => "0000000000111100111101",
			896 => "0000000000111100111101",
			897 => "0011001110111100000100",
			898 => "0000000000111100111101",
			899 => "0000000000111100111101",
			900 => "0001111100001000010000",
			901 => "0010101100011100001000",
			902 => "0011010000001100000100",
			903 => "0000001000111100111101",
			904 => "0000001000111100111101",
			905 => "0001000100001100000100",
			906 => "0000000000111100111101",
			907 => "0000001000111100111101",
			908 => "0001110100000000001000",
			909 => "0001010100001000000100",
			910 => "0000000000111100111101",
			911 => "0000001000111100111101",
			912 => "0011101000111000000100",
			913 => "0000001000111100111101",
			914 => "0000000000111100111101",
			915 => "0000100011001000011100",
			916 => "0001101010011000010000",
			917 => "0010101000010100001000",
			918 => "0001001000000100000100",
			919 => "0000000000111100111101",
			920 => "0000001000111100111101",
			921 => "0011000100000000000100",
			922 => "1111111000111100111101",
			923 => "0000000000111100111101",
			924 => "0000100101110000000100",
			925 => "0000010000111100111101",
			926 => "0010111101100000000100",
			927 => "0000000000111100111101",
			928 => "0000000000111100111101",
			929 => "0001101100011000001100",
			930 => "0000011100110100000100",
			931 => "1111111000111100111101",
			932 => "0010110101101100000100",
			933 => "0000010000111100111101",
			934 => "0000000000111100111101",
			935 => "0011001000111000001000",
			936 => "0001101001100100000100",
			937 => "0000000000111100111101",
			938 => "1111111000111100111101",
			939 => "0000011011101000000100",
			940 => "0000001000111100111101",
			941 => "1111111000111100111101",
			942 => "0010001001101000001100",
			943 => "0000011011101000001000",
			944 => "0000011011101000000100",
			945 => "1111111000111100111101",
			946 => "0000001000111100111101",
			947 => "1111111000111100111101",
			948 => "0001000010010000101000",
			949 => "0010000001110100011000",
			950 => "0011101011110000001100",
			951 => "0001001011100000001000",
			952 => "0001001000001000000100",
			953 => "0000000000111100111101",
			954 => "0000001000111100111101",
			955 => "1111111000111100111101",
			956 => "0001101001111100000100",
			957 => "1111111000111100111101",
			958 => "0001100100101100000100",
			959 => "0000000000111100111101",
			960 => "1111111000111100111101",
			961 => "0001001101110100001000",
			962 => "0001111111011100000100",
			963 => "0000001000111100111101",
			964 => "0000001000111100111101",
			965 => "0010001010101100000100",
			966 => "1111111000111100111101",
			967 => "0000001000111100111101",
			968 => "0001000000000000001100",
			969 => "0010000000110000000100",
			970 => "1111111000111100111101",
			971 => "0010100001110100000100",
			972 => "0000001000111100111101",
			973 => "1111111000111100111101",
			974 => "1111111000111100111101",
			975 => "0011011011000010011100",
			976 => "0001110111111001000000",
			977 => "0001111110111100101000",
			978 => "0011001010000000010000",
			979 => "0010110111111000001100",
			980 => "0001001011100000001000",
			981 => "0000000011111100000100",
			982 => "1111111001000100011001",
			983 => "0000001001000100011001",
			984 => "1111111001000100011001",
			985 => "1111111001000100011001",
			986 => "0001000011010100001000",
			987 => "0000100101001000000100",
			988 => "0000001001000100011001",
			989 => "0000000001000100011001",
			990 => "0010100110011100001000",
			991 => "0001011000111000000100",
			992 => "0000000001000100011001",
			993 => "1111111001000100011001",
			994 => "0000110010011000000100",
			995 => "1111111001000100011001",
			996 => "0000001001000100011001",
			997 => "0010101010110000010000",
			998 => "0001101011111100001000",
			999 => "0011110111010000000100",
			1000 => "0000001001000100011001",
			1001 => "0000000001000100011001",
			1002 => "0000011110100000000100",
			1003 => "1111110001000100011001",
			1004 => "1111111001000100011001",
			1005 => "0010000111000000000100",
			1006 => "0000001001000100011001",
			1007 => "1111111001000100011001",
			1008 => "0010101001000100111000",
			1009 => "0000101110000100011100",
			1010 => "0001010011011100001100",
			1011 => "0000111000111000001000",
			1012 => "0001110100010100000100",
			1013 => "1111111001000100011001",
			1014 => "0000000001000100011001",
			1015 => "1111110001000100011001",
			1016 => "0000111101100000001000",
			1017 => "0001010101101100000100",
			1018 => "0000000001000100011001",
			1019 => "0000001001000100011001",
			1020 => "0010000001110000000100",
			1021 => "0000000001000100011001",
			1022 => "0000000001000100011001",
			1023 => "0001001100001100010000",
			1024 => "0010101000010100001000",
			1025 => "0001001011110000000100",
			1026 => "0000000001000100011001",
			1027 => "0000001001000100011001",
			1028 => "0001000010010100000100",
			1029 => "0000010001000100011001",
			1030 => "0000000001000100011001",
			1031 => "0010000001110000000100",
			1032 => "1111111001000100011001",
			1033 => "0011111011011100000100",
			1034 => "0000000001000100011001",
			1035 => "0000001001000100011001",
			1036 => "0000001111000100000100",
			1037 => "0000010001000100011001",
			1038 => "0001000010110000010000",
			1039 => "0001110100010100001000",
			1040 => "0000100010011100000100",
			1041 => "0000000001000100011001",
			1042 => "0000010001000100011001",
			1043 => "0001011010111000000100",
			1044 => "0000000001000100011001",
			1045 => "0000001001000100011001",
			1046 => "0001111100001000001000",
			1047 => "0001111100001000000100",
			1048 => "0000000001000100011001",
			1049 => "0000000001000100011001",
			1050 => "0001111100001000000100",
			1051 => "0000000001000100011001",
			1052 => "0000000001000100011001",
			1053 => "0000000111000000011000",
			1054 => "0001011000000000010000",
			1055 => "0001111101100000001000",
			1056 => "0011011001001000000100",
			1057 => "0000000001000100011001",
			1058 => "0000000001000100011001",
			1059 => "0000001010100000000100",
			1060 => "0000000001000100011001",
			1061 => "0000001001000100011001",
			1062 => "0010000001110000000100",
			1063 => "1111111001000100011001",
			1064 => "0000000001000100011001",
			1065 => "0001000000000000111000",
			1066 => "0010111100101100011100",
			1067 => "0000110100000100001100",
			1068 => "0000011001111000000100",
			1069 => "1111111001000100011001",
			1070 => "0011110111100000000100",
			1071 => "0000000001000100011001",
			1072 => "0000001001000100011001",
			1073 => "0010100001010000001000",
			1074 => "0011111001010000000100",
			1075 => "1111111001000100011001",
			1076 => "0000001001000100011001",
			1077 => "0001101011001100000100",
			1078 => "1111110001000100011001",
			1079 => "1111111001000100011001",
			1080 => "0000110100000100001100",
			1081 => "0001011001001000001000",
			1082 => "0000111010001100000100",
			1083 => "0000000001000100011001",
			1084 => "1111111001000100011001",
			1085 => "1111111001000100011001",
			1086 => "0001100100111100001000",
			1087 => "0001111101100000000100",
			1088 => "0000000001000100011001",
			1089 => "0000000001000100011001",
			1090 => "0010001001101000000100",
			1091 => "1111111001000100011001",
			1092 => "0000000001000100011001",
			1093 => "1111111001000100011001",
			1094 => "0001000001001110111100",
			1095 => "0000111011000101010000",
			1096 => "0001100001111000100100",
			1097 => "0000100010110100010000",
			1098 => "0010111110111100000100",
			1099 => "1111111001001010111101",
			1100 => "0001001110000000000100",
			1101 => "0000000001001010111101",
			1102 => "0011001110111100000100",
			1103 => "0000000001001010111101",
			1104 => "0000001001001010111101",
			1105 => "0010000110001000001100",
			1106 => "0010110111111000001000",
			1107 => "0000110100010100000100",
			1108 => "0000000001001010111101",
			1109 => "1111110001001010111101",
			1110 => "1111110001001010111101",
			1111 => "0011000000111000000100",
			1112 => "0000000001001010111101",
			1113 => "0000001001001010111101",
			1114 => "0001000000010100011000",
			1115 => "0011110001101000010000",
			1116 => "0001101101111100001000",
			1117 => "0000100110100000000100",
			1118 => "0000001001001010111101",
			1119 => "0000000001001010111101",
			1120 => "0011101000110000000100",
			1121 => "0000001001001010111101",
			1122 => "0000000001001010111101",
			1123 => "0010000110001000000100",
			1124 => "0000000001001010111101",
			1125 => "0000001001001010111101",
			1126 => "0000000111111000001000",
			1127 => "0011101111000100000100",
			1128 => "0000000001001010111101",
			1129 => "1111110001001010111101",
			1130 => "0011110001011000001000",
			1131 => "0000100101110000000100",
			1132 => "0000000001001010111101",
			1133 => "1111111001001010111101",
			1134 => "0000001001001010111101",
			1135 => "0001010011011100101100",
			1136 => "0011100010011000001100",
			1137 => "0001011001110000001000",
			1138 => "0000111100001000000100",
			1139 => "0000000001001010111101",
			1140 => "1111111001001010111101",
			1141 => "1111101001001010111101",
			1142 => "0000011110100000010000",
			1143 => "0000010110000000001000",
			1144 => "0000001011000100000100",
			1145 => "1111111001001010111101",
			1146 => "0000000001001010111101",
			1147 => "0001100100110100000100",
			1148 => "0000000001001010111101",
			1149 => "1111111001001010111101",
			1150 => "0010110100010100001000",
			1151 => "0001110111111000000100",
			1152 => "0000000001001010111101",
			1153 => "1111110001001010111101",
			1154 => "0000111000111000000100",
			1155 => "0000001001001010111101",
			1156 => "1111111001001010111101",
			1157 => "0010111011000100100000",
			1158 => "0010110100010100010000",
			1159 => "0001000101010100001000",
			1160 => "0001100001111000000100",
			1161 => "0000001001001010111101",
			1162 => "1111111001001010111101",
			1163 => "0010110111111000000100",
			1164 => "0000001001001010111101",
			1165 => "0000000001001010111101",
			1166 => "0011001110111100001000",
			1167 => "0010100110011000000100",
			1168 => "0000001001001010111101",
			1169 => "1111111001001010111101",
			1170 => "0011110101110100000100",
			1171 => "0000000001001010111101",
			1172 => "0000001001001010111101",
			1173 => "0001110100010100010000",
			1174 => "0011111010010100001000",
			1175 => "0001011101100000000100",
			1176 => "0000000001001010111101",
			1177 => "1111111001001010111101",
			1178 => "0000100011001000000100",
			1179 => "0000010001001010111101",
			1180 => "0000000001001010111101",
			1181 => "0000111100001000001000",
			1182 => "0011111000011000000100",
			1183 => "1111111001001010111101",
			1184 => "0000000001001010111101",
			1185 => "0000110100000000000100",
			1186 => "0000001001001010111101",
			1187 => "0000000001001010111101",
			1188 => "0001111100001000010100",
			1189 => "0011000111111000001100",
			1190 => "0001011001110000000100",
			1191 => "1111111001001010111101",
			1192 => "0001010011011100000100",
			1193 => "0000000001001010111101",
			1194 => "1111111001001010111101",
			1195 => "0000101111010000000100",
			1196 => "0000000001001010111101",
			1197 => "0000001001001010111101",
			1198 => "1111111001001010111101",
			1199 => "0011000100000010010000",
			1200 => "0001111001110001100100",
			1201 => "0001011010111100110000",
			1202 => "0011000100000000010100",
			1203 => "0010011111001100010000",
			1204 => "0010010110101000001000",
			1205 => "0000110011011100000100",
			1206 => "0000000001010011010001",
			1207 => "0000000001010011010001",
			1208 => "0000011110100000000100",
			1209 => "0000001001010011010001",
			1210 => "0000000001010011010001",
			1211 => "0000001001010011010001",
			1212 => "0010111000111000010000",
			1213 => "0010101010110000001000",
			1214 => "0010001011010100000100",
			1215 => "0000000001010011010001",
			1216 => "0000001001010011010001",
			1217 => "0001000100001100000100",
			1218 => "1111111001010011010001",
			1219 => "0000001001010011010001",
			1220 => "0010000001110100001000",
			1221 => "0010101001000100000100",
			1222 => "0000000001010011010001",
			1223 => "0000001001010011010001",
			1224 => "0000000001010011010001",
			1225 => "0010011101011100100000",
			1226 => "0010111101100000010000",
			1227 => "0011000100000000001000",
			1228 => "0001110100000000000100",
			1229 => "1111111001010011010001",
			1230 => "0000000001010011010001",
			1231 => "0001111000111000000100",
			1232 => "0000001001010011010001",
			1233 => "1111111001010011010001",
			1234 => "0011111110101100001000",
			1235 => "0010011011101000000100",
			1236 => "1111111001010011010001",
			1237 => "0000001001010011010001",
			1238 => "0010111100110000000100",
			1239 => "1111111001010011010001",
			1240 => "0000000001010011010001",
			1241 => "0011000000101000000100",
			1242 => "0000001001010011010001",
			1243 => "0011101000000000001000",
			1244 => "0000100010000000000100",
			1245 => "0000000001010011010001",
			1246 => "0000001001010011010001",
			1247 => "0000101110110100000100",
			1248 => "1111111001010011010001",
			1249 => "0000000001010011010001",
			1250 => "0010000001110100100100",
			1251 => "0001011010111000001100",
			1252 => "0000100101110000000100",
			1253 => "0000000001010011010001",
			1254 => "0010000111000100000100",
			1255 => "0000001001010011010001",
			1256 => "0000001001010011010001",
			1257 => "0011010110100100001100",
			1258 => "0010101010110000001000",
			1259 => "0010111100101100000100",
			1260 => "0000001001010011010001",
			1261 => "1111111001010011010001",
			1262 => "1111111001010011010001",
			1263 => "0010011011111100001000",
			1264 => "0000101100010000000100",
			1265 => "0000000001010011010001",
			1266 => "0000001001010011010001",
			1267 => "0000000001010011010001",
			1268 => "0010000010101000000100",
			1269 => "1111111001010011010001",
			1270 => "0000000001010011010001",
			1271 => "0011000100000000100000",
			1272 => "0001011010111000011000",
			1273 => "0011010001111100001000",
			1274 => "0011111110101100000100",
			1275 => "1111111001010011010001",
			1276 => "0000000001010011010001",
			1277 => "0010101100011100001100",
			1278 => "0000011001111000001000",
			1279 => "0000100100101000000100",
			1280 => "0000000001010011010001",
			1281 => "1111111001010011010001",
			1282 => "0000000001010011010001",
			1283 => "0000000001010011010001",
			1284 => "0011101000011000000100",
			1285 => "0000001001010011010001",
			1286 => "1111111001010011010001",
			1287 => "0011001000111100100100",
			1288 => "0011001000111100010100",
			1289 => "0001111001110000001100",
			1290 => "0011110100010000000100",
			1291 => "0000001001010011010001",
			1292 => "0000101010001000000100",
			1293 => "1111111001010011010001",
			1294 => "0000000001010011010001",
			1295 => "0010000111000100000100",
			1296 => "1111111001010011010001",
			1297 => "0000000001010011010001",
			1298 => "0010001011010100001000",
			1299 => "0010100110011000000100",
			1300 => "0000001001010011010001",
			1301 => "1111111001010011010001",
			1302 => "0000101100000000000100",
			1303 => "0000001001010011010001",
			1304 => "0000000001010011010001",
			1305 => "0000010010001100011000",
			1306 => "0011110010001000001100",
			1307 => "0011111011011100001000",
			1308 => "0011111011011100000100",
			1309 => "0000000001010011010001",
			1310 => "0000000001010011010001",
			1311 => "1111111001010011010001",
			1312 => "0001011110110000001000",
			1313 => "0001111000111000000100",
			1314 => "0000001001010011010001",
			1315 => "0000001001010011010001",
			1316 => "0000000001010011010001",
			1317 => "0000011001111000010000",
			1318 => "0011001000111000001000",
			1319 => "0000010010001100000100",
			1320 => "0000000001010011010001",
			1321 => "1111111001010011010001",
			1322 => "0011100001111100000100",
			1323 => "0000000001010011010001",
			1324 => "0000001001010011010001",
			1325 => "0010100001010000001000",
			1326 => "0011100101100100000100",
			1327 => "1111111001010011010001",
			1328 => "0000000001010011010001",
			1329 => "0011011000000000000100",
			1330 => "0000001001010011010001",
			1331 => "0000000001010011010001",
			1332 => "0000001100001010110000",
			1333 => "0010101100011101010100",
			1334 => "0000100010110100101000",
			1335 => "0000100001001000010100",
			1336 => "0000001000110000001100",
			1337 => "0010111011000100000100",
			1338 => "1111111001011011110101",
			1339 => "0011000100010100000100",
			1340 => "0000000001011011110101",
			1341 => "1111111001011011110101",
			1342 => "0011001010000000000100",
			1343 => "0000000001011011110101",
			1344 => "0000001001011011110101",
			1345 => "0010000001110100010000",
			1346 => "0010101000010100001000",
			1347 => "0000101110101100000100",
			1348 => "0000000001011011110101",
			1349 => "1111111001011011110101",
			1350 => "0010101001000100000100",
			1351 => "0000001001011011110101",
			1352 => "0000000001011011110101",
			1353 => "1111111001011011110101",
			1354 => "0010000010101000100000",
			1355 => "0001000010100100010000",
			1356 => "0000111000111100001000",
			1357 => "0010110100010100000100",
			1358 => "0000000001011011110101",
			1359 => "0000000001011011110101",
			1360 => "0011011100101100000100",
			1361 => "0000000001011011110101",
			1362 => "0000000001011011110101",
			1363 => "0011010011011100001000",
			1364 => "0000001011000100000100",
			1365 => "0000000001011011110101",
			1366 => "0000001001011011110101",
			1367 => "0001100100110100000100",
			1368 => "1111111001011011110101",
			1369 => "0000000001011011110101",
			1370 => "0011010011011100000100",
			1371 => "0000000001011011110101",
			1372 => "0000111000111000000100",
			1373 => "0000001001011011110101",
			1374 => "0000001001011011110101",
			1375 => "0010010111100100101100",
			1376 => "0000110101101100011000",
			1377 => "0010010110101000010000",
			1378 => "0001000011110100001000",
			1379 => "0000001011000100000100",
			1380 => "1111111001011011110101",
			1381 => "0000000001011011110101",
			1382 => "0011000100010100000100",
			1383 => "0000001001011011110101",
			1384 => "0000000001011011110101",
			1385 => "0010010111100100000100",
			1386 => "0000001001011011110101",
			1387 => "0000000001011011110101",
			1388 => "0011100000101000001000",
			1389 => "0011101011000100000100",
			1390 => "0000000001011011110101",
			1391 => "1111110001011011110101",
			1392 => "0011100100000000000100",
			1393 => "0000001001011011110101",
			1394 => "0010100110011100000100",
			1395 => "1111111001011011110101",
			1396 => "0000000001011011110101",
			1397 => "0001101101011000011000",
			1398 => "0000110001111100001100",
			1399 => "0011101100110000001000",
			1400 => "0011000000101000000100",
			1401 => "0000001001011011110101",
			1402 => "0000000001011011110101",
			1403 => "1111111001011011110101",
			1404 => "0011111101000100000100",
			1405 => "0000001001011011110101",
			1406 => "0011010001111100000100",
			1407 => "0000001001011011110101",
			1408 => "0000000001011011110101",
			1409 => "0001111000111000001100",
			1410 => "0000111010111100000100",
			1411 => "0000000001011011110101",
			1412 => "0011011010111100000100",
			1413 => "1111111001011011110101",
			1414 => "0000000001011011110101",
			1415 => "0011010111001000000100",
			1416 => "0000001001011011110101",
			1417 => "0001000010100100000100",
			1418 => "0000000001011011110101",
			1419 => "0000000001011011110101",
			1420 => "0011000111111000101100",
			1421 => "0000110100000000101000",
			1422 => "0000110100010100011100",
			1423 => "0010100110011100001100",
			1424 => "0011000000111000000100",
			1425 => "0000000001011011110101",
			1426 => "0001101101111100000100",
			1427 => "0000000001011011110101",
			1428 => "0000001001011011110101",
			1429 => "0011011000111100001000",
			1430 => "0011001010000000000100",
			1431 => "0000000001011011110101",
			1432 => "1111111001011011110101",
			1433 => "0000110000111000000100",
			1434 => "0000001001011011110101",
			1435 => "0000000001011011110101",
			1436 => "0000000100000000000100",
			1437 => "0000000001011011110101",
			1438 => "0011011000111000000100",
			1439 => "0000000001011011110101",
			1440 => "1111111001011011110101",
			1441 => "0000001001011011110101",
			1442 => "0001110100010100010000",
			1443 => "0010011100110100001100",
			1444 => "0011110100011000001000",
			1445 => "0010010000011000000100",
			1446 => "0000000001011011110101",
			1447 => "0000001001011011110101",
			1448 => "1111111001011011110101",
			1449 => "0000001001011011110101",
			1450 => "0010110000101000010100",
			1451 => "0010010110101000001100",
			1452 => "0001000011011000000100",
			1453 => "0000001001011011110101",
			1454 => "0001100100110100000100",
			1455 => "0000001001011011110101",
			1456 => "0000000001011011110101",
			1457 => "0000100011001000000100",
			1458 => "1111111001011011110101",
			1459 => "0000000001011011110101",
			1460 => "0011011110001100000100",
			1461 => "0000001001011011110101",
			1462 => "0010010110101000001000",
			1463 => "0001101101111100000100",
			1464 => "0000000001011011110101",
			1465 => "1111111001011011110101",
			1466 => "0010000111000000000100",
			1467 => "0000000001011011110101",
			1468 => "0000001001011011110101",
			1469 => "0011100101101110011000",
			1470 => "0011110101100101011100",
			1471 => "0001100111101000101000",
			1472 => "0011010110000100011000",
			1473 => "0000111000111000010000",
			1474 => "0000000011111100001000",
			1475 => "0010000101000100000100",
			1476 => "1111111001100101010001",
			1477 => "0000001001100101010001",
			1478 => "0001110100010100000100",
			1479 => "0000000001100101010001",
			1480 => "0000001001100101010001",
			1481 => "0011101110111100000100",
			1482 => "1111111001100101010001",
			1483 => "1111111001100101010001",
			1484 => "0001010101101100000100",
			1485 => "0000000001100101010001",
			1486 => "0000001001101000000100",
			1487 => "0000000001100101010001",
			1488 => "0010001100000100000100",
			1489 => "0000001001100101010001",
			1490 => "0000000001100101010001",
			1491 => "0000111100110000100000",
			1492 => "0010111100001000010000",
			1493 => "0001011101100000001000",
			1494 => "0010110100010100000100",
			1495 => "0000000001100101010001",
			1496 => "0000000001100101010001",
			1497 => "0001011101100000000100",
			1498 => "1111111001100101010001",
			1499 => "0000000001100101010001",
			1500 => "0011110100000100001000",
			1501 => "0000000011010000000100",
			1502 => "1111111001100101010001",
			1503 => "0000000001100101010001",
			1504 => "0000011110100000000100",
			1505 => "0000000001100101010001",
			1506 => "0000001001100101010001",
			1507 => "0000101111010000010000",
			1508 => "0000100111100000001000",
			1509 => "0000101101000100000100",
			1510 => "1111111001100101010001",
			1511 => "0000000001100101010001",
			1512 => "0001011110001100000100",
			1513 => "1111111001100101010001",
			1514 => "1111111001100101010001",
			1515 => "0000000001100101010001",
			1516 => "0010000111000000101100",
			1517 => "0001000011011000011100",
			1518 => "0011010011011100001100",
			1519 => "0001001001001100000100",
			1520 => "1111110001100101010001",
			1521 => "0001000011010100000100",
			1522 => "0000001001100101010001",
			1523 => "1111111001100101010001",
			1524 => "0000111001110000001000",
			1525 => "0000000000101000000100",
			1526 => "0000000001100101010001",
			1527 => "0000000001100101010001",
			1528 => "0000000000110000000100",
			1529 => "0000000001100101010001",
			1530 => "0000000001100101010001",
			1531 => "0011111010010100001000",
			1532 => "0001110111111000000100",
			1533 => "0000000001100101010001",
			1534 => "1111110001100101010001",
			1535 => "0010000001110100000100",
			1536 => "0000000001100101010001",
			1537 => "0000001001100101010001",
			1538 => "0001000001001100001000",
			1539 => "0000100010000100000100",
			1540 => "0000001001100101010001",
			1541 => "0000000001100101010001",
			1542 => "0001011101111000000100",
			1543 => "0000000001100101010001",
			1544 => "1111111001100101010001",
			1545 => "0000110111001001001000",
			1546 => "0011000000101000100000",
			1547 => "0011000100010100010000",
			1548 => "0011111110101000001100",
			1549 => "0001001100111000000100",
			1550 => "0000011001100101010001",
			1551 => "0011111101000100000100",
			1552 => "0000000001100101010001",
			1553 => "1111111001100101010001",
			1554 => "0000001001100101010001",
			1555 => "0011000100010100001000",
			1556 => "0001001100001100000100",
			1557 => "0000000001100101010001",
			1558 => "1111111001100101010001",
			1559 => "0011111110101100000100",
			1560 => "1111111001100101010001",
			1561 => "0000000001100101010001",
			1562 => "0010111000111100010100",
			1563 => "0010001001101000000100",
			1564 => "1111111001100101010001",
			1565 => "0011101100101100001000",
			1566 => "0010000110001000000100",
			1567 => "0000001001100101010001",
			1568 => "0000000001100101010001",
			1569 => "0011000000101000000100",
			1570 => "0000000001100101010001",
			1571 => "0000001001100101010001",
			1572 => "0000101100100100001000",
			1573 => "0001101101011100000100",
			1574 => "0000000001100101010001",
			1575 => "0000010001100101010001",
			1576 => "0011000000101000000100",
			1577 => "0000000001100101010001",
			1578 => "0011100000001100000100",
			1579 => "0000000001100101010001",
			1580 => "1111111001100101010001",
			1581 => "0000110111001000010100",
			1582 => "0000001010000000001100",
			1583 => "0011010001111100000100",
			1584 => "0000010001100101010001",
			1585 => "0001000010110000000100",
			1586 => "0000000001100101010001",
			1587 => "0000001001100101010001",
			1588 => "0011110010110100000100",
			1589 => "1111111001100101010001",
			1590 => "0000001001100101010001",
			1591 => "0001101010011000100000",
			1592 => "0000100010000100010000",
			1593 => "0001001110111000001000",
			1594 => "0001100100110100000100",
			1595 => "0000000001100101010001",
			1596 => "0000000001100101010001",
			1597 => "0001000011010100000100",
			1598 => "0000001001100101010001",
			1599 => "0000000001100101010001",
			1600 => "0001110100000000001000",
			1601 => "0011010100001000000100",
			1602 => "0000000001100101010001",
			1603 => "0000001001100101010001",
			1604 => "0001101010011000000100",
			1605 => "0000000001100101010001",
			1606 => "0000001001100101010001",
			1607 => "0001010100001000001100",
			1608 => "0000100110111100001000",
			1609 => "0011101010111100000100",
			1610 => "1111111001100101010001",
			1611 => "0000000001100101010001",
			1612 => "0000000001100101010001",
			1613 => "0011110001000000001000",
			1614 => "0000100010000100000100",
			1615 => "0000000001100101010001",
			1616 => "0000001001100101010001",
			1617 => "0011100100000100000100",
			1618 => "0000000001100101010001",
			1619 => "0000000001100101010001",
			1620 => "0011011011000010111100",
			1621 => "0011110101100101000100",
			1622 => "0011100100000000110100",
			1623 => "0001000110110000100000",
			1624 => "0000110000110000010000",
			1625 => "0001110111111000001000",
			1626 => "0000110011111100000100",
			1627 => "0000001001101101010101",
			1628 => "0000000001101101010101",
			1629 => "0011111010111000000100",
			1630 => "0000000001101101010101",
			1631 => "0000001001101101010101",
			1632 => "0001111100001000001000",
			1633 => "0011000100010100000100",
			1634 => "0000000001101101010101",
			1635 => "0000000001101101010101",
			1636 => "0001111100001000000100",
			1637 => "0000001001101101010101",
			1638 => "0000000001101101010101",
			1639 => "0001101010011000001100",
			1640 => "0001000011111000000100",
			1641 => "1111111001101101010101",
			1642 => "0001000101100000000100",
			1643 => "0000000001101101010101",
			1644 => "1111111001101101010101",
			1645 => "0010101000110000000100",
			1646 => "0000001001101101010101",
			1647 => "0000000001101101010101",
			1648 => "0001100111101000001000",
			1649 => "0000100001001000000100",
			1650 => "1111111001101101010101",
			1651 => "0000001001101101010101",
			1652 => "0011000100010100000100",
			1653 => "0000000001101101010101",
			1654 => "1111111001101101010101",
			1655 => "0010100110011000111100",
			1656 => "0000100100101000100000",
			1657 => "0000110110000100010000",
			1658 => "0010010110101000001000",
			1659 => "0000111101100000000100",
			1660 => "0000000001101101010101",
			1661 => "1111111001101101010101",
			1662 => "0011000111111000000100",
			1663 => "0000010001101101010101",
			1664 => "0000001001101101010101",
			1665 => "0010010110101000001000",
			1666 => "0011110101110100000100",
			1667 => "1111111001101101010101",
			1668 => "0000000001101101010101",
			1669 => "0010101000010100000100",
			1670 => "0000000001101101010101",
			1671 => "0000000001101101010101",
			1672 => "0000100100101000001100",
			1673 => "0000110100001000001000",
			1674 => "0001001000001000000100",
			1675 => "0000010001101101010101",
			1676 => "0000001001101101010101",
			1677 => "0000000001101101010101",
			1678 => "0001100001111000001000",
			1679 => "0011101001110000000100",
			1680 => "0000000001101101010101",
			1681 => "1111111001101101010101",
			1682 => "0011001000111100000100",
			1683 => "0000000001101101010101",
			1684 => "1111111001101101010101",
			1685 => "0011100100010100011100",
			1686 => "0011001110111100010000",
			1687 => "0001100100110100001000",
			1688 => "0011110110110100000100",
			1689 => "0000000001101101010101",
			1690 => "1111111001101101010101",
			1691 => "0000100011001000000100",
			1692 => "0000001001101101010101",
			1693 => "0000000001101101010101",
			1694 => "0000000000111000000100",
			1695 => "0000000001101101010101",
			1696 => "0010100001010000000100",
			1697 => "0000001001101101010101",
			1698 => "0000000001101101010101",
			1699 => "0010010110101000010000",
			1700 => "0011110111110000001000",
			1701 => "0000111101100000000100",
			1702 => "0000000001101101010101",
			1703 => "1111111001101101010101",
			1704 => "0010100001010000000100",
			1705 => "0000001001101101010101",
			1706 => "0000000001101101010101",
			1707 => "0011101100001000001000",
			1708 => "0001100100110100000100",
			1709 => "0000001001101101010101",
			1710 => "0000000001101101010101",
			1711 => "0001000011010100000100",
			1712 => "0000000001101101010101",
			1713 => "0000000001101101010101",
			1714 => "0000000111000000010100",
			1715 => "0010110000001100010000",
			1716 => "0010001100011100001100",
			1717 => "0001110101101100000100",
			1718 => "1111111001101101010101",
			1719 => "0001110101101100000100",
			1720 => "0000000001101101010101",
			1721 => "0000000001101101010101",
			1722 => "0000000001101101010101",
			1723 => "1111111001101101010101",
			1724 => "0001000000000000110000",
			1725 => "0010011101011100010100",
			1726 => "0011001000111000001100",
			1727 => "0011011000000000000100",
			1728 => "0000000001101101010101",
			1729 => "0001111101100000000100",
			1730 => "1111111001101101010101",
			1731 => "1111111001101101010101",
			1732 => "0001101101011000000100",
			1733 => "0000000001101101010101",
			1734 => "0000001001101101010101",
			1735 => "0001111101100000001100",
			1736 => "0011100001101000000100",
			1737 => "0000001001101101010101",
			1738 => "0001000011110000000100",
			1739 => "1111111001101101010101",
			1740 => "0000000001101101010101",
			1741 => "0011100011100000001000",
			1742 => "0010101010110000000100",
			1743 => "1111111001101101010101",
			1744 => "0000000001101101010101",
			1745 => "0011011001001000000100",
			1746 => "0000001001101101010101",
			1747 => "0000000001101101010101",
			1748 => "1111111001101101010101",
			1749 => "0011000111111010001000",
			1750 => "0010010110101001001100",
			1751 => "0000111001110000110000",
			1752 => "0001111011000100100000",
			1753 => "0000000010111100010000",
			1754 => "0001010011011100001000",
			1755 => "0001000101000000000100",
			1756 => "1111111001110110110001",
			1757 => "1111101001110110110001",
			1758 => "0011000111111000000100",
			1759 => "0000001001110110110001",
			1760 => "0000000001110110110001",
			1761 => "0000010110000000001000",
			1762 => "0000110011010000000100",
			1763 => "0000000001110110110001",
			1764 => "0000000001110110110001",
			1765 => "0000111011000100000100",
			1766 => "0000000001110110110001",
			1767 => "0000000001110110110001",
			1768 => "0011000111111000000100",
			1769 => "0000001001110110110001",
			1770 => "0001101101111100001000",
			1771 => "0001100001111000000100",
			1772 => "0000001001110110110001",
			1773 => "0000000001110110110001",
			1774 => "0000001001110110110001",
			1775 => "0010000010101000011000",
			1776 => "0011100111111000001100",
			1777 => "0011000111111000001000",
			1778 => "0000100011001000000100",
			1779 => "0000000001110110110001",
			1780 => "1111111001110110110001",
			1781 => "1111111001110110110001",
			1782 => "0001001111100000001000",
			1783 => "0000000011010000000100",
			1784 => "1111111001110110110001",
			1785 => "0000000001110110110001",
			1786 => "1111111001110110110001",
			1787 => "0000001001110110110001",
			1788 => "0001011100110000010100",
			1789 => "0010110000101000010000",
			1790 => "0011101000111100001100",
			1791 => "0011101110111100000100",
			1792 => "0000000001110110110001",
			1793 => "0001101101111100000100",
			1794 => "0000001001110110110001",
			1795 => "0000001001110110110001",
			1796 => "0000000001110110110001",
			1797 => "0000010001110110110001",
			1798 => "0011001110111100010000",
			1799 => "0010101001000100000100",
			1800 => "0000001001110110110001",
			1801 => "0011001010000000000100",
			1802 => "0000000001110110110001",
			1803 => "0000110110000100000100",
			1804 => "1111111001110110110001",
			1805 => "1111111001110110110001",
			1806 => "0001111100001000010000",
			1807 => "0011101001110000001000",
			1808 => "0010010111100100000100",
			1809 => "0000000001110110110001",
			1810 => "0000001001110110110001",
			1811 => "0000110100001000000100",
			1812 => "0000000001110110110001",
			1813 => "0000001001110110110001",
			1814 => "0001011110001100000100",
			1815 => "1111111001110110110001",
			1816 => "0000000001110110110001",
			1817 => "0011000100010100110100",
			1818 => "0010101001000100010100",
			1819 => "0001110100010100000100",
			1820 => "1111111001110110110001",
			1821 => "0000011110100000001000",
			1822 => "0001100001111000000100",
			1823 => "0000000001110110110001",
			1824 => "0000001001110110110001",
			1825 => "0011000111111000000100",
			1826 => "0000000001110110110001",
			1827 => "1111111001110110110001",
			1828 => "0000100011001000011000",
			1829 => "0001110100010100001100",
			1830 => "0010111110111100000100",
			1831 => "0000001001110110110001",
			1832 => "0000110000110000000100",
			1833 => "1111111001110110110001",
			1834 => "0000000001110110110001",
			1835 => "0000010110000000000100",
			1836 => "0000001001110110110001",
			1837 => "0011100100010100000100",
			1838 => "1111111001110110110001",
			1839 => "1111111001110110110001",
			1840 => "0001101100011000000100",
			1841 => "0000001001110110110001",
			1842 => "1111111001110110110001",
			1843 => "0000111100110000111000",
			1844 => "0010010110101000011100",
			1845 => "0000011110100000010000",
			1846 => "0001010101101100001000",
			1847 => "0000110011011100000100",
			1848 => "0000000001110110110001",
			1849 => "1111111001110110110001",
			1850 => "0000100111100000000100",
			1851 => "0000000001110110110001",
			1852 => "0000000001110110110001",
			1853 => "0001101100011000001000",
			1854 => "0001111100001000000100",
			1855 => "0000000001110110110001",
			1856 => "1111111001110110110001",
			1857 => "0000001001110110110001",
			1858 => "0010001011010100001100",
			1859 => "0001001100001100001000",
			1860 => "0000100110100000000100",
			1861 => "0000000001110110110001",
			1862 => "0000001001110110110001",
			1863 => "1111111001110110110001",
			1864 => "0001001110111000001000",
			1865 => "0001000010111000000100",
			1866 => "0000001001110110110001",
			1867 => "0000001001110110110001",
			1868 => "0001101010011000000100",
			1869 => "0000000001110110110001",
			1870 => "0000001001110110110001",
			1871 => "0010010111100100011100",
			1872 => "0000111101111000010000",
			1873 => "0000101100010100001000",
			1874 => "0000111100110000000100",
			1875 => "1111111001110110110001",
			1876 => "0000000001110110110001",
			1877 => "0010100110011100000100",
			1878 => "0000001001110110110001",
			1879 => "0000000001110110110001",
			1880 => "0001001011100000001000",
			1881 => "0010101100011100000100",
			1882 => "1111111001110110110001",
			1883 => "1111110001110110110001",
			1884 => "0000001001110110110001",
			1885 => "0000011100110100010000",
			1886 => "0000110000001100001000",
			1887 => "0000101001010000000100",
			1888 => "0000000001110110110001",
			1889 => "0000001001110110110001",
			1890 => "0010111100001000000100",
			1891 => "0000001001110110110001",
			1892 => "0000000001110110110001",
			1893 => "0010010111100100001000",
			1894 => "0010000111000100000100",
			1895 => "0000000001110110110001",
			1896 => "0000000001110110110001",
			1897 => "0010110100000000000100",
			1898 => "0000001001110110110001",
			1899 => "0000000001110110110001",
			1900 => "0011100101101110100000",
			1901 => "0011110101100101011100",
			1902 => "0001100111101000101000",
			1903 => "0011010110000100011000",
			1904 => "0000111000111000010000",
			1905 => "0001011000111000001000",
			1906 => "0011111011000000000100",
			1907 => "0000000010000000010101",
			1908 => "1111110010000000010101",
			1909 => "0010101001000100000100",
			1910 => "0000000010000000010101",
			1911 => "1111111010000000010101",
			1912 => "0000001101010000000100",
			1913 => "1111110010000000010101",
			1914 => "1111111010000000010101",
			1915 => "0001010101101100000100",
			1916 => "0000000010000000010101",
			1917 => "0000001001101000000100",
			1918 => "0000000010000000010101",
			1919 => "0011110000011100000100",
			1920 => "0000001010000000010101",
			1921 => "0000000010000000010101",
			1922 => "0000111100110000100000",
			1923 => "0010111100001000010000",
			1924 => "0001011101100000001000",
			1925 => "0001010011011100000100",
			1926 => "0000000010000000010101",
			1927 => "0000001010000000010101",
			1928 => "0011101011000100000100",
			1929 => "0000000010000000010101",
			1930 => "0000001010000000010101",
			1931 => "0011110111010000001000",
			1932 => "0000111001110000000100",
			1933 => "0000000010000000010101",
			1934 => "1111111010000000010101",
			1935 => "0000111001110000000100",
			1936 => "0000001010000000010101",
			1937 => "0000000010000000010101",
			1938 => "0011011101010100010000",
			1939 => "0000011100110100001000",
			1940 => "0011011100101000000100",
			1941 => "1111111010000000010101",
			1942 => "0000000010000000010101",
			1943 => "0000010010001100000100",
			1944 => "1111111010000000010101",
			1945 => "1111111010000000010101",
			1946 => "0000000010000000010101",
			1947 => "0010011011101000101100",
			1948 => "0010111101100000100000",
			1949 => "0000111001110000010000",
			1950 => "0011010011011100001000",
			1951 => "0011110101110100000100",
			1952 => "1111111010000000010101",
			1953 => "0000001010000000010101",
			1954 => "0000000000101000000100",
			1955 => "0000001010000000010101",
			1956 => "0000000010000000010101",
			1957 => "0010011001111000001000",
			1958 => "0010110000101000000100",
			1959 => "1111111010000000010101",
			1960 => "0000001010000000010101",
			1961 => "0010010110101000000100",
			1962 => "0000000010000000010101",
			1963 => "0000000010000000010101",
			1964 => "0001111001110000000100",
			1965 => "1111110010000000010101",
			1966 => "0001010000011100000100",
			1967 => "0000001010000000010101",
			1968 => "0000000010000000010101",
			1969 => "0001101010011000001000",
			1970 => "0011101100110000000100",
			1971 => "0000001010000000010101",
			1972 => "0000001010000000010101",
			1973 => "0011110000110100001000",
			1974 => "0000111010111100000100",
			1975 => "0000001010000000010101",
			1976 => "0000000010000000010101",
			1977 => "0000101011101100000100",
			1978 => "1111110010000000010101",
			1979 => "0000000010000000010101",
			1980 => "0000001111000100111000",
			1981 => "0010010100110100110000",
			1982 => "0001001000000100011100",
			1983 => "0000001101010000001100",
			1984 => "0001001011110000001000",
			1985 => "0001101010011000000100",
			1986 => "0000000010000000010101",
			1987 => "0000001010000000010101",
			1988 => "0000001010000000010101",
			1989 => "0010101001000100001000",
			1990 => "0001011100101000000100",
			1991 => "0000000010000000010101",
			1992 => "1111111010000000010101",
			1993 => "0001101001100100000100",
			1994 => "0000001010000000010101",
			1995 => "0000000010000000010101",
			1996 => "0001101101111100000100",
			1997 => "1111111010000000010101",
			1998 => "0000101100010100001000",
			1999 => "0000100100101000000100",
			2000 => "0000001010000000010101",
			2001 => "0000010010000000010101",
			2002 => "0011100101100100000100",
			2003 => "0000000010000000010101",
			2004 => "0000001010000000010101",
			2005 => "0010101010110000000100",
			2006 => "1111111010000000010101",
			2007 => "0000000010000000010101",
			2008 => "0000101110010000100000",
			2009 => "0000110000001100000100",
			2010 => "0000001010000000010101",
			2011 => "0001101010011000010000",
			2012 => "0011010001111100001000",
			2013 => "0011011100101000000100",
			2014 => "1111111010000000010101",
			2015 => "0000000010000000010101",
			2016 => "0010100001010000000100",
			2017 => "1111111010000000010101",
			2018 => "0000000010000000010101",
			2019 => "0010011101101000000100",
			2020 => "0000001010000000010101",
			2021 => "0010011011101000000100",
			2022 => "1111111010000000010101",
			2023 => "0000000010000000010101",
			2024 => "0001101100011000011100",
			2025 => "0011110010110100001100",
			2026 => "0010111000111100000100",
			2027 => "1111111010000000010101",
			2028 => "0011111110101100000100",
			2029 => "0000001010000000010101",
			2030 => "0000000010000000010101",
			2031 => "0011101110001100001000",
			2032 => "0010100001010000000100",
			2033 => "0000001010000000010101",
			2034 => "0000000010000000010101",
			2035 => "0000100110010000000100",
			2036 => "0000000010000000010101",
			2037 => "0000001010000000010101",
			2038 => "0010011011101000010000",
			2039 => "0011111110101100001000",
			2040 => "0001001010110100000100",
			2041 => "0000000010000000010101",
			2042 => "0000001010000000010101",
			2043 => "0001010111001000000100",
			2044 => "0000000010000000010101",
			2045 => "0000001010000000010101",
			2046 => "0000111011000000001000",
			2047 => "0000101100010100000100",
			2048 => "0000000010000000010101",
			2049 => "0000001010000000010101",
			2050 => "0001000101000000000100",
			2051 => "1111111010000000010101",
			2052 => "0000000010000000010101",
			2053 => "0010001001101010110000",
			2054 => "0010001001101001011100",
			2055 => "0011010101101100101000",
			2056 => "0001110100010100011000",
			2057 => "0000111000111000010000",
			2058 => "0000000011111100001000",
			2059 => "0010110100010100000100",
			2060 => "0000000010001010011001",
			2061 => "0000001010001010011001",
			2062 => "0011110000011100000100",
			2063 => "1111111010001010011001",
			2064 => "0000001010001010011001",
			2065 => "0000000011111100000100",
			2066 => "1111111010001010011001",
			2067 => "0000000010001010011001",
			2068 => "0000101101000100001100",
			2069 => "0000110100010100000100",
			2070 => "0000000010001010011001",
			2071 => "0011011100110000000100",
			2072 => "1111110010001010011001",
			2073 => "1111111010001010011001",
			2074 => "0000000010001010011001",
			2075 => "0000010010001100011100",
			2076 => "0010111001110000010000",
			2077 => "0001110100010100001000",
			2078 => "0000011110100000000100",
			2079 => "0000000010001010011001",
			2080 => "1111111010001010011001",
			2081 => "0010110000101000000100",
			2082 => "0000001010001010011001",
			2083 => "0000000010001010011001",
			2084 => "0000101110101000000100",
			2085 => "1111111010001010011001",
			2086 => "0001001110100100000100",
			2087 => "0000001010001010011001",
			2088 => "0000000010001010011001",
			2089 => "0011010001111100001000",
			2090 => "0001010000001100000100",
			2091 => "0000000010001010011001",
			2092 => "1111111010001010011001",
			2093 => "0001000110001100001000",
			2094 => "0000001111000100000100",
			2095 => "0000000010001010011001",
			2096 => "1111111010001010011001",
			2097 => "0011000110000100000100",
			2098 => "0000001010001010011001",
			2099 => "1111111010001010011001",
			2100 => "0000100101110000110000",
			2101 => "0000011100110100100000",
			2102 => "0011110100000100010000",
			2103 => "0011111111011100001000",
			2104 => "0001011100110000000100",
			2105 => "0000001010001010011001",
			2106 => "0000000010001010011001",
			2107 => "0001011101100000000100",
			2108 => "0000000010001010011001",
			2109 => "1111111010001010011001",
			2110 => "0000111101100000001000",
			2111 => "0001100001111000000100",
			2112 => "0000000010001010011001",
			2113 => "0000001010001010011001",
			2114 => "0001111100001000000100",
			2115 => "0000000010001010011001",
			2116 => "0000001010001010011001",
			2117 => "0010011101101000001100",
			2118 => "0010001001101000000100",
			2119 => "0000000010001010011001",
			2120 => "0000111110001100000100",
			2121 => "1111110010001010011001",
			2122 => "1111111010001010011001",
			2123 => "0000001010001010011001",
			2124 => "0000011001111000010100",
			2125 => "0000111011000000010000",
			2126 => "0000010010001100001000",
			2127 => "0011011100101000000100",
			2128 => "0000000010001010011001",
			2129 => "0000001010001010011001",
			2130 => "0000010010001100000100",
			2131 => "1111111010001010011001",
			2132 => "0000000010001010011001",
			2133 => "0000010010001010011001",
			2134 => "0001101010011000000100",
			2135 => "1111111010001010011001",
			2136 => "0011000100000000000100",
			2137 => "0000001010001010011001",
			2138 => "0001111001110000000100",
			2139 => "0000000010001010011001",
			2140 => "0000000010001010011001",
			2141 => "0000100111111101001000",
			2142 => "0010001011010100010100",
			2143 => "0011111010010100010000",
			2144 => "0011001010000000000100",
			2145 => "1111111010001010011001",
			2146 => "0000000011111100000100",
			2147 => "1111111010001010011001",
			2148 => "0010001001101000000100",
			2149 => "1111111010001010011001",
			2150 => "0000000010001010011001",
			2151 => "0000000010001010011001",
			2152 => "0010001011010100010100",
			2153 => "0011000100010100001100",
			2154 => "0000100001000000000100",
			2155 => "0000000010001010011001",
			2156 => "0000111101100000000100",
			2157 => "0000001010001010011001",
			2158 => "0000001010001010011001",
			2159 => "0011011101111000000100",
			2160 => "1111111010001010011001",
			2161 => "0000001010001010011001",
			2162 => "0000111101111000010000",
			2163 => "0011010000001100001000",
			2164 => "0001110100010100000100",
			2165 => "0000000010001010011001",
			2166 => "0000000010001010011001",
			2167 => "0011000000101000000100",
			2168 => "0000000010001010011001",
			2169 => "0000001010001010011001",
			2170 => "0010011011101000001000",
			2171 => "0010001011010100000100",
			2172 => "0000000010001010011001",
			2173 => "1111111010001010011001",
			2174 => "0000010010001100000100",
			2175 => "0000001010001010011001",
			2176 => "0000000010001010011001",
			2177 => "0000100111111100001100",
			2178 => "0001101100011000001000",
			2179 => "0010111000111100000100",
			2180 => "0000001010001010011001",
			2181 => "0000000010001010011001",
			2182 => "1111111010001010011001",
			2183 => "0001000100001100100000",
			2184 => "0010000001110100010000",
			2185 => "0001110100000000001000",
			2186 => "0001110100000000000100",
			2187 => "0000000010001010011001",
			2188 => "0000000010001010011001",
			2189 => "0001010001111100000100",
			2190 => "0000000010001010011001",
			2191 => "0000000010001010011001",
			2192 => "0010011101101000001000",
			2193 => "0010010110101000000100",
			2194 => "0000001010001010011001",
			2195 => "1111111010001010011001",
			2196 => "0011110110100000000100",
			2197 => "0000001010001010011001",
			2198 => "0000000010001010011001",
			2199 => "0010001111001000010000",
			2200 => "0010111000111100001000",
			2201 => "0000001110111100000100",
			2202 => "1111001010001010011001",
			2203 => "0000000010001010011001",
			2204 => "0010000110001000000100",
			2205 => "1111111010001010011001",
			2206 => "0000000010001010011001",
			2207 => "0011000111111000001000",
			2208 => "0011001010000000000100",
			2209 => "0000000010001010011001",
			2210 => "1111111010001010011001",
			2211 => "0010000010101000000100",
			2212 => "0000000010001010011001",
			2213 => "0000000010001010011001",
			2214 => "0000100110010010110000",
			2215 => "0011000100000001100100",
			2216 => "0010111000111100110000",
			2217 => "0011010000001100010100",
			2218 => "0010011101101000010000",
			2219 => "0011011101111000001000",
			2220 => "0011000000101000000100",
			2221 => "0000000010010101000101",
			2222 => "0000000010010101000101",
			2223 => "0011000111111000000100",
			2224 => "0000001010010101000101",
			2225 => "0000000010010101000101",
			2226 => "0000001010010101000101",
			2227 => "0001011101111000001100",
			2228 => "0010010111100100000100",
			2229 => "0000000010010101000101",
			2230 => "0001000011110000000100",
			2231 => "0000000010010101000101",
			2232 => "0000001010010101000101",
			2233 => "0010110100000000001000",
			2234 => "0011011100101000000100",
			2235 => "1111111010010101000101",
			2236 => "0000000010010101000101",
			2237 => "0011101101100000000100",
			2238 => "0000000010010101000101",
			2239 => "0000000010010101000101",
			2240 => "0011000000101000010100",
			2241 => "0001100001111000001000",
			2242 => "0001001011110000000100",
			2243 => "0000000010010101000101",
			2244 => "0000001010010101000101",
			2245 => "0001000100001100001000",
			2246 => "0000001110111100000100",
			2247 => "1111111010010101000101",
			2248 => "0000000010010101000101",
			2249 => "1111110010010101000101",
			2250 => "0011000000101000010000",
			2251 => "0000101001011100001000",
			2252 => "0011101000111000000100",
			2253 => "0000001010010101000101",
			2254 => "0000000010010101000101",
			2255 => "0010100001010000000100",
			2256 => "0000001010010101000101",
			2257 => "0000000010010101000101",
			2258 => "0001101101011000001000",
			2259 => "0011000000101000000100",
			2260 => "0000000010010101000101",
			2261 => "0000000010010101000101",
			2262 => "0001101101011000000100",
			2263 => "0000001010010101000101",
			2264 => "0000000010010101000101",
			2265 => "0011000100000000100000",
			2266 => "0010101010110000010000",
			2267 => "0000101100010100001100",
			2268 => "0001101100011000001000",
			2269 => "0000011100110100000100",
			2270 => "0000001010010101000101",
			2271 => "0000000010010101000101",
			2272 => "0000010010010101000101",
			2273 => "0000000010010101000101",
			2274 => "0010101100011100001000",
			2275 => "0011101100101100000100",
			2276 => "1111111010010101000101",
			2277 => "0000000010010101000101",
			2278 => "0001110100000000000100",
			2279 => "0000000010010101000101",
			2280 => "0000001010010101000101",
			2281 => "0001101100011000011100",
			2282 => "0001100100110100001100",
			2283 => "0001010000001100000100",
			2284 => "1111111010010101000101",
			2285 => "0001000000010000000100",
			2286 => "0000000010010101000101",
			2287 => "0000001010010101000101",
			2288 => "0001001001001100001000",
			2289 => "0001011010111100000100",
			2290 => "0000000010010101000101",
			2291 => "1111111010010101000101",
			2292 => "0000100010000000000100",
			2293 => "1111111010010101000101",
			2294 => "1111110010010101000101",
			2295 => "0001101100011000000100",
			2296 => "0000001010010101000101",
			2297 => "0001010000001100000100",
			2298 => "1111111010010101000101",
			2299 => "0000010010001100000100",
			2300 => "0000001010010101000101",
			2301 => "0000000010010101000101",
			2302 => "0011000100000001001100",
			2303 => "0010011101101000101000",
			2304 => "0010111001110000100000",
			2305 => "0001101010011000010000",
			2306 => "0011101101111000001000",
			2307 => "0011000100010100000100",
			2308 => "0000000010010101000101",
			2309 => "0000001010010101000101",
			2310 => "0011000100010100000100",
			2311 => "0000000010010101000101",
			2312 => "1111111010010101000101",
			2313 => "0001111100001000001000",
			2314 => "0000110000001100000100",
			2315 => "0000000010010101000101",
			2316 => "1111111010010101000101",
			2317 => "0001110100000000000100",
			2318 => "0000000010010101000101",
			2319 => "0000000010010101000101",
			2320 => "0011101110001100000100",
			2321 => "0000000010010101000101",
			2322 => "1111111010010101000101",
			2323 => "0000110010001000100000",
			2324 => "0010101010110000010000",
			2325 => "0000111000000000001000",
			2326 => "0010011011101000000100",
			2327 => "0000001010010101000101",
			2328 => "0000010010010101000101",
			2329 => "0001011101010100000100",
			2330 => "0000000010010101000101",
			2331 => "0000001010010101000101",
			2332 => "0001110100000000001000",
			2333 => "0010101100011100000100",
			2334 => "1111111010010101000101",
			2335 => "0000000010010101000101",
			2336 => "0001000100001100000100",
			2337 => "0000000010010101000101",
			2338 => "0000001010010101000101",
			2339 => "1111111010010101000101",
			2340 => "0001111001110000100100",
			2341 => "0011101101111000010000",
			2342 => "0010101010110000000100",
			2343 => "1111111010010101000101",
			2344 => "0000000100010100000100",
			2345 => "0000001010010101000101",
			2346 => "0000001011000100000100",
			2347 => "0000000010010101000101",
			2348 => "0000001010010101000101",
			2349 => "0010100110011000000100",
			2350 => "0000001010010101000101",
			2351 => "0001001010110100001000",
			2352 => "0000000000111000000100",
			2353 => "1111111010010101000101",
			2354 => "1111111010010101000101",
			2355 => "0001000101010100000100",
			2356 => "0000001010010101000101",
			2357 => "0000000010010101000101",
			2358 => "0001001110100100011000",
			2359 => "0010011110010100001100",
			2360 => "0011001000111100000100",
			2361 => "1111111010010101000101",
			2362 => "0001101001100100000100",
			2363 => "0000000010010101000101",
			2364 => "0000001010010101000101",
			2365 => "0001011111011100000100",
			2366 => "1111111010010101000101",
			2367 => "0001010110110100000100",
			2368 => "0000000010010101000101",
			2369 => "1111111010010101000101",
			2370 => "0000000010111100010000",
			2371 => "0010011010100000001000",
			2372 => "0000001000101100000100",
			2373 => "0000011010010101000101",
			2374 => "0000001010010101000101",
			2375 => "0001110100010000000100",
			2376 => "1111111010010101000101",
			2377 => "0000000010010101000101",
			2378 => "0010110101101100001000",
			2379 => "0000001010000000000100",
			2380 => "0000001010010101000101",
			2381 => "0000000010010101000101",
			2382 => "0010101010110000000100",
			2383 => "1111111010010101000101",
			2384 => "0000000010010101000101",
			2385 => "0011101100001010111000",
			2386 => "0011110010001001110000",
			2387 => "0001000100001100110000",
			2388 => "0000011110100000011000",
			2389 => "0010101010110000010000",
			2390 => "0001101101111100001000",
			2391 => "0000100101110000000100",
			2392 => "0000000010100000110001",
			2393 => "0000000010100000110001",
			2394 => "0000000000110000000100",
			2395 => "0000000010100000110001",
			2396 => "0000001010100000110001",
			2397 => "0011101101010000000100",
			2398 => "1111111010100000110001",
			2399 => "0000000010100000110001",
			2400 => "0001111011000100001100",
			2401 => "0000000100010100001000",
			2402 => "0011011101100000000100",
			2403 => "1111111010100000110001",
			2404 => "0000000010100000110001",
			2405 => "0000001010100000110001",
			2406 => "0001000100001100001000",
			2407 => "0011110110110100000100",
			2408 => "0000000010100000110001",
			2409 => "0000000010100000110001",
			2410 => "1111111010100000110001",
			2411 => "0010000001110100100000",
			2412 => "0001100001111000010000",
			2413 => "0000110100010100001000",
			2414 => "0000110000111000000100",
			2415 => "0000000010100000110001",
			2416 => "1111111010100000110001",
			2417 => "0000010110000000000100",
			2418 => "0000000010100000110001",
			2419 => "0000001010100000110001",
			2420 => "0011100000111000001000",
			2421 => "0011011100110000000100",
			2422 => "1111111010100000110001",
			2423 => "0000001010100000110001",
			2424 => "0000000111111000000100",
			2425 => "0000000010100000110001",
			2426 => "1111111010100000110001",
			2427 => "0011011100101100010000",
			2428 => "0001000010100100001000",
			2429 => "0000010110000000000100",
			2430 => "0000000010100000110001",
			2431 => "0000000010100000110001",
			2432 => "0011110110110100000100",
			2433 => "0000000010100000110001",
			2434 => "1111111010100000110001",
			2435 => "0010101100011100001000",
			2436 => "0010110100000000000100",
			2437 => "1111111010100000110001",
			2438 => "0000000010100000110001",
			2439 => "0001000001101100000100",
			2440 => "0000001010100000110001",
			2441 => "1111111010100000110001",
			2442 => "0011011100101100100100",
			2443 => "0000110101101100011000",
			2444 => "0000011100110100010000",
			2445 => "0011100000101000001000",
			2446 => "0000101100010100000100",
			2447 => "0000000010100000110001",
			2448 => "0000000010100000110001",
			2449 => "0000000100010100000100",
			2450 => "0000001010100000110001",
			2451 => "0000000010100000110001",
			2452 => "0010111100001000000100",
			2453 => "0000000010100000110001",
			2454 => "1111111010100000110001",
			2455 => "0011110001001000001000",
			2456 => "0011100000101000000100",
			2457 => "1111110010100000110001",
			2458 => "1111111010100000110001",
			2459 => "0000000010100000110001",
			2460 => "0001011101111000011000",
			2461 => "0001010110000100001100",
			2462 => "0010110100000000001000",
			2463 => "0001111011000100000100",
			2464 => "0000000010100000110001",
			2465 => "0000001010100000110001",
			2466 => "1111111010100000110001",
			2467 => "0010001011010100000100",
			2468 => "0000000010100000110001",
			2469 => "0010001010101100000100",
			2470 => "0000001010100000110001",
			2471 => "0000000010100000110001",
			2472 => "0000011100110100000100",
			2473 => "1111110010100000110001",
			2474 => "0001001011100000000100",
			2475 => "0000001010100000110001",
			2476 => "0000000010100000110001",
			2477 => "0011010000001101011000",
			2478 => "0001011101111000111000",
			2479 => "0000011100110100100000",
			2480 => "0011111011110100010000",
			2481 => "0010110100000000001000",
			2482 => "0000100100101000000100",
			2483 => "0000000010100000110001",
			2484 => "1111111010100000110001",
			2485 => "0011011101111000000100",
			2486 => "0000001010100000110001",
			2487 => "0000000010100000110001",
			2488 => "0000011100110100001000",
			2489 => "0000110100001000000100",
			2490 => "0000000010100000110001",
			2491 => "1111111010100000110001",
			2492 => "0001011110001100000100",
			2493 => "0000000010100000110001",
			2494 => "1111111010100000110001",
			2495 => "0011101000111000001100",
			2496 => "0000111110001100000100",
			2497 => "0000001010100000110001",
			2498 => "0000111101111000000100",
			2499 => "0000000010100000110001",
			2500 => "0000001010100000110001",
			2501 => "0001000100001100001000",
			2502 => "0001101010011000000100",
			2503 => "0000000010100000110001",
			2504 => "1111111010100000110001",
			2505 => "0000001010100000110001",
			2506 => "0000110001111100011000",
			2507 => "0000011100110100001100",
			2508 => "0001111100001000000100",
			2509 => "0000000010100000110001",
			2510 => "0011010000001100000100",
			2511 => "1111111010100000110001",
			2512 => "0000000010100000110001",
			2513 => "0001000000010100001000",
			2514 => "0000111101111000000100",
			2515 => "0000000010100000110001",
			2516 => "1111111010100000110001",
			2517 => "1111110010100000110001",
			2518 => "0011110010110100000100",
			2519 => "0000001010100000110001",
			2520 => "0000000010100000110001",
			2521 => "0010111000111100101000",
			2522 => "0001100001111000001000",
			2523 => "0000011100110100000100",
			2524 => "1111111010100000110001",
			2525 => "0000000010100000110001",
			2526 => "0011010001111100010000",
			2527 => "0010111000111100001000",
			2528 => "0000111101111000000100",
			2529 => "0000001010100000110001",
			2530 => "0000000010100000110001",
			2531 => "0000111101111000000100",
			2532 => "0000000010100000110001",
			2533 => "0000001010100000110001",
			2534 => "0010101010110000001000",
			2535 => "0010000110001000000100",
			2536 => "0000000010100000110001",
			2537 => "0000001010100000110001",
			2538 => "0001000000010100000100",
			2539 => "1111111010100000110001",
			2540 => "0000000010100000110001",
			2541 => "0010111000111000100000",
			2542 => "0010101010110000010000",
			2543 => "0000101100010100001000",
			2544 => "0000010010001100000100",
			2545 => "0000000010100000110001",
			2546 => "1111111010100000110001",
			2547 => "0000110100011000000100",
			2548 => "0000000010100000110001",
			2549 => "0000001010100000110001",
			2550 => "0001001111100000001000",
			2551 => "0001010000001100000100",
			2552 => "1111110010100000110001",
			2553 => "1111111010100000110001",
			2554 => "0000110001111100000100",
			2555 => "1111111010100000110001",
			2556 => "0000000010100000110001",
			2557 => "0001011100101000010000",
			2558 => "0001111000111000001000",
			2559 => "0010000111000100000100",
			2560 => "0000000010100000110001",
			2561 => "0000000010100000110001",
			2562 => "0011010001111100000100",
			2563 => "0000001010100000110001",
			2564 => "0000000010100000110001",
			2565 => "0011010001111100001000",
			2566 => "0000100010000100000100",
			2567 => "0000000010100000110001",
			2568 => "0000001010100000110001",
			2569 => "0000110100001000000100",
			2570 => "0000001010100000110001",
			2571 => "0000000010100000110001",
			2572 => "0011110000110111010100",
			2573 => "0011101010000001110100",
			2574 => "0010110100010100110100",
			2575 => "0000011110100000011100",
			2576 => "0010011001111000010000",
			2577 => "0011000111111000001000",
			2578 => "0001110111111000000100",
			2579 => "0000000010101100000111",
			2580 => "0000000010101100000111",
			2581 => "0011100011111100000100",
			2582 => "0000000010101100000111",
			2583 => "1111111010101100000111",
			2584 => "0010110100010100001000",
			2585 => "0011000111111000000100",
			2586 => "0000000010101100000111",
			2587 => "0000001010101100000111",
			2588 => "0000000010101100000111",
			2589 => "0011000111111000001100",
			2590 => "0010011001111000000100",
			2591 => "1111111010101100000111",
			2592 => "0000111100001000000100",
			2593 => "0000001010101100000111",
			2594 => "0000000010101100000111",
			2595 => "0001111011000100001000",
			2596 => "0011010101101100000100",
			2597 => "1111111010101100000111",
			2598 => "0000000010101100000111",
			2599 => "0000000010101100000111",
			2600 => "0001100100110100100000",
			2601 => "0011100000111000010000",
			2602 => "0010010010001100001000",
			2603 => "0000010110000000000100",
			2604 => "0000000010101100000111",
			2605 => "1111110010101100000111",
			2606 => "0010001011010100000100",
			2607 => "0000000010101100000111",
			2608 => "0000001010101100000111",
			2609 => "0010011001111000001000",
			2610 => "0001011101100000000100",
			2611 => "0000000010101100000111",
			2612 => "1111111010101100000111",
			2613 => "0011110111010000000100",
			2614 => "0000000010101100000111",
			2615 => "0000000010101100000111",
			2616 => "0011110100000100010000",
			2617 => "0011111000011000001000",
			2618 => "0001000000101100000100",
			2619 => "0000001010101100000111",
			2620 => "1111111010101100000111",
			2621 => "0001111100001000000100",
			2622 => "1111111010101100000111",
			2623 => "0000001010101100000111",
			2624 => "0011011110001100001000",
			2625 => "0001011101100000000100",
			2626 => "0000000010101100000111",
			2627 => "0000001010101100000111",
			2628 => "0010010110101000000100",
			2629 => "1111111010101100000111",
			2630 => "0000001010101100000111",
			2631 => "0011011100101100100100",
			2632 => "0011000000101000100000",
			2633 => "0000110101101100010000",
			2634 => "0011111011011100001000",
			2635 => "0010110100010100000100",
			2636 => "0000001010101100000111",
			2637 => "0000000010101100000111",
			2638 => "0000111001110000000100",
			2639 => "0000000010101100000111",
			2640 => "0000000010101100000111",
			2641 => "0011110111110000001000",
			2642 => "0001000010110000000100",
			2643 => "0000000010101100000111",
			2644 => "1111111010101100000111",
			2645 => "0010000110001000000100",
			2646 => "0000001010101100000111",
			2647 => "0000000010101100000111",
			2648 => "1111111010101100000111",
			2649 => "0011101101100000100000",
			2650 => "0010010111100100010000",
			2651 => "0000011100110100001000",
			2652 => "0010010110101000000100",
			2653 => "0000000010101100000111",
			2654 => "0000000010101100000111",
			2655 => "0011000100000000000100",
			2656 => "0000000010101100000111",
			2657 => "1111111010101100000111",
			2658 => "0001000011001100001000",
			2659 => "0000111110001100000100",
			2660 => "0000001010101100000111",
			2661 => "0000000010101100000111",
			2662 => "0001101010011000000100",
			2663 => "0000001010101100000111",
			2664 => "0000000010101100000111",
			2665 => "0010011011101000010000",
			2666 => "0011000100010100001000",
			2667 => "0011000100010100000100",
			2668 => "0000000010101100000111",
			2669 => "0000001010101100000111",
			2670 => "0010110100000000000100",
			2671 => "1111111010101100000111",
			2672 => "0000000010101100000111",
			2673 => "0010000111000100001000",
			2674 => "0000011001111000000100",
			2675 => "0000000010101100000111",
			2676 => "0000000010101100000111",
			2677 => "0000001010101100000111",
			2678 => "0001110100000001100000",
			2679 => "0010101100011100110100",
			2680 => "0001001010110100011100",
			2681 => "0011000100000000010000",
			2682 => "0001101101111100001000",
			2683 => "0000011110100000000100",
			2684 => "0000000010101100000111",
			2685 => "0000001010101100000111",
			2686 => "0001001011110000000100",
			2687 => "1111111010101100000111",
			2688 => "0000000010101100000111",
			2689 => "0011011010111000001000",
			2690 => "0010000110001000000100",
			2691 => "0000001010101100000111",
			2692 => "0000000010101100000111",
			2693 => "0000000010101100000111",
			2694 => "0011010101101100001100",
			2695 => "0001110111111000001000",
			2696 => "0011111110101100000100",
			2697 => "0000001010101100000111",
			2698 => "0000000010101100000111",
			2699 => "1111111010101100000111",
			2700 => "0011000100000000001000",
			2701 => "0011010000001100000100",
			2702 => "0000000010101100000111",
			2703 => "0000001010101100000111",
			2704 => "0000000010101100000111",
			2705 => "0010111001110000100000",
			2706 => "0001000011010100010000",
			2707 => "0001010000001100001000",
			2708 => "0010010111100100000100",
			2709 => "1111111010101100000111",
			2710 => "0000000010101100000111",
			2711 => "0001101010011000000100",
			2712 => "1111111010101100000111",
			2713 => "1111111010101100000111",
			2714 => "0001111100001000001000",
			2715 => "0011101000111000000100",
			2716 => "0000001010101100000111",
			2717 => "0000000010101100000111",
			2718 => "0011000100010100000100",
			2719 => "0000000010101100000111",
			2720 => "0000001010101100000111",
			2721 => "0011000000101000000100",
			2722 => "1111111010101100000111",
			2723 => "0011101100101100000100",
			2724 => "0000000010101100000111",
			2725 => "0000001010101100000111",
			2726 => "0001111000111000011100",
			2727 => "0011110000110100000100",
			2728 => "0000001010101100000111",
			2729 => "0011000100000000001100",
			2730 => "0001111000111100001000",
			2731 => "0010011011101000000100",
			2732 => "1111111010101100000111",
			2733 => "0000000010101100000111",
			2734 => "1111111010101100000111",
			2735 => "0011001000111000001000",
			2736 => "0001010100001000000100",
			2737 => "0000001010101100000111",
			2738 => "0000000010101100000111",
			2739 => "1111111010101100000111",
			2740 => "0000110100001000000100",
			2741 => "1111111010101100000111",
			2742 => "0010010111100100001000",
			2743 => "0011111110101100000100",
			2744 => "0000001010101100000111",
			2745 => "0000010010101100000111",
			2746 => "0011000000101000001000",
			2747 => "0001101010011000000100",
			2748 => "0000000010101100000111",
			2749 => "0000001010101100000111",
			2750 => "0011000000101000000100",
			2751 => "1111111010101100000111",
			2752 => "0000000010101100000111",
			2753 => "0001000001001101001000",
			2754 => "0001000110111100001000",
			2755 => "0001110100010100000100",
			2756 => "0000000010101111010001",
			2757 => "1111111010101111010001",
			2758 => "0000110011111100001100",
			2759 => "0010111010000000000100",
			2760 => "0000000010101111010001",
			2761 => "0010011100110100000100",
			2762 => "0000001010101111010001",
			2763 => "0000000010101111010001",
			2764 => "0010011100110100011000",
			2765 => "0000110000111000001000",
			2766 => "0011100111000100000100",
			2767 => "1111111010101111010001",
			2768 => "0000001010101111010001",
			2769 => "0011000000111000001000",
			2770 => "0011000011111100000100",
			2771 => "0000000010101111010001",
			2772 => "0000001010101111010001",
			2773 => "0001110111111000000100",
			2774 => "1111111010101111010001",
			2775 => "0000000010101111010001",
			2776 => "0011101000110000001100",
			2777 => "0000101111010000001000",
			2778 => "0000110011010000000100",
			2779 => "1111111010101111010001",
			2780 => "0000001010101111010001",
			2781 => "1111111010101111010001",
			2782 => "0011110010001000001000",
			2783 => "0011100111111000000100",
			2784 => "0000000010101111010001",
			2785 => "0000000010101111010001",
			2786 => "0000111100101100000100",
			2787 => "0000000010101111010001",
			2788 => "0000000010101111010001",
			2789 => "0001111100001000011100",
			2790 => "0011000111111000010100",
			2791 => "0011010100000000000100",
			2792 => "1111111010101111010001",
			2793 => "0011010011011100001100",
			2794 => "0000100111111100001000",
			2795 => "0000101101000100000100",
			2796 => "0000000010101111010001",
			2797 => "0000000010101111010001",
			2798 => "0000000010101111010001",
			2799 => "1111111010101111010001",
			2800 => "0000101111010000000100",
			2801 => "0000000010101111010001",
			2802 => "0000001010101111010001",
			2803 => "1111111010101111010001",
			2804 => "0010011001111000111100",
			2805 => "0001111100001000110100",
			2806 => "0001111100001000110000",
			2807 => "0000111100001000011100",
			2808 => "0000100111111100010000",
			2809 => "0001000011010100001000",
			2810 => "0000101111010000000100",
			2811 => "0000000010110011101101",
			2812 => "0000001010110011101101",
			2813 => "0011100011111100000100",
			2814 => "0000000010110011101101",
			2815 => "1111111010110011101101",
			2816 => "0010011100110100000100",
			2817 => "1111111010110011101101",
			2818 => "0001010011011100000100",
			2819 => "0000001010110011101101",
			2820 => "0000000010110011101101",
			2821 => "0001010110000100010000",
			2822 => "0000101110101000001000",
			2823 => "0010001100000100000100",
			2824 => "0000000010110011101101",
			2825 => "1111111010110011101101",
			2826 => "0011000100010100000100",
			2827 => "0000000010110011101101",
			2828 => "0000000010110011101101",
			2829 => "0000001010110011101101",
			2830 => "1111111010110011101101",
			2831 => "0001000010010000000100",
			2832 => "0000001010110011101101",
			2833 => "1111111010110011101101",
			2834 => "0011100011010000010000",
			2835 => "0000101010010100000100",
			2836 => "0000000010110011101101",
			2837 => "0010011001111000001000",
			2838 => "0001001001001100000100",
			2839 => "0000001010110011101101",
			2840 => "0000000010110011101101",
			2841 => "0000001010110011101101",
			2842 => "0011001010000000010100",
			2843 => "0011100100000000001100",
			2844 => "0010100110011000000100",
			2845 => "0000001010110011101101",
			2846 => "0001000100001100000100",
			2847 => "0000000010110011101101",
			2848 => "0000001010110011101101",
			2849 => "0000101010001000000100",
			2850 => "1111111010110011101101",
			2851 => "0000001010110011101101",
			2852 => "0011001110111100010000",
			2853 => "0000101100010100001100",
			2854 => "0011010101101100000100",
			2855 => "1111111010110011101101",
			2856 => "0010001111001000000100",
			2857 => "0000000010110011101101",
			2858 => "0000001010110011101101",
			2859 => "1111111010110011101101",
			2860 => "0001000100001100010000",
			2861 => "0000000100010100001000",
			2862 => "0010000001110100000100",
			2863 => "0000000010110011101101",
			2864 => "0000000010110011101101",
			2865 => "0011101100110000000100",
			2866 => "0000001010110011101101",
			2867 => "0000000010110011101101",
			2868 => "0010000111000100001000",
			2869 => "0001111100001000000100",
			2870 => "0000000010110011101101",
			2871 => "1111111010110011101101",
			2872 => "0010000010101000000100",
			2873 => "0000000010110011101101",
			2874 => "0000000010110011101101",
			2875 => "0011001110001101011100",
			2876 => "0001001011100101010000",
			2877 => "0001000000010000010000",
			2878 => "0011101000111000000100",
			2879 => "0000000010111000101001",
			2880 => "0010111110001100000100",
			2881 => "1111111010111000101001",
			2882 => "0010111101111000000100",
			2883 => "0000000010111000101001",
			2884 => "1111111010111000101001",
			2885 => "0011000000101000100000",
			2886 => "0011100000001100010000",
			2887 => "0010011101101000001000",
			2888 => "0011101100001000000100",
			2889 => "0000000010111000101001",
			2890 => "0000000010111000101001",
			2891 => "0011111001010100000100",
			2892 => "0000000010111000101001",
			2893 => "0000001010111000101001",
			2894 => "0011000100010100001000",
			2895 => "0001101101011000000100",
			2896 => "0000000010111000101001",
			2897 => "1111111010111000101001",
			2898 => "0010110101101100000100",
			2899 => "1111111010111000101001",
			2900 => "0000001010111000101001",
			2901 => "0011000000101000010000",
			2902 => "0010100110011000001000",
			2903 => "0000100111111100000100",
			2904 => "0000001010111000101001",
			2905 => "0000010010111000101001",
			2906 => "0010001011010100000100",
			2907 => "1111111010111000101001",
			2908 => "0000001010111000101001",
			2909 => "0011000000101000001000",
			2910 => "0000100101110000000100",
			2911 => "0000000010111000101001",
			2912 => "1111111010111000101001",
			2913 => "0011111101000100000100",
			2914 => "0000000010111000101001",
			2915 => "0000000010111000101001",
			2916 => "0010010110000000000100",
			2917 => "1111111010111000101001",
			2918 => "0011111001001000000100",
			2919 => "0000001010111000101001",
			2920 => "1111111010111000101001",
			2921 => "0010001001101000001100",
			2922 => "0011101010001100001000",
			2923 => "0001010100000100000100",
			2924 => "0000000010111000101001",
			2925 => "0000001010111000101001",
			2926 => "1111111010111000101001",
			2927 => "0001000110110000101100",
			2928 => "0010000110001000010000",
			2929 => "0000100101000000001100",
			2930 => "0001011111010000001000",
			2931 => "0011110110111000000100",
			2932 => "0000001010111000101001",
			2933 => "1111111010111000101001",
			2934 => "0000001010111000101001",
			2935 => "1111111010111000101001",
			2936 => "0001000011101100010000",
			2937 => "0001001001001100001000",
			2938 => "0010101100011100000100",
			2939 => "0000000010111000101001",
			2940 => "1111111010111000101001",
			2941 => "0011101000001000000100",
			2942 => "0000001010111000101001",
			2943 => "0000000010111000101001",
			2944 => "0010000001110100000100",
			2945 => "1111111010111000101001",
			2946 => "0001101001111100000100",
			2947 => "0000000010111000101001",
			2948 => "0000001010111000101001",
			2949 => "0011000000001100001000",
			2950 => "0001000011000100000100",
			2951 => "0000001010111000101001",
			2952 => "1111111010111000101001",
			2953 => "1111111010111000101001",
			2954 => "0001000001001101111000",
			2955 => "0010001101010001101000",
			2956 => "0001000011011001000000",
			2957 => "0011100011010000100000",
			2958 => "0011110001101000010000",
			2959 => "0011101000110000001000",
			2960 => "0001011000111000000100",
			2961 => "0000000010111101000101",
			2962 => "0000001010111101000101",
			2963 => "0001110000101000000100",
			2964 => "1111111010111101000101",
			2965 => "0000001010111101000101",
			2966 => "0010010010001100001000",
			2967 => "0011101111000100000100",
			2968 => "0000001010111101000101",
			2969 => "0000000010111101000101",
			2970 => "0001110000101000000100",
			2971 => "0000001010111101000101",
			2972 => "0000000010111101000101",
			2973 => "0001110111111000010000",
			2974 => "0001111110111100001000",
			2975 => "0011001010000000000100",
			2976 => "1111111010111101000101",
			2977 => "0000001010111101000101",
			2978 => "0011000000110000000100",
			2979 => "0000000010111101000101",
			2980 => "1111111010111101000101",
			2981 => "0011110101100100001000",
			2982 => "0010110100010100000100",
			2983 => "1111111010111101000101",
			2984 => "0000000010111101000101",
			2985 => "0001101010011000000100",
			2986 => "0000000010111101000101",
			2987 => "0000000010111101000101",
			2988 => "0011111001001000001000",
			2989 => "0011000111111000000100",
			2990 => "0000000010111101000101",
			2991 => "0000001010111101000101",
			2992 => "0010000111000000010000",
			2993 => "0010100110011100001000",
			2994 => "0010000010101000000100",
			2995 => "1111111010111101000101",
			2996 => "0000000010111101000101",
			2997 => "0000101111010100000100",
			2998 => "1111110010111101000101",
			2999 => "1111111010111101000101",
			3000 => "0011000100010100001000",
			3001 => "0001111011000100000100",
			3002 => "0000000010111101000101",
			3003 => "1111111010111101000101",
			3004 => "0010100001010100000100",
			3005 => "0000001010111101000101",
			3006 => "0000000010111101000101",
			3007 => "0001101010011000000100",
			3008 => "0000000010111101000101",
			3009 => "0010101001101000001000",
			3010 => "0010101100000100000100",
			3011 => "0000001010111101000101",
			3012 => "0000000010111101000101",
			3013 => "0000001010111101000101",
			3014 => "0001111100001000010100",
			3015 => "0011000111111000001100",
			3016 => "0001011001110000000100",
			3017 => "1111111010111101000101",
			3018 => "0001010011011100000100",
			3019 => "0000000010111101000101",
			3020 => "1111111010111101000101",
			3021 => "0001000100100000000100",
			3022 => "0000000010111101000101",
			3023 => "0000000010111101000101",
			3024 => "1111111010111101000101",
			3025 => "0011100011111101010100",
			3026 => "0001001001000000101000",
			3027 => "0000101111010000011100",
			3028 => "0000000000101000010100",
			3029 => "0001000010100100001100",
			3030 => "0010000010101000001000",
			3031 => "0000000100010100000100",
			3032 => "0000000011000011110001",
			3033 => "0000001011000011110001",
			3034 => "1111111011000011110001",
			3035 => "0011011101100000000100",
			3036 => "0000000011000011110001",
			3037 => "1111110011000011110001",
			3038 => "0010101100011100000100",
			3039 => "0000000011000011110001",
			3040 => "0000001011000011110001",
			3041 => "0010011100110100000100",
			3042 => "1111111011000011110001",
			3043 => "0000000100010100000100",
			3044 => "0000000011000011110001",
			3045 => "0000001011000011110001",
			3046 => "0010010010001100100100",
			3047 => "0011011101100000011000",
			3048 => "0001010011011100010000",
			3049 => "0001100100110100001000",
			3050 => "0001110100010100000100",
			3051 => "1111111011000011110001",
			3052 => "0000000011000011110001",
			3053 => "0001011001110000000100",
			3054 => "0000000011000011110001",
			3055 => "0000001011000011110001",
			3056 => "0010010000011000000100",
			3057 => "0000000011000011110001",
			3058 => "1111110011000011110001",
			3059 => "0001000110110000000100",
			3060 => "0000001011000011110001",
			3061 => "0001110100010100000100",
			3062 => "0000000011000011110001",
			3063 => "1111111011000011110001",
			3064 => "0001001100111100000100",
			3065 => "0000001011000011110001",
			3066 => "0000000011000011110001",
			3067 => "0010011001111000111100",
			3068 => "0011111010001100011000",
			3069 => "0001001101001000010000",
			3070 => "0001000110001100001000",
			3071 => "0011110001101000000100",
			3072 => "0000000011000011110001",
			3073 => "1111111011000011110001",
			3074 => "0011100011010000000100",
			3075 => "0000001011000011110001",
			3076 => "0000000011000011110001",
			3077 => "0010101010110000000100",
			3078 => "1111110011000011110001",
			3079 => "1111111011000011110001",
			3080 => "0000110000101000000100",
			3081 => "0000001011000011110001",
			3082 => "0010101001000100010000",
			3083 => "0000110100000000001000",
			3084 => "0010010010001100000100",
			3085 => "1111111011000011110001",
			3086 => "0000001011000011110001",
			3087 => "0000000011010000000100",
			3088 => "0000000011000011110001",
			3089 => "0000001011000011110001",
			3090 => "0011110110110100001000",
			3091 => "0000111000111100000100",
			3092 => "0000000011000011110001",
			3093 => "1111111011000011110001",
			3094 => "0000100100101000000100",
			3095 => "0000001011000011110001",
			3096 => "0000000011000011110001",
			3097 => "0001010011011100010100",
			3098 => "0001101101111100001100",
			3099 => "0000000011111100000100",
			3100 => "1111111011000011110001",
			3101 => "0011110110110100000100",
			3102 => "0000001011000011110001",
			3103 => "0000000011000011110001",
			3104 => "0010110100010100000100",
			3105 => "1111111011000011110001",
			3106 => "0000000011000011110001",
			3107 => "0000111100110000010100",
			3108 => "0011011101111000010000",
			3109 => "0011111111011100001000",
			3110 => "0000111000111100000100",
			3111 => "0000000011000011110001",
			3112 => "1111111011000011110001",
			3113 => "0001110111111000000100",
			3114 => "1111111011000011110001",
			3115 => "0000000011000011110001",
			3116 => "0000001011000011110001",
			3117 => "0011111010010100010000",
			3118 => "0010010110101000001000",
			3119 => "0011110111110000000100",
			3120 => "1111111011000011110001",
			3121 => "0000000011000011110001",
			3122 => "0011110111110000000100",
			3123 => "0000000011000011110001",
			3124 => "0000000011000011110001",
			3125 => "0000111101111000001000",
			3126 => "0000000000110000000100",
			3127 => "0000001011000011110001",
			3128 => "0000000011000011110001",
			3129 => "0010010111100100000100",
			3130 => "0000000011000011110001",
			3131 => "0000000011000011110001",
			3132 => "0010000111000001101100",
			3133 => "0010100110011101001100",
			3134 => "0000110000110000001100",
			3135 => "0001101110010100000100",
			3136 => "1111111011001001110101",
			3137 => "0010111110111100000100",
			3138 => "0000000011001001110101",
			3139 => "0000001011001001110101",
			3140 => "0010011001111000100000",
			3141 => "0000111000111100010000",
			3142 => "0000101111010000001000",
			3143 => "0001000010111000000100",
			3144 => "0000000011001001110101",
			3145 => "0000000011001001110101",
			3146 => "0011000111111000000100",
			3147 => "0000000011001001110101",
			3148 => "0000001011001001110101",
			3149 => "0001011101100000001000",
			3150 => "0001100100110100000100",
			3151 => "0000000011001001110101",
			3152 => "0000001011001001110101",
			3153 => "0011101110111100000100",
			3154 => "0000000011001001110101",
			3155 => "1111111011001001110101",
			3156 => "0000011110100000010000",
			3157 => "0001011100110000001000",
			3158 => "0001010011011100000100",
			3159 => "0000000011001001110101",
			3160 => "0000000011001001110101",
			3161 => "0001110100010100000100",
			3162 => "1111111011001001110101",
			3163 => "0000000011001001110101",
			3164 => "0010010110101000001000",
			3165 => "0001110100010100000100",
			3166 => "0000000011001001110101",
			3167 => "0000000011001001110101",
			3168 => "0011100000101000000100",
			3169 => "0000000011001001110101",
			3170 => "0000000011001001110101",
			3171 => "0010010110101000000100",
			3172 => "1111110011001001110101",
			3173 => "0010111000111100001000",
			3174 => "0001001111100000000100",
			3175 => "1111111011001001110101",
			3176 => "0000001011001001110101",
			3177 => "0010011011101000001000",
			3178 => "0011101101100000000100",
			3179 => "0000000011001001110101",
			3180 => "1111111011001001110101",
			3181 => "0011101010111000000100",
			3182 => "0000001011001001110101",
			3183 => "0000011001111000000100",
			3184 => "1111111011001001110101",
			3185 => "0000000011001001110101",
			3186 => "0001000011011000010100",
			3187 => "0001001001000000010000",
			3188 => "0010111011000100000100",
			3189 => "0000001011001001110101",
			3190 => "0010111100001000000100",
			3191 => "1111111011001001110101",
			3192 => "0001101011001100000100",
			3193 => "0000001011001001110101",
			3194 => "0000000011001001110101",
			3195 => "0000001011001001110101",
			3196 => "0011000111111000011000",
			3197 => "0010110100010100010000",
			3198 => "0001110111111000000100",
			3199 => "1111111011001001110101",
			3200 => "0001000110110000000100",
			3201 => "0000001011001001110101",
			3202 => "0010100110001000000100",
			3203 => "1111111011001001110101",
			3204 => "0000000011001001110101",
			3205 => "0000111000101100000100",
			3206 => "0000000011001001110101",
			3207 => "1111110011001001110101",
			3208 => "0001111011000100010100",
			3209 => "0001000010010000001000",
			3210 => "0001011101100000000100",
			3211 => "0000001011001001110101",
			3212 => "0000000011001001110101",
			3213 => "0001100100110100001000",
			3214 => "0010101100000100000100",
			3215 => "1111111011001001110101",
			3216 => "0000000011001001110101",
			3217 => "0000000011001001110101",
			3218 => "0011000100010100001000",
			3219 => "0001111100001000000100",
			3220 => "1111111011001001110101",
			3221 => "0000000011001001110101",
			3222 => "0000001100101100001000",
			3223 => "0010010110101000000100",
			3224 => "0000001011001001110101",
			3225 => "0000000011001001110101",
			3226 => "0000101110110100000100",
			3227 => "0000000011001001110101",
			3228 => "1111111011001001110101",
			3229 => "0001111100101001100100",
			3230 => "0001000110110001000100",
			3231 => "0001100001000100000100",
			3232 => "1111111011001111011001",
			3233 => "0011100100010100100000",
			3234 => "0001010110000100010000",
			3235 => "0000110111111000001000",
			3236 => "0010011100110100000100",
			3237 => "0000000011001111011001",
			3238 => "0000001011001111011001",
			3239 => "0010011100110100000100",
			3240 => "1111111011001111011001",
			3241 => "0000000011001111011001",
			3242 => "0010110100000000001000",
			3243 => "0011111000011000000100",
			3244 => "0000000011001111011001",
			3245 => "0000001011001111011001",
			3246 => "0001111100001000000100",
			3247 => "0000000011001111011001",
			3248 => "0000001011001111011001",
			3249 => "0000101010001000010000",
			3250 => "0001100001111000001000",
			3251 => "0001011110001100000100",
			3252 => "0000000011001111011001",
			3253 => "0000001011001111011001",
			3254 => "0000101110000100000100",
			3255 => "0000000011001111011001",
			3256 => "0000000011001111011001",
			3257 => "0001101100011000001000",
			3258 => "0011010101101100000100",
			3259 => "0000000011001111011001",
			3260 => "0000001011001111011001",
			3261 => "0001000100001100000100",
			3262 => "0000000011001111011001",
			3263 => "0000000011001111011001",
			3264 => "0000100010010100011100",
			3265 => "0000011110100000010100",
			3266 => "0011101000101100001100",
			3267 => "0000011100100000000100",
			3268 => "1111111011001111011001",
			3269 => "0001000011111000000100",
			3270 => "1111111011001111011001",
			3271 => "0000000011001111011001",
			3272 => "0000010000011000000100",
			3273 => "1111111011001111011001",
			3274 => "1111110011001111011001",
			3275 => "0011100100000000000100",
			3276 => "0000000011001111011001",
			3277 => "1111111011001111011001",
			3278 => "0000000011001111011001",
			3279 => "0010001001101000010100",
			3280 => "0011000110000100001000",
			3281 => "0011000110000100000100",
			3282 => "1111111011001111011001",
			3283 => "0000001011001111011001",
			3284 => "0011101010001100001000",
			3285 => "0001010100000100000100",
			3286 => "1111111011001111011001",
			3287 => "0000001011001111011001",
			3288 => "1111111011001111011001",
			3289 => "0001000010010000100100",
			3290 => "0010000111000000100000",
			3291 => "0011111011110000010000",
			3292 => "0001000011110100001000",
			3293 => "0011000100001000000100",
			3294 => "0000000011001111011001",
			3295 => "0000001011001111011001",
			3296 => "0010011101011000000100",
			3297 => "0000000011001111011001",
			3298 => "1111111011001111011001",
			3299 => "0011000111010000001000",
			3300 => "0010000111000100000100",
			3301 => "1111111011001111011001",
			3302 => "0000000011001111011001",
			3303 => "0011110010111000000100",
			3304 => "0000010011001111011001",
			3305 => "0000000011001111011001",
			3306 => "0000001011001111011001",
			3307 => "0001000000000000010100",
			3308 => "0010000000110000001100",
			3309 => "0001000011111000001000",
			3310 => "0001001011100100000100",
			3311 => "1111111011001111011001",
			3312 => "0000000011001111011001",
			3313 => "1111111011001111011001",
			3314 => "0010001010000000000100",
			3315 => "0000001011001111011001",
			3316 => "1111111011001111011001",
			3317 => "1111111011001111011001",
			3318 => "0001111110001110000000",
			3319 => "0000010000011000010000",
			3320 => "0000011100100000000100",
			3321 => "1111111011010101001101",
			3322 => "0000111000110000000100",
			3323 => "0000001011010101001101",
			3324 => "0001110111111000000100",
			3325 => "1111111011010101001101",
			3326 => "0000000011010101001101",
			3327 => "0011101101100000111100",
			3328 => "0000000100010100100000",
			3329 => "0000110100000000010000",
			3330 => "0010011100110100001000",
			3331 => "0000110000111000000100",
			3332 => "0000010011010101001101",
			3333 => "1111111011010101001101",
			3334 => "0001000011010100000100",
			3335 => "0000001011010101001101",
			3336 => "0000000011010101001101",
			3337 => "0010010010001100001000",
			3338 => "0011000111111000000100",
			3339 => "1111111011010101001101",
			3340 => "1111111011010101001101",
			3341 => "0000101010001000000100",
			3342 => "0000001011010101001101",
			3343 => "0000001011010101001101",
			3344 => "0001000110110000010000",
			3345 => "0001110111111000001000",
			3346 => "0000101110000100000100",
			3347 => "0000001011010101001101",
			3348 => "0000000011010101001101",
			3349 => "0010000111000000000100",
			3350 => "0000001011010101001101",
			3351 => "0000001011010101001101",
			3352 => "0000001101111000000100",
			3353 => "1111111011010101001101",
			3354 => "0011111110101100000100",
			3355 => "0000001011010101001101",
			3356 => "1111111011010101001101",
			3357 => "0001001101001000011000",
			3358 => "0001000000010000001000",
			3359 => "0011000100000000000100",
			3360 => "0000000011010101001101",
			3361 => "1111111011010101001101",
			3362 => "0011001000111000001000",
			3363 => "0010100111110100000100",
			3364 => "0000001011010101001101",
			3365 => "0000000011010101001101",
			3366 => "0001111001110000000100",
			3367 => "0000000011010101001101",
			3368 => "0000001011010101001101",
			3369 => "0011011000000000010000",
			3370 => "0001111100001000001000",
			3371 => "0011110010110100000100",
			3372 => "1111111011010101001101",
			3373 => "0000001011010101001101",
			3374 => "0001111001110000000100",
			3375 => "0000001011010101001101",
			3376 => "0000001011010101001101",
			3377 => "0000000011010000000100",
			3378 => "0000001011010101001101",
			3379 => "0000011001111000000100",
			3380 => "0000001011010101001101",
			3381 => "0000000011010101001101",
			3382 => "0001111100101000011000",
			3383 => "0001000111011100001100",
			3384 => "0010101001000100000100",
			3385 => "1111111011010101001101",
			3386 => "0011000110000100000100",
			3387 => "0000000011010101001101",
			3388 => "0000010011010101001101",
			3389 => "0001111101111000001000",
			3390 => "0011101000000000000100",
			3391 => "1111111011010101001101",
			3392 => "0000001011010101001101",
			3393 => "1111111011010101001101",
			3394 => "0010001001101000000100",
			3395 => "1111111011010101001101",
			3396 => "0001000110110000011100",
			3397 => "0010001111001000001100",
			3398 => "0010011101011000000100",
			3399 => "0000001011010101001101",
			3400 => "0011001011011100000100",
			3401 => "1111111011010101001101",
			3402 => "0000000011010101001101",
			3403 => "0000101110111000001000",
			3404 => "0001001001001100000100",
			3405 => "1111111011010101001101",
			3406 => "0000001011010101001101",
			3407 => "0001010110111100000100",
			3408 => "1111111011010101001101",
			3409 => "0000001011010101001101",
			3410 => "1111111011010101001101",
			3411 => "0001111101111010001000",
			3412 => "0000010000011000011000",
			3413 => "0000101010010100001000",
			3414 => "0001011000111100000100",
			3415 => "1111111011011011101001",
			3416 => "0000001011011011101001",
			3417 => "0001101100011000001000",
			3418 => "0000100001001000000100",
			3419 => "0000000011011011101001",
			3420 => "1111111011011011101001",
			3421 => "0010101000101100000100",
			3422 => "0000000011011011101001",
			3423 => "1111111011011011101001",
			3424 => "0011101101111001000000",
			3425 => "0001111100001000100000",
			3426 => "0000111101100000010000",
			3427 => "0001110111111000001000",
			3428 => "0000100001000000000100",
			3429 => "0000000011011011101001",
			3430 => "1111111011011011101001",
			3431 => "0000111011000100000100",
			3432 => "0000001011011011101001",
			3433 => "0000000011011011101001",
			3434 => "0000100100101000001000",
			3435 => "0010010110101000000100",
			3436 => "1111111011011011101001",
			3437 => "0000000011011011101001",
			3438 => "0010011001111000000100",
			3439 => "0000000011011011101001",
			3440 => "0000000011011011101001",
			3441 => "0011011110110000010000",
			3442 => "0000101100010100001000",
			3443 => "0001100001111000000100",
			3444 => "0000001011011011101001",
			3445 => "0000000011011011101001",
			3446 => "0010000111000100000100",
			3447 => "0000001011011011101001",
			3448 => "0000001011011011101001",
			3449 => "0001101010011000001000",
			3450 => "0000100001001000000100",
			3451 => "1111111011011011101001",
			3452 => "1111111011011011101001",
			3453 => "0000100111011000000100",
			3454 => "0000001011011011101001",
			3455 => "1111111011011011101001",
			3456 => "0000100011001000010100",
			3457 => "0001011000000000010000",
			3458 => "0001111000111000001000",
			3459 => "0000011001111000000100",
			3460 => "0000000011011011101001",
			3461 => "0000001011011011101001",
			3462 => "0001101100011000000100",
			3463 => "0000000011011011101001",
			3464 => "0000001011011011101001",
			3465 => "1111111011011011101001",
			3466 => "0001101100011000001100",
			3467 => "0001101101111100000100",
			3468 => "0000000011011011101001",
			3469 => "0010001001101000000100",
			3470 => "0000000011011011101001",
			3471 => "0000010011011011101001",
			3472 => "0001111001110000001000",
			3473 => "0001000000010100000100",
			3474 => "0000000011011011101001",
			3475 => "0000000011011011101001",
			3476 => "0011011000000000000100",
			3477 => "0000001011011011101001",
			3478 => "0000000011011011101001",
			3479 => "0010001001101000001100",
			3480 => "0000011011101000001000",
			3481 => "0000011011101000000100",
			3482 => "1111111011011011101001",
			3483 => "0000001011011011101001",
			3484 => "1111111011011011101001",
			3485 => "0001000010010000101100",
			3486 => "0010000001110100011000",
			3487 => "0011101011110000001100",
			3488 => "0001001011100000001000",
			3489 => "0001000010111000000100",
			3490 => "0000000011011011101001",
			3491 => "0000001011011011101001",
			3492 => "1111111011011011101001",
			3493 => "0001101001111100000100",
			3494 => "1111111011011011101001",
			3495 => "0001100100101100000100",
			3496 => "0000000011011011101001",
			3497 => "1111111011011011101001",
			3498 => "0001001101110100001100",
			3499 => "0000101101001000001000",
			3500 => "0000101100001100000100",
			3501 => "0000001011011011101001",
			3502 => "0000000011011011101001",
			3503 => "0000001011011011101001",
			3504 => "0010001010101100000100",
			3505 => "1111111011011011101001",
			3506 => "0000001011011011101001",
			3507 => "0001000000000000001100",
			3508 => "0010000000110000000100",
			3509 => "1111111011011011101001",
			3510 => "0010001010000000000100",
			3511 => "0000000011011011101001",
			3512 => "1111111011011011101001",
			3513 => "1111111011011011101001",
			3514 => "0000000010101000110000",
			3515 => "0001100111101000010000",
			3516 => "0011111000000000000100",
			3517 => "1111111011100010011101",
			3518 => "0010001000010100000100",
			3519 => "0000000011100010011101",
			3520 => "0000011110100000000100",
			3521 => "0000000011100010011101",
			3522 => "0000001011100010011101",
			3523 => "0010000110011100011000",
			3524 => "0001100111101000001000",
			3525 => "0010000011101000000100",
			3526 => "0000000011100010011101",
			3527 => "1111110011100010011101",
			3528 => "0001100001111000001100",
			3529 => "0001100001111000000100",
			3530 => "1111111011100010011101",
			3531 => "0001100001111000000100",
			3532 => "0000000011100010011101",
			3533 => "0000000011100010011101",
			3534 => "1111111011100010011101",
			3535 => "0001101011001100000100",
			3536 => "0000001011100010011101",
			3537 => "1111111011100010011101",
			3538 => "0010011111001101100000",
			3539 => "0001110100000000101000",
			3540 => "0001110100000000011100",
			3541 => "0001110100000000010000",
			3542 => "0001111100001000001000",
			3543 => "0001111100001000000100",
			3544 => "0000000011100010011101",
			3545 => "0000000011100010011101",
			3546 => "0010110100000000000100",
			3547 => "1111111011100010011101",
			3548 => "0000000011100010011101",
			3549 => "0011000100010100000100",
			3550 => "1111111011100010011101",
			3551 => "0011011101111000000100",
			3552 => "0000001011100010011101",
			3553 => "0000000011100010011101",
			3554 => "0011101110001100001000",
			3555 => "0001101100011000000100",
			3556 => "0000001011100010011101",
			3557 => "0000001011100010011101",
			3558 => "0000000011100010011101",
			3559 => "0001111000111000011100",
			3560 => "0010000110001000001100",
			3561 => "0001000010111000001000",
			3562 => "0000000011111100000100",
			3563 => "0000000011100010011101",
			3564 => "1111111011100010011101",
			3565 => "0000001011100010011101",
			3566 => "0000110000001100001000",
			3567 => "0000111101111000000100",
			3568 => "0000000011100010011101",
			3569 => "0000001011100010011101",
			3570 => "0000010010001100000100",
			3571 => "1111111011100010011101",
			3572 => "0000000011100010011101",
			3573 => "0011111001010000010000",
			3574 => "0010010111100100001000",
			3575 => "0010111101100000000100",
			3576 => "0000000011100010011101",
			3577 => "1111110011100010011101",
			3578 => "0010010111100100000100",
			3579 => "0000001011100010011101",
			3580 => "0000000011100010011101",
			3581 => "0000011001111000001000",
			3582 => "0001111001110000000100",
			3583 => "1111111011100010011101",
			3584 => "0000000011100010011101",
			3585 => "0000000011100010011101",
			3586 => "0011000000101000001100",
			3587 => "0011000000101000001000",
			3588 => "0010111101100000000100",
			3589 => "0000001011100010011101",
			3590 => "1111111011100010011101",
			3591 => "0000001011100010011101",
			3592 => "0011101010111000100000",
			3593 => "0000100110010000010000",
			3594 => "0011101101010100001000",
			3595 => "0010000110001000000100",
			3596 => "0000000011100010011101",
			3597 => "0000001011100010011101",
			3598 => "0000111001001000000100",
			3599 => "0000010011100010011101",
			3600 => "0000001011100010011101",
			3601 => "0011101101010100001000",
			3602 => "0011011001001000000100",
			3603 => "0000001011100010011101",
			3604 => "0000000011100010011101",
			3605 => "0001101011001100000100",
			3606 => "1111111011100010011101",
			3607 => "0000001011100010011101",
			3608 => "0011111110101000010000",
			3609 => "0001000110111000001000",
			3610 => "0010000001110000000100",
			3611 => "0000000011100010011101",
			3612 => "0000001011100010011101",
			3613 => "0001111001110000000100",
			3614 => "1111111011100010011101",
			3615 => "1111111011100010011101",
			3616 => "0001111000111000001000",
			3617 => "0000101100010000000100",
			3618 => "1111111011100010011101",
			3619 => "0000000011100010011101",
			3620 => "0000111111011100000100",
			3621 => "0000001011100010011101",
			3622 => "0000000011100010011101",
			3623 => "0001010100011001111000",
			3624 => "0000010000011000011100",
			3625 => "0001101101111100010000",
			3626 => "0001101101111100001000",
			3627 => "0000100101110100000100",
			3628 => "1110011011101010010001",
			3629 => "1110010011101010010001",
			3630 => "0001011000111100000100",
			3631 => "1110011011101010010001",
			3632 => "1110011011101010010001",
			3633 => "0000111000110000000100",
			3634 => "1110111011101010010001",
			3635 => "0000100001000000000100",
			3636 => "1110101011101010010001",
			3637 => "1110011011101010010001",
			3638 => "0000111101100000101000",
			3639 => "0001100001000100001000",
			3640 => "0001011001110000000100",
			3641 => "1110010011101010010001",
			3642 => "1110011011101010010001",
			3643 => "0000111001110000010000",
			3644 => "0001110111111000001000",
			3645 => "0011000000110000000100",
			3646 => "1110100011101010010001",
			3647 => "1110110011101010010001",
			3648 => "0000110100010100000100",
			3649 => "1110111011101010010001",
			3650 => "1110110011101010010001",
			3651 => "0011011100101100001000",
			3652 => "0001110000101000000100",
			3653 => "1110100011101010010001",
			3654 => "1110110011101010010001",
			3655 => "0010010110101000000100",
			3656 => "1110101011101010010001",
			3657 => "1110111011101010010001",
			3658 => "0000000000110000011000",
			3659 => "0001101011111100001000",
			3660 => "0001100001000100000100",
			3661 => "1110010011101010010001",
			3662 => "1110011011101010010001",
			3663 => "0001101101111100001000",
			3664 => "0001111011000100000100",
			3665 => "1110100011101010010001",
			3666 => "1110110011101010010001",
			3667 => "0000000011111100000100",
			3668 => "1110100011101010010001",
			3669 => "1110100011101010010001",
			3670 => "0001101011001100010000",
			3671 => "0000000111111000001000",
			3672 => "0001110000101000000100",
			3673 => "1110100011101010010001",
			3674 => "1110110011101010010001",
			3675 => "0010011001111000000100",
			3676 => "1110101011101010010001",
			3677 => "1110110011101010010001",
			3678 => "0001111101100000001000",
			3679 => "0000111010111100000100",
			3680 => "1110101011101010010001",
			3681 => "1110011011101010010001",
			3682 => "1110101011101010010001",
			3683 => "0001111110001101001000",
			3684 => "0000110001101000010100",
			3685 => "0011000110000100010000",
			3686 => "0011011001001000001000",
			3687 => "0000111001110100000100",
			3688 => "1110010011101010010001",
			3689 => "1110101011101010010001",
			3690 => "0011001100110000000100",
			3691 => "1110010011101010010001",
			3692 => "1110011011101010010001",
			3693 => "1110100011101010010001",
			3694 => "0001101001100100011000",
			3695 => "0000000001110100001000",
			3696 => "0001110101101100000100",
			3697 => "1110011011101010010001",
			3698 => "1110010011101010010001",
			3699 => "0010000010101000001000",
			3700 => "0001111001110000000100",
			3701 => "1110011011101010010001",
			3702 => "1110110011101010010001",
			3703 => "0000001100110000000100",
			3704 => "1110011011101010010001",
			3705 => "1110011011101010010001",
			3706 => "0001110110000100010000",
			3707 => "0000010111100100001000",
			3708 => "0000000011010000000100",
			3709 => "1110100011101010010001",
			3710 => "1110011011101010010001",
			3711 => "0010000111000100000100",
			3712 => "1110010011101010010001",
			3713 => "1110011011101010010001",
			3714 => "0000101000100000000100",
			3715 => "1110111011101010010001",
			3716 => "0000111101000100000100",
			3717 => "1110010011101010010001",
			3718 => "1110100011101010010001",
			3719 => "0010011000010100110100",
			3720 => "0001111101111000011000",
			3721 => "0011110110010000010000",
			3722 => "0011011000011000001000",
			3723 => "0011111110101100000100",
			3724 => "1110010011101010010001",
			3725 => "1110101011101010010001",
			3726 => "0000110000110100000100",
			3727 => "1110010011101010010001",
			3728 => "1110011011101010010001",
			3729 => "0011001100110000000100",
			3730 => "1110010011101010010001",
			3731 => "1110110011101010010001",
			3732 => "0010001001101000001100",
			3733 => "0011000110000100001000",
			3734 => "0011000110000100000100",
			3735 => "1110010011101010010001",
			3736 => "1110011011101010010001",
			3737 => "1110010011101010010001",
			3738 => "0000001000111100001000",
			3739 => "0000011101101000000100",
			3740 => "1110111011101010010001",
			3741 => "1110011011101010010001",
			3742 => "0010100001010100000100",
			3743 => "1110011011101010010001",
			3744 => "1110010011101010010001",
			3745 => "0000000011010000000100",
			3746 => "1110010011101010010001",
			3747 => "1110101011101010010001",
			3748 => "0001000110110010101000",
			3749 => "0000011011101001110100",
			3750 => "0000011001111001000000",
			3751 => "0011101101111000100000",
			3752 => "0010010111100100010000",
			3753 => "0000111101111000001000",
			3754 => "0010010110101000000100",
			3755 => "0000000011110000010101",
			3756 => "0000000011110000010101",
			3757 => "0000100110010000000100",
			3758 => "0000000011110000010101",
			3759 => "0000000011110000010101",
			3760 => "0000101110101000001000",
			3761 => "0010000101000100000100",
			3762 => "0000000011110000010101",
			3763 => "1111111011110000010101",
			3764 => "0010101000100100000100",
			3765 => "0000001011110000010101",
			3766 => "0000000011110000010101",
			3767 => "0010111100001000010000",
			3768 => "0001111011000100001000",
			3769 => "0011011100101100000100",
			3770 => "0000001011110000010101",
			3771 => "1111111011110000010101",
			3772 => "0001101100011000000100",
			3773 => "0000010011110000010101",
			3774 => "0000000011110000010101",
			3775 => "0000011100110100001000",
			3776 => "0011110001000000000100",
			3777 => "1111111011110000010101",
			3778 => "0000000011110000010101",
			3779 => "0000100010000000000100",
			3780 => "0000000011110000010101",
			3781 => "0000000011110000010101",
			3782 => "0011101010111000011000",
			3783 => "0010001011010100001100",
			3784 => "0001111000111000000100",
			3785 => "0000001011110000010101",
			3786 => "0011100000001100000100",
			3787 => "0000000011110000010101",
			3788 => "1111111011110000010101",
			3789 => "0010111101100000000100",
			3790 => "0000000011110000010101",
			3791 => "0001101010011000000100",
			3792 => "0000001011110000010101",
			3793 => "0000001011110000010101",
			3794 => "0001111101100000010000",
			3795 => "0000010110101000001000",
			3796 => "0011000000101000000100",
			3797 => "0000001011110000010101",
			3798 => "0000000011110000010101",
			3799 => "0001001110000000000100",
			3800 => "0000000011110000010101",
			3801 => "1111111011110000010101",
			3802 => "0010001010110000000100",
			3803 => "1111111011110000010101",
			3804 => "0011010000011100000100",
			3805 => "0000000011110000010101",
			3806 => "0000001011110000010101",
			3807 => "0010000110001000010100",
			3808 => "0011001011011100010000",
			3809 => "0001001000001000000100",
			3810 => "1111111011110000010101",
			3811 => "0001001000001000001000",
			3812 => "0010001100000100000100",
			3813 => "0000000011110000010101",
			3814 => "0000000011110000010101",
			3815 => "1111111011110000010101",
			3816 => "0000000011110000010101",
			3817 => "0010111000000000000100",
			3818 => "1111111011110000010101",
			3819 => "0001101001111100010000",
			3820 => "0001001011100000001000",
			3821 => "0010101100011100000100",
			3822 => "0000001011110000010101",
			3823 => "0000000011110000010101",
			3824 => "0010100001010100000100",
			3825 => "1111111011110000010101",
			3826 => "0000001011110000010101",
			3827 => "0011100011010100001000",
			3828 => "0001001110111000000100",
			3829 => "0000000011110000010101",
			3830 => "0000001011110000010101",
			3831 => "0000000011110000010101",
			3832 => "0001101011001100000100",
			3833 => "1111111011110000010101",
			3834 => "0000100010000100001000",
			3835 => "0000011110011100000100",
			3836 => "0000000011110000010101",
			3837 => "0000001011110000010101",
			3838 => "0010101100000100001100",
			3839 => "0010001111000100000100",
			3840 => "1111111011110000010101",
			3841 => "0001000101100000000100",
			3842 => "0000001011110000010101",
			3843 => "0000000011110000010101",
			3844 => "1111111011110000010101",
			3845 => "0011000000001110010000",
			3846 => "0001000110110001111000",
			3847 => "0011101000111100111100",
			3848 => "0010010110101000011100",
			3849 => "0010110100000000010000",
			3850 => "0011011100101100001000",
			3851 => "0000111001110000000100",
			3852 => "0000000011110110011001",
			3853 => "0000000011110110011001",
			3854 => "0000100111111100000100",
			3855 => "0000000011110110011001",
			3856 => "0000001011110110011001",
			3857 => "0010101100011100001000",
			3858 => "0000100101110000000100",
			3859 => "0000000011110110011001",
			3860 => "1111110011110110011001",
			3861 => "0000001011110110011001",
			3862 => "0000011100110100010000",
			3863 => "0011101100001000001000",
			3864 => "0001010110000100000100",
			3865 => "0000000011110110011001",
			3866 => "0000001011110110011001",
			3867 => "0011111011110100000100",
			3868 => "0000000011110110011001",
			3869 => "0000001011110110011001",
			3870 => "0010010111100100001000",
			3871 => "0010111100001000000100",
			3872 => "0000000011110110011001",
			3873 => "0000000011110110011001",
			3874 => "0011110101100100000100",
			3875 => "0000000011110110011001",
			3876 => "0000001011110110011001",
			3877 => "0011110010001000011100",
			3878 => "0010011101101000010000",
			3879 => "0010110000101000001000",
			3880 => "0011000111111000000100",
			3881 => "0000010011110110011001",
			3882 => "0000000011110110011001",
			3883 => "0010000001010100000100",
			3884 => "1111111011110110011001",
			3885 => "1111111011110110011001",
			3886 => "0001011101111000000100",
			3887 => "1111111011110110011001",
			3888 => "0011100101101100000100",
			3889 => "0000000011110110011001",
			3890 => "1111111011110110011001",
			3891 => "0010011101101000010000",
			3892 => "0000100010000000001000",
			3893 => "0011100101101100000100",
			3894 => "0000000011110110011001",
			3895 => "1111111011110110011001",
			3896 => "0001011010111100000100",
			3897 => "0000000011110110011001",
			3898 => "1111111011110110011001",
			3899 => "0011101101111000001000",
			3900 => "0011011101111000000100",
			3901 => "1111111011110110011001",
			3902 => "0000000011110110011001",
			3903 => "0010011111001100000100",
			3904 => "0000000011110110011001",
			3905 => "0000000011110110011001",
			3906 => "0010110100011000010100",
			3907 => "0000011100100000000100",
			3908 => "1111111011110110011001",
			3909 => "0011111001001000000100",
			3910 => "0000000011110110011001",
			3911 => "0000101010001000000100",
			3912 => "1111111011110110011001",
			3913 => "0000101001100000000100",
			3914 => "0000001011110110011001",
			3915 => "1111111011110110011001",
			3916 => "0000001011110110011001",
			3917 => "0010001001101000001000",
			3918 => "0011101010001100000100",
			3919 => "0000001011110110011001",
			3920 => "1111111011110110011001",
			3921 => "0001000011111000101000",
			3922 => "0011101100111000010100",
			3923 => "0000101011110000001100",
			3924 => "0010011011001100001000",
			3925 => "0001001101110100000100",
			3926 => "0000001011110110011001",
			3927 => "0000000011110110011001",
			3928 => "1111111011110110011001",
			3929 => "0000100101000000000100",
			3930 => "0000001011110110011001",
			3931 => "0000000011110110011001",
			3932 => "0011001011011100001100",
			3933 => "0010000110001000000100",
			3934 => "1111111011110110011001",
			3935 => "0000000000111000000100",
			3936 => "0000001011110110011001",
			3937 => "1111111011110110011001",
			3938 => "0000011100011000000100",
			3939 => "1111111011110110011001",
			3940 => "0000001011110110011001",
			3941 => "1111111011110110011001",
			3942 => "0001010100011010101100",
			3943 => "0010101001000101011100",
			3944 => "0010110100010100011100",
			3945 => "0000001111000100001000",
			3946 => "0011101010000000000100",
			3947 => "1111110011111101111101",
			3948 => "1111111011111101111101",
			3949 => "0001001100001100000100",
			3950 => "0000001011111101111101",
			3951 => "0011100011010000001000",
			3952 => "0010101000010100000100",
			3953 => "1111111011111101111101",
			3954 => "0000000011111101111101",
			3955 => "0010001001101000000100",
			3956 => "1111101011111101111101",
			3957 => "1111111011111101111101",
			3958 => "0000100100101000100000",
			3959 => "0001001100001100010000",
			3960 => "0011100000110000001000",
			3961 => "0001000101000000000100",
			3962 => "0000001011111101111101",
			3963 => "0000000011111101111101",
			3964 => "0010011001111000000100",
			3965 => "1111111011111101111101",
			3966 => "0000000011111101111101",
			3967 => "0011111011011100001000",
			3968 => "0000101001010000000100",
			3969 => "0000000011111101111101",
			3970 => "1111111011111101111101",
			3971 => "0000101111010000000100",
			3972 => "0000000011111101111101",
			3973 => "0000001011111101111101",
			3974 => "0010001001101000010000",
			3975 => "0010101000010100001000",
			3976 => "0001001110000000000100",
			3977 => "0000000011111101111101",
			3978 => "0000001011111101111101",
			3979 => "0000100011001000000100",
			3980 => "1111111011111101111101",
			3981 => "0000001011111101111101",
			3982 => "0001101101111100001000",
			3983 => "0001010110000100000100",
			3984 => "0000001011111101111101",
			3985 => "0000000011111101111101",
			3986 => "0001111100001000000100",
			3987 => "0000010011111101111101",
			3988 => "0000001011111101111101",
			3989 => "0001000011001100011000",
			3990 => "0000000000110000010000",
			3991 => "0000001111000100000100",
			3992 => "0000001011111101111101",
			3993 => "0000010110000000000100",
			3994 => "0000001011111101111101",
			3995 => "0001011101010100000100",
			3996 => "0000000011111101111101",
			3997 => "0000000011111101111101",
			3998 => "0000101001011100000100",
			3999 => "0000010011111101111101",
			4000 => "0000001011111101111101",
			4001 => "0001100001111000011000",
			4002 => "0001111011000100010000",
			4003 => "0001110100010100001000",
			4004 => "0010000110001000000100",
			4005 => "0000001011111101111101",
			4006 => "1111111011111101111101",
			4007 => "0011111001110100000100",
			4008 => "0000000011111101111101",
			4009 => "1111110011111101111101",
			4010 => "0001010011011100000100",
			4011 => "1111111011111101111101",
			4012 => "0000001011111101111101",
			4013 => "0010100001010000010000",
			4014 => "0010010111100100001000",
			4015 => "0011101100001000000100",
			4016 => "0000000011111101111101",
			4017 => "0000000011111101111101",
			4018 => "0011001000111000000100",
			4019 => "0000001011111101111101",
			4020 => "1111111011111101111101",
			4021 => "0001001001001100001000",
			4022 => "0010011011101000000100",
			4023 => "0000000011111101111101",
			4024 => "0000000011111101111101",
			4025 => "0011001110111100000100",
			4026 => "0000000011111101111101",
			4027 => "0000000011111101111101",
			4028 => "0010000001010100011000",
			4029 => "0001011000000000010100",
			4030 => "0001111101100000001100",
			4031 => "0001101101111100001000",
			4032 => "0011001000111000000100",
			4033 => "0000000011111101111101",
			4034 => "0000000011111101111101",
			4035 => "1111111011111101111101",
			4036 => "0011111010111000000100",
			4037 => "0000000011111101111101",
			4038 => "0000001011111101111101",
			4039 => "1111111011111101111101",
			4040 => "0001000000000000101100",
			4041 => "0010110110000100010000",
			4042 => "0000000010111100000100",
			4043 => "0000001011111101111101",
			4044 => "0010011111001100000100",
			4045 => "1111110011111101111101",
			4046 => "0000101100000000000100",
			4047 => "0000000011111101111101",
			4048 => "1111111011111101111101",
			4049 => "0011100001011100001100",
			4050 => "0010000001010100000100",
			4051 => "0000010011111101111101",
			4052 => "0010101100000100000100",
			4053 => "0000000011111101111101",
			4054 => "0000001011111101111101",
			4055 => "0001101001111100001000",
			4056 => "0011001011011100000100",
			4057 => "1111111011111101111101",
			4058 => "0000000011111101111101",
			4059 => "0011110000010100000100",
			4060 => "0000000011111101111101",
			4061 => "0000000011111101111101",
			4062 => "1111111011111101111101",
			4063 => "0010011001111010001000",
			4064 => "0001011101100001000100",
			4065 => "0001010011011100111100",
			4066 => "0000101001010000011100",
			4067 => "0000111100001000010000",
			4068 => "0001000000010100001000",
			4069 => "0010001100000100000100",
			4070 => "1111111100000110101001",
			4071 => "0000000100000110101001",
			4072 => "0010101010110000000100",
			4073 => "1111111100000110101001",
			4074 => "0000000100000110101001",
			4075 => "0010001011010100001000",
			4076 => "0000110100000000000100",
			4077 => "0000001100000110101001",
			4078 => "1111111100000110101001",
			4079 => "1111111100000110101001",
			4080 => "0010101010110000010000",
			4081 => "0010101010110000001000",
			4082 => "0011011001110000000100",
			4083 => "1111111100000110101001",
			4084 => "0000000100000110101001",
			4085 => "0001111110111100000100",
			4086 => "0000000100000110101001",
			4087 => "0000001100000110101001",
			4088 => "0001101101111100001000",
			4089 => "0000101110010000000100",
			4090 => "0000000100000110101001",
			4091 => "1111111100000110101001",
			4092 => "0000101110010000000100",
			4093 => "0000000100000110101001",
			4094 => "0000001100000110101001",
			4095 => "0001001011100000000100",
			4096 => "0000001100000110101001",
			4097 => "0000000100000110101001",
			4098 => "0001101101111100100100",
			4099 => "0011011101100000001100",
			4100 => "0011000100010100001000",
			4101 => "0001000101010100000100",
			4102 => "1111111100000110101001",
			4103 => "0000001100000110101001",
			4104 => "1111111100000110101001",
			4105 => "0000000011010000001100",
			4106 => "0000111100001000000100",
			4107 => "0000001100000110101001",
			4108 => "0000101110101000000100",
			4109 => "1111111100000110101001",
			4110 => "0000000100000110101001",
			4111 => "0000101100010100001000",
			4112 => "0010011100110100000100",
			4113 => "0000000100000110101001",
			4114 => "0000001100000110101001",
			4115 => "0000000100000110101001",
			4116 => "0011100000111000010100",
			4117 => "0011100011111100010000",
			4118 => "0010110100010100001000",
			4119 => "0000110100010100000100",
			4120 => "0000000100000110101001",
			4121 => "1111111100000110101001",
			4122 => "0001101101111100000100",
			4123 => "0000001100000110101001",
			4124 => "0000000100000110101001",
			4125 => "0000000100000110101001",
			4126 => "0011100111111000001000",
			4127 => "0000101010001000000100",
			4128 => "1111111100000110101001",
			4129 => "1111111100000110101001",
			4130 => "0000000100000110101001",
			4131 => "0000110101101101001100",
			4132 => "0000110101101100110100",
			4133 => "0000111100110000100000",
			4134 => "0000111100110000010000",
			4135 => "0000111100110000001000",
			4136 => "0011011101111000000100",
			4137 => "0000000100000110101001",
			4138 => "0000001100000110101001",
			4139 => "0011000111111000000100",
			4140 => "0000001100000110101001",
			4141 => "1111111100000110101001",
			4142 => "0010101100011100001000",
			4143 => "0001010110000100000100",
			4144 => "0000000100000110101001",
			4145 => "0000001100000110101001",
			4146 => "0010000010101000000100",
			4147 => "1111111100000110101001",
			4148 => "0000001100000110101001",
			4149 => "0010101001000100001000",
			4150 => "0011011100101100000100",
			4151 => "0000001100000110101001",
			4152 => "0000000100000110101001",
			4153 => "0000101110010000001000",
			4154 => "0011011110001100000100",
			4155 => "1111111100000110101001",
			4156 => "0000000100000110101001",
			4157 => "0000000100000110101001",
			4158 => "0010111100001000001100",
			4159 => "0001111011000100000100",
			4160 => "0000000100000110101001",
			4161 => "0011101011000100000100",
			4162 => "0000001100000110101001",
			4163 => "0000001100000110101001",
			4164 => "0010010111100100000100",
			4165 => "0000000100000110101001",
			4166 => "0001111100001000000100",
			4167 => "0000000100000110101001",
			4168 => "0000001100000110101001",
			4169 => "0011010101101100001100",
			4170 => "0011101001110000001000",
			4171 => "0000101110010000000100",
			4172 => "0000000100000110101001",
			4173 => "1111111100000110101001",
			4174 => "0000000100000110101001",
			4175 => "0000110110000100011100",
			4176 => "0000110101101100010000",
			4177 => "0010101001000100001000",
			4178 => "0010111100001000000100",
			4179 => "1111111100000110101001",
			4180 => "0000001100000110101001",
			4181 => "0000000000110000000100",
			4182 => "1111111100000110101001",
			4183 => "0000000100000110101001",
			4184 => "0011011101111000001000",
			4185 => "0000100100101000000100",
			4186 => "1111111100000110101001",
			4187 => "1111111100000110101001",
			4188 => "0000000100000110101001",
			4189 => "0000110110000100001100",
			4190 => "0010101100011100001000",
			4191 => "0000101001010000000100",
			4192 => "0000000100000110101001",
			4193 => "0000001100000110101001",
			4194 => "1111111100000110101001",
			4195 => "0011000000101000001000",
			4196 => "0011000000101000000100",
			4197 => "0000000100000110101001",
			4198 => "0000000100000110101001",
			4199 => "0001111100001000000100",
			4200 => "0000000100000110101001",
			4201 => "0000000100000110101001",
			4202 => "0000110100000010001100",
			4203 => "0001000011010101000100",
			4204 => "0000000100010100110100",
			4205 => "0000110100000000100000",
			4206 => "0000111100001000010000",
			4207 => "0001100100110100001000",
			4208 => "0011100011111100000100",
			4209 => "0000000100001111001101",
			4210 => "0000000100001111001101",
			4211 => "0010011001111000000100",
			4212 => "1111111100001111001101",
			4213 => "0000000100001111001101",
			4214 => "0001001010110100001000",
			4215 => "0001111011000100000100",
			4216 => "1111111100001111001101",
			4217 => "0000000100001111001101",
			4218 => "0011100011010000000100",
			4219 => "0000000100001111001101",
			4220 => "0000001100001111001101",
			4221 => "0010110100010100001100",
			4222 => "0001001010110100000100",
			4223 => "0000001100001111001101",
			4224 => "0001000000010100000100",
			4225 => "1111111100001111001101",
			4226 => "0000000100001111001101",
			4227 => "0010010110101000000100",
			4228 => "0000001100001111001101",
			4229 => "0000000100001111001101",
			4230 => "0001100100110100000100",
			4231 => "0000001100001111001101",
			4232 => "0011011101100000000100",
			4233 => "1111111100001111001101",
			4234 => "0011011100101100000100",
			4235 => "0000001100001111001101",
			4236 => "0000000100001111001101",
			4237 => "0001000011110100011000",
			4238 => "0000011110100000010100",
			4239 => "0001101101111100000100",
			4240 => "1111111100001111001101",
			4241 => "0000111100001000001000",
			4242 => "0010110100010100000100",
			4243 => "0000000100001111001101",
			4244 => "0000000100001111001101",
			4245 => "0001100100110100000100",
			4246 => "0000000100001111001101",
			4247 => "1111110100001111001101",
			4248 => "0000001100001111001101",
			4249 => "0000010110000000011100",
			4250 => "0011111110110000001100",
			4251 => "0001000110110000000100",
			4252 => "0000001100001111001101",
			4253 => "0001101011001100000100",
			4254 => "0000000100001111001101",
			4255 => "0000000100001111001101",
			4256 => "0010111110111100001000",
			4257 => "0001011000111000000100",
			4258 => "0000000100001111001101",
			4259 => "0000001100001111001101",
			4260 => "0011000100010100000100",
			4261 => "1111111100001111001101",
			4262 => "0000000100001111001101",
			4263 => "0000010110000000001000",
			4264 => "0000001000111000000100",
			4265 => "0000001100001111001101",
			4266 => "0000000100001111001101",
			4267 => "0010110111111000000100",
			4268 => "1111111100001111001101",
			4269 => "0011110101100100000100",
			4270 => "0000000100001111001101",
			4271 => "0000001100001111001101",
			4272 => "0010010010001100011100",
			4273 => "0001100001111000001100",
			4274 => "0011100000110000001000",
			4275 => "0001001101110100000100",
			4276 => "0000001100001111001101",
			4277 => "0000000100001111001101",
			4278 => "0000000100001111001101",
			4279 => "0001101101111100000100",
			4280 => "1111111100001111001101",
			4281 => "0011101010000000001000",
			4282 => "0011110110110100000100",
			4283 => "0000001100001111001101",
			4284 => "0000000100001111001101",
			4285 => "1111111100001111001101",
			4286 => "0011110001011000110000",
			4287 => "0010010110101000010100",
			4288 => "0000011110100000010000",
			4289 => "0011100000110000001000",
			4290 => "0001110100010100000100",
			4291 => "0000000100001111001101",
			4292 => "0000001100001111001101",
			4293 => "0001010101101100000100",
			4294 => "1111111100001111001101",
			4295 => "0000000100001111001101",
			4296 => "1111111100001111001101",
			4297 => "0011011110001100010000",
			4298 => "0011110000011100001000",
			4299 => "0010001001101000000100",
			4300 => "0000001100001111001101",
			4301 => "0000000100001111001101",
			4302 => "0000110011011100000100",
			4303 => "1111111100001111001101",
			4304 => "0000000100001111001101",
			4305 => "0011100000110000000100",
			4306 => "1111111100001111001101",
			4307 => "0001001010110100000100",
			4308 => "0000000100001111001101",
			4309 => "0000001100001111001101",
			4310 => "0010000110001000100000",
			4311 => "0001000011001100010000",
			4312 => "0011100111111000001000",
			4313 => "0011010110000100000100",
			4314 => "1111111100001111001101",
			4315 => "0000000100001111001101",
			4316 => "0001011101111000000100",
			4317 => "0000000100001111001101",
			4318 => "0000000100001111001101",
			4319 => "0011111010010100001000",
			4320 => "0010001001101000000100",
			4321 => "0000001100001111001101",
			4322 => "0000000100001111001101",
			4323 => "0011011100101000000100",
			4324 => "0000001100001111001101",
			4325 => "0000000100001111001101",
			4326 => "0001110111111000001100",
			4327 => "0001011100110000001000",
			4328 => "0001011101100000000100",
			4329 => "0000000100001111001101",
			4330 => "0000001100001111001101",
			4331 => "0000000100001111001101",
			4332 => "0000000100010100001000",
			4333 => "0010000111000100000100",
			4334 => "0000000100001111001101",
			4335 => "0000000100001111001101",
			4336 => "0001000000010100000100",
			4337 => "0000001100001111001101",
			4338 => "0000000100001111001101",
			4339 => "0000100010110101110000",
			4340 => "0000100001001000100100",
			4341 => "0000001000110000010000",
			4342 => "0010111011000100000100",
			4343 => "1111111100011000100001",
			4344 => "0011000100010100001000",
			4345 => "0000000110001000000100",
			4346 => "0000000100011000100001",
			4347 => "0000001100011000100001",
			4348 => "1111111100011000100001",
			4349 => "0011001010000000010000",
			4350 => "0001110111111000001000",
			4351 => "0001111010000000000100",
			4352 => "0000000100011000100001",
			4353 => "1111111100011000100001",
			4354 => "0000011100100000000100",
			4355 => "0000000100011000100001",
			4356 => "0000001100011000100001",
			4357 => "0000001100011000100001",
			4358 => "0010110100010100101000",
			4359 => "0001110111111000011100",
			4360 => "0001111110111100001100",
			4361 => "0001100001111000000100",
			4362 => "0000000100011000100001",
			4363 => "0010101100000100000100",
			4364 => "0000001100011000100001",
			4365 => "0000000100011000100001",
			4366 => "0011001010000000001000",
			4367 => "0000101110101100000100",
			4368 => "0000000100011000100001",
			4369 => "0000000100011000100001",
			4370 => "0001100001111000000100",
			4371 => "0000000100011000100001",
			4372 => "1111111100011000100001",
			4373 => "0011110110100100001000",
			4374 => "0000010000011000000100",
			4375 => "0000000100011000100001",
			4376 => "0000001100011000100001",
			4377 => "0000000100011000100001",
			4378 => "0001011100110000010000",
			4379 => "0000100000110100000100",
			4380 => "0000000100011000100001",
			4381 => "0011000100010100001000",
			4382 => "0000001110111100000100",
			4383 => "1111111100011000100001",
			4384 => "1111110100011000100001",
			4385 => "0000000100011000100001",
			4386 => "0000000000111000010000",
			4387 => "0001100111101000001000",
			4388 => "0011111111011100000100",
			4389 => "0000001100011000100001",
			4390 => "0000000100011000100001",
			4391 => "0010010110101000000100",
			4392 => "1111111100011000100001",
			4393 => "0000000100011000100001",
			4394 => "0000001100011000100001",
			4395 => "0000000010111101011000",
			4396 => "0001000110001100110100",
			4397 => "0010100110011000100000",
			4398 => "0010101000010100010000",
			4399 => "0010001001101000001000",
			4400 => "0001001100001100000100",
			4401 => "0000000100011000100001",
			4402 => "1111111100011000100001",
			4403 => "0010111100001000000100",
			4404 => "0000001100011000100001",
			4405 => "0000000100011000100001",
			4406 => "0001001000110100001000",
			4407 => "0000010010001100000100",
			4408 => "0000001100011000100001",
			4409 => "0000000100011000100001",
			4410 => "0011000100000000000100",
			4411 => "1111111100011000100001",
			4412 => "0000000100011000100001",
			4413 => "0001010100011000001000",
			4414 => "0000011001111000000100",
			4415 => "0000000100011000100001",
			4416 => "0000001100011000100001",
			4417 => "0001111101100000000100",
			4418 => "1111111100011000100001",
			4419 => "0010001011010100000100",
			4420 => "1111111100011000100001",
			4421 => "0000001100011000100001",
			4422 => "0000010110000000000100",
			4423 => "1111111100011000100001",
			4424 => "0000000010011000010000",
			4425 => "0010001001101000001000",
			4426 => "0000001111000100000100",
			4427 => "0000000100011000100001",
			4428 => "1111110100011000100001",
			4429 => "0011001001110100000100",
			4430 => "0000000100011000100001",
			4431 => "0000001100011000100001",
			4432 => "0011000100000000001000",
			4433 => "0010111000111100000100",
			4434 => "0000000100011000100001",
			4435 => "0000001100011000100001",
			4436 => "0010001001101000000100",
			4437 => "0000001100011000100001",
			4438 => "1111111100011000100001",
			4439 => "0000111100001000111000",
			4440 => "0001001110111000011000",
			4441 => "0010111011000100010000",
			4442 => "0001110100010100001000",
			4443 => "0001100001111000000100",
			4444 => "0000000100011000100001",
			4445 => "0000001100011000100001",
			4446 => "0001001101001000000100",
			4447 => "0000001100011000100001",
			4448 => "0000000100011000100001",
			4449 => "0010110000101000000100",
			4450 => "0000001100011000100001",
			4451 => "0000000100011000100001",
			4452 => "0000000111111000010000",
			4453 => "0011001010000000001000",
			4454 => "0010110111111000000100",
			4455 => "1111111100011000100001",
			4456 => "0000001100011000100001",
			4457 => "0001100001111000000100",
			4458 => "0000000100011000100001",
			4459 => "1111111100011000100001",
			4460 => "0011000111111000001000",
			4461 => "0011000111111000000100",
			4462 => "0000000100011000100001",
			4463 => "1111111100011000100001",
			4464 => "0011000111111000000100",
			4465 => "0000001100011000100001",
			4466 => "0000000100011000100001",
			4467 => "0010001001101000011000",
			4468 => "0000111101111000001100",
			4469 => "0011000000101000001000",
			4470 => "0010111011000100000100",
			4471 => "0000000100011000100001",
			4472 => "1111111100011000100001",
			4473 => "0000001100011000100001",
			4474 => "0000110100011000001000",
			4475 => "0000000010111100000100",
			4476 => "1111111100011000100001",
			4477 => "1111111100011000100001",
			4478 => "0000000100011000100001",
			4479 => "0010001001101000000100",
			4480 => "0000001100011000100001",
			4481 => "0011000111111000001000",
			4482 => "0011001010000000000100",
			4483 => "0000000100011000100001",
			4484 => "0000000100011000100001",
			4485 => "0011000111111000000100",
			4486 => "0000000100011000100001",
			4487 => "0000000100011000100001",
			4488 => "0001110100010110010000",
			4489 => "0000110000101000111000",
			4490 => "0010001100000100010000",
			4491 => "0000100010110100001000",
			4492 => "0011000111111000000100",
			4493 => "1111111100100010101101",
			4494 => "0000001100100010101101",
			4495 => "0011101101010000000100",
			4496 => "0000000100100010101101",
			4497 => "1111110100100010101101",
			4498 => "0001000000010100010000",
			4499 => "0001101101111100001100",
			4500 => "0011000000110000000100",
			4501 => "0000000100100010101101",
			4502 => "0000010110000000000100",
			4503 => "0000000100100010101101",
			4504 => "0000001100100010101101",
			4505 => "0000000100100010101101",
			4506 => "0000001110111100001000",
			4507 => "0000111110111100000100",
			4508 => "0000000100100010101101",
			4509 => "1111110100100010101101",
			4510 => "0010010010001100001000",
			4511 => "0000101101000100000100",
			4512 => "0000001100100010101101",
			4513 => "0000000100100010101101",
			4514 => "0011101101010000000100",
			4515 => "0000000100100010101101",
			4516 => "0000001100100010101101",
			4517 => "0011000111111000101000",
			4518 => "0011000000110000010000",
			4519 => "0001000011010100001100",
			4520 => "0000111101100000001000",
			4521 => "0001110111111000000100",
			4522 => "0000000100100010101101",
			4523 => "0000001100100010101101",
			4524 => "1111111100100010101101",
			4525 => "1111111100100010101101",
			4526 => "0000101110101000001000",
			4527 => "0010001001101000000100",
			4528 => "0000000100100010101101",
			4529 => "1111110100100010101101",
			4530 => "0010100110011000001000",
			4531 => "0000000010111100000100",
			4532 => "1111111100100010101101",
			4533 => "0000000100100010101101",
			4534 => "0010000111000100000100",
			4535 => "1111111100100010101101",
			4536 => "0000000100100010101101",
			4537 => "0001110111111000011000",
			4538 => "0000111100001000001000",
			4539 => "0000101001010000000100",
			4540 => "0000001100100010101101",
			4541 => "0000000100100010101101",
			4542 => "0011110111110000001000",
			4543 => "0011000100010100000100",
			4544 => "1111110100100010101101",
			4545 => "1111111100100010101101",
			4546 => "0000101100010100000100",
			4547 => "0000001100100010101101",
			4548 => "0000000100100010101101",
			4549 => "0011101110111100001100",
			4550 => "0011110000011100000100",
			4551 => "0000000100100010101101",
			4552 => "0000110100000000000100",
			4553 => "0000001100100010101101",
			4554 => "0000001100100010101101",
			4555 => "0001110111111000000100",
			4556 => "0000001100100010101101",
			4557 => "0011011110001100000100",
			4558 => "0000000100100010101101",
			4559 => "0000000100100010101101",
			4560 => "0001110000101001001100",
			4561 => "0001110000101000111000",
			4562 => "0011110001101000011100",
			4563 => "0010101000100100001100",
			4564 => "0001101011111100000100",
			4565 => "1111111100100010101101",
			4566 => "0011000100010100000100",
			4567 => "0000001100100010101101",
			4568 => "0000000100100010101101",
			4569 => "0011100010011000001000",
			4570 => "0011011100110000000100",
			4571 => "0000000100100010101101",
			4572 => "0000001100100010101101",
			4573 => "0011110110100100000100",
			4574 => "1111110100100010101101",
			4575 => "1111111100100010101101",
			4576 => "0011000000101000010000",
			4577 => "0001111011000100001000",
			4578 => "0001110100010100000100",
			4579 => "0000000100100010101101",
			4580 => "0000000100100010101101",
			4581 => "0010100110011100000100",
			4582 => "0000000100100010101101",
			4583 => "1111111100100010101101",
			4584 => "0000011100110100000100",
			4585 => "0000000100100010101101",
			4586 => "0010010111100100000100",
			4587 => "1111111100100010101101",
			4588 => "0000000100100010101101",
			4589 => "0010010111100100010000",
			4590 => "0011011100101100001000",
			4591 => "0011000100010100000100",
			4592 => "0000001100100010101101",
			4593 => "0000000100100010101101",
			4594 => "0000111100110000000100",
			4595 => "0000000100100010101101",
			4596 => "0000001100100010101101",
			4597 => "0000001100100010101101",
			4598 => "0001111100001000110000",
			4599 => "0010101100011100011100",
			4600 => "0000001110111100010000",
			4601 => "0010010110101000001000",
			4602 => "0000011110100000000100",
			4603 => "0000000100100010101101",
			4604 => "1111111100100010101101",
			4605 => "0010100001010000000100",
			4606 => "0000000100100010101101",
			4607 => "1111111100100010101101",
			4608 => "0011011101111000001000",
			4609 => "0011010110000100000100",
			4610 => "0000000100100010101101",
			4611 => "0000001100100010101101",
			4612 => "0000000100100010101101",
			4613 => "0010100110011100001000",
			4614 => "0010000010101000000100",
			4615 => "1111110100100010101101",
			4616 => "1111111100100010101101",
			4617 => "0011000100010100001000",
			4618 => "0011000100010100000100",
			4619 => "0000000100100010101101",
			4620 => "1111111100100010101101",
			4621 => "0000000100100010101101",
			4622 => "0001111100001000100000",
			4623 => "0001111100001000010000",
			4624 => "0000101100010100001000",
			4625 => "0001111100001000000100",
			4626 => "0000000100100010101101",
			4627 => "0000000100100010101101",
			4628 => "0001101010011000000100",
			4629 => "0000001100100010101101",
			4630 => "0000000100100010101101",
			4631 => "0001001100001100001000",
			4632 => "0010001001101000000100",
			4633 => "0000001100100010101101",
			4634 => "0000010100100010101101",
			4635 => "0000000011010000000100",
			4636 => "0000000100100010101101",
			4637 => "0000001100100010101101",
			4638 => "0001110100000000001100",
			4639 => "0001000010100100001000",
			4640 => "0010100110011100000100",
			4641 => "0000000100100010101101",
			4642 => "1111110100100010101101",
			4643 => "0000001100100010101101",
			4644 => "0010011101101000001000",
			4645 => "0011101100101100000100",
			4646 => "0000000100100010101101",
			4647 => "0000000100100010101101",
			4648 => "0001110100000000000100",
			4649 => "0000001100100010101101",
			4650 => "0000000100100010101101",
			4651 => "0001000110111100000100",
			4652 => "1111111100101000010001",
			4653 => "0001110000101001011000",
			4654 => "0001110100010100110000",
			4655 => "0001110100010100010000",
			4656 => "0000011100110100001100",
			4657 => "0010010111100100001000",
			4658 => "0001011100101100000100",
			4659 => "0000000100101000010001",
			4660 => "0000001100101000010001",
			4661 => "0000001100101000010001",
			4662 => "1111111100101000010001",
			4663 => "0010110100010100010000",
			4664 => "0011111010111000001000",
			4665 => "0011000111111000000100",
			4666 => "0000000100101000010001",
			4667 => "1111110100101000010001",
			4668 => "0010110100010100000100",
			4669 => "0000000100101000010001",
			4670 => "0000001100101000010001",
			4671 => "0010111011000100001000",
			4672 => "0011000111111000000100",
			4673 => "1111111100101000010001",
			4674 => "0000000100101000010001",
			4675 => "0011111011110100000100",
			4676 => "0000000100101000010001",
			4677 => "0000001100101000010001",
			4678 => "0001010011011100010100",
			4679 => "0001001001001100001000",
			4680 => "0001111011000100000100",
			4681 => "1111111100101000010001",
			4682 => "0000001100101000010001",
			4683 => "0000100010011100001000",
			4684 => "0000111011000100000100",
			4685 => "1111111100101000010001",
			4686 => "1111110100101000010001",
			4687 => "0000000100101000010001",
			4688 => "0000100010000100010000",
			4689 => "0001001111100000001000",
			4690 => "0000010010001100000100",
			4691 => "0000000100101000010001",
			4692 => "0000001100101000010001",
			4693 => "0011010110000100000100",
			4694 => "0000000100101000010001",
			4695 => "0000001100101000010001",
			4696 => "1111111100101000010001",
			4697 => "0001110000101000011000",
			4698 => "0001100111101000000100",
			4699 => "1111111100101000010001",
			4700 => "0001011110001100010000",
			4701 => "0001010110000100001000",
			4702 => "0011000100010100000100",
			4703 => "0000001100101000010001",
			4704 => "0000000100101000010001",
			4705 => "0001101101111100000100",
			4706 => "0000000100101000010001",
			4707 => "0000001100101000010001",
			4708 => "0000000100101000010001",
			4709 => "0010100111110100100000",
			4710 => "0011000100000000010000",
			4711 => "0000111010111100001000",
			4712 => "0000110000001100000100",
			4713 => "0000001100101000010001",
			4714 => "1111111100101000010001",
			4715 => "0001101101111100000100",
			4716 => "0000001100101000010001",
			4717 => "0000000100101000010001",
			4718 => "0001001111101000001000",
			4719 => "0001001011101100000100",
			4720 => "0000000100101000010001",
			4721 => "1111111100101000010001",
			4722 => "0000100111011000000100",
			4723 => "0000001100101000010001",
			4724 => "0000000100101000010001",
			4725 => "0001000100001100010000",
			4726 => "0011000111111000001000",
			4727 => "0001001000001000000100",
			4728 => "0000000100101000010001",
			4729 => "0000001100101000010001",
			4730 => "0010011011101000000100",
			4731 => "0000000100101000010001",
			4732 => "0000000100101000010001",
			4733 => "0010001111001000001000",
			4734 => "0001001111100000000100",
			4735 => "1111110100101000010001",
			4736 => "0000000100101000010001",
			4737 => "0010000010101000000100",
			4738 => "0000000100101000010001",
			4739 => "0000000100101000010001",
			4740 => "0010010110101010110000",
			4741 => "0000110011011101001100",
			4742 => "0011110110110100100100",
			4743 => "0000111001110000100000",
			4744 => "0011100011010000010000",
			4745 => "0011000100010100001000",
			4746 => "0011001010000000000100",
			4747 => "0000000100110010100101",
			4748 => "0000000100110010100101",
			4749 => "0000110100010100000100",
			4750 => "0000000100110010100101",
			4751 => "0000001100110010100101",
			4752 => "0001101101111100001000",
			4753 => "0010011001111000000100",
			4754 => "0000000100110010100101",
			4755 => "0000000100110010100101",
			4756 => "0001100100110100000100",
			4757 => "1111111100110010100101",
			4758 => "0000000100110010100101",
			4759 => "0000001100110010100101",
			4760 => "0010011001111000011000",
			4761 => "0001110100010100001100",
			4762 => "0001011101100000001000",
			4763 => "0000111001110000000100",
			4764 => "0000000100110010100101",
			4765 => "0000000100110010100101",
			4766 => "1111111100110010100101",
			4767 => "0010000110001000000100",
			4768 => "0000000100110010100101",
			4769 => "0000001000011000000100",
			4770 => "0000001100110010100101",
			4771 => "0000000100110010100101",
			4772 => "0001001010110100000100",
			4773 => "0000000100110010100101",
			4774 => "0010010110101000001000",
			4775 => "0001111100001000000100",
			4776 => "0000001100110010100101",
			4777 => "0000000100110010100101",
			4778 => "0000000100110010100101",
			4779 => "0000100101110000101000",
			4780 => "0001010101101100010000",
			4781 => "0011011100110000000100",
			4782 => "0000000100110010100101",
			4783 => "0000101101000100000100",
			4784 => "0000001100110010100101",
			4785 => "0010011001111000000100",
			4786 => "0000000100110010100101",
			4787 => "1111111100110010100101",
			4788 => "0001010101101100001000",
			4789 => "0011111011011100000100",
			4790 => "0000001100110010100101",
			4791 => "0000000100110010100101",
			4792 => "0000000000111000001000",
			4793 => "0001000101000000000100",
			4794 => "1111111100110010100101",
			4795 => "0000000100110010100101",
			4796 => "0011000100010100000100",
			4797 => "0000000100110010100101",
			4798 => "1111111100110010100101",
			4799 => "0001001001001100011100",
			4800 => "0000110101101100001100",
			4801 => "0001010101101100001000",
			4802 => "0000001010000000000100",
			4803 => "0000000100110010100101",
			4804 => "0000001100110010100101",
			4805 => "0000001100110010100101",
			4806 => "0011110001001000001000",
			4807 => "0001001101001000000100",
			4808 => "0000000100110010100101",
			4809 => "1111111100110010100101",
			4810 => "0011100101101100000100",
			4811 => "0000001100110010100101",
			4812 => "0000000100110010100101",
			4813 => "0011000100010100010000",
			4814 => "0011010110000100001000",
			4815 => "0001011100110000000100",
			4816 => "0000000100110010100101",
			4817 => "1111111100110010100101",
			4818 => "0010111100001000000100",
			4819 => "0000001100110010100101",
			4820 => "0000000100110010100101",
			4821 => "0010110000101000001000",
			4822 => "0001110100010100000100",
			4823 => "1111111100110010100101",
			4824 => "0000001100110010100101",
			4825 => "0001101101111100000100",
			4826 => "0000001100110010100101",
			4827 => "1111111100110010100101",
			4828 => "0000110101101101100000",
			4829 => "0010111100001000100100",
			4830 => "0001100001111000010000",
			4831 => "0001001011110000000100",
			4832 => "1111111100110010100101",
			4833 => "0000111100110000001000",
			4834 => "0011110000011100000100",
			4835 => "0000001100110010100101",
			4836 => "0000000100110010100101",
			4837 => "0000001100110010100101",
			4838 => "0010001001101000000100",
			4839 => "1111111100110010100101",
			4840 => "0000001010000000001000",
			4841 => "0000000000110000000100",
			4842 => "0000000100110010100101",
			4843 => "1111111100110010100101",
			4844 => "0011000000101000000100",
			4845 => "0000000100110010100101",
			4846 => "0000000100110010100101",
			4847 => "0011111011011100100000",
			4848 => "0000111101100000010000",
			4849 => "0011100000111000001000",
			4850 => "0001101100011000000100",
			4851 => "0000000100110010100101",
			4852 => "1111111100110010100101",
			4853 => "0011100111111000000100",
			4854 => "0000001100110010100101",
			4855 => "0000000100110010100101",
			4856 => "0010010111100100001000",
			4857 => "0011000100010100000100",
			4858 => "1111111100110010100101",
			4859 => "0000000100110010100101",
			4860 => "0001001010110100000100",
			4861 => "0000000100110010100101",
			4862 => "0000001100110010100101",
			4863 => "0011110010001000001100",
			4864 => "0010111100001000000100",
			4865 => "0000001100110010100101",
			4866 => "0011101011000100000100",
			4867 => "0000001100110010100101",
			4868 => "0000010100110010100101",
			4869 => "0011110101110100001000",
			4870 => "0011110100010000000100",
			4871 => "0000000100110010100101",
			4872 => "1111111100110010100101",
			4873 => "0001101010011000000100",
			4874 => "0000001100110010100101",
			4875 => "0000000100110010100101",
			4876 => "0000110110000100010000",
			4877 => "0000100100101000001000",
			4878 => "0011011110001100000100",
			4879 => "0000001100110010100101",
			4880 => "1111111100110010100101",
			4881 => "0010000111000100000100",
			4882 => "1111111100110010100101",
			4883 => "0000000100110010100101",
			4884 => "0000110110000100001100",
			4885 => "0010000111000100001000",
			4886 => "0001011100101100000100",
			4887 => "0000001100110010100101",
			4888 => "0000001100110010100101",
			4889 => "0000000100110010100101",
			4890 => "0000100101110000010000",
			4891 => "0010000110001000001000",
			4892 => "0011101011000100000100",
			4893 => "0000001100110010100101",
			4894 => "0000000100110010100101",
			4895 => "0000111110001100000100",
			4896 => "1111111100110010100101",
			4897 => "0000000100110010100101",
			4898 => "0001111100001000001000",
			4899 => "0000110000001100000100",
			4900 => "0000000100110010100101",
			4901 => "0000000100110010100101",
			4902 => "0010111100001000000100",
			4903 => "1111111100110010100101",
			4904 => "0000000100110010100101",
			4905 => "0010010010001110010100",
			4906 => "0011101111000101011100",
			4907 => "0010100101000100101100",
			4908 => "0010000111000100010100",
			4909 => "0000010110000000010000",
			4910 => "0011001010000000001000",
			4911 => "0001100001111000000100",
			4912 => "1111111100111101011001",
			4913 => "0000000100111101011001",
			4914 => "0001110111111000000100",
			4915 => "1111111100111101011001",
			4916 => "0000001100111101011001",
			4917 => "1111111100111101011001",
			4918 => "0010011110100000001100",
			4919 => "0011101011010100001000",
			4920 => "0000101111010000000100",
			4921 => "0000001100111101011001",
			4922 => "0000000100111101011001",
			4923 => "1111111100111101011001",
			4924 => "0000101111010000001000",
			4925 => "0000010000011000000100",
			4926 => "0000000100111101011001",
			4927 => "0000001100111101011001",
			4928 => "0000000100111101011001",
			4929 => "0001010011011100011100",
			4930 => "0001110111111000001100",
			4931 => "0000101010010100000100",
			4932 => "0000001100111101011001",
			4933 => "0011111010001100000100",
			4934 => "1111111100111101011001",
			4935 => "0000000100111101011001",
			4936 => "0001101101111100001000",
			4937 => "0001100001111000000100",
			4938 => "1111111100111101011001",
			4939 => "1111110100111101011001",
			4940 => "0011000111111000000100",
			4941 => "0000001100111101011001",
			4942 => "0000000100111101011001",
			4943 => "0011011101100000001000",
			4944 => "0011010011011100000100",
			4945 => "1111111100111101011001",
			4946 => "1111110100111101011001",
			4947 => "0011000100010100000100",
			4948 => "0000001100111101011001",
			4949 => "0000101110101000000100",
			4950 => "0000000100111101011001",
			4951 => "1111111100111101011001",
			4952 => "0010001111001000100000",
			4953 => "0010001011010100010000",
			4954 => "0001110100010100001100",
			4955 => "0010101000100100000100",
			4956 => "0000000100111101011001",
			4957 => "0001011000111000000100",
			4958 => "0000000100111101011001",
			4959 => "1111110100111101011001",
			4960 => "0000001100111101011001",
			4961 => "0000010000011000000100",
			4962 => "1111111100111101011001",
			4963 => "0010110111111000000100",
			4964 => "0000000100111101011001",
			4965 => "0011110111010000000100",
			4966 => "0000000100111101011001",
			4967 => "0000001100111101011001",
			4968 => "0011100010011000000100",
			4969 => "1111111100111101011001",
			4970 => "0010010010001100010000",
			4971 => "0010000010101000001000",
			4972 => "0010101010110000000100",
			4973 => "0000000100111101011001",
			4974 => "1111111100111101011001",
			4975 => "0001000001101100000100",
			4976 => "0000000100111101011001",
			4977 => "1111111100111101011001",
			4978 => "0000000100111101011001",
			4979 => "0011000111111001101000",
			4980 => "0001111011000100111100",
			4981 => "0001100001111000011100",
			4982 => "0001010011011100001100",
			4983 => "0011000111111000001000",
			4984 => "0010000110001000000100",
			4985 => "1111111100111101011001",
			4986 => "0000001100111101011001",
			4987 => "1111110100111101011001",
			4988 => "0011100100010100001000",
			4989 => "0001010101101100000100",
			4990 => "0000000100111101011001",
			4991 => "1111111100111101011001",
			4992 => "0001100001111000000100",
			4993 => "0000000100111101011001",
			4994 => "1111111100111101011001",
			4995 => "0011000111111000010000",
			4996 => "0010101001000100001000",
			4997 => "0000011110100000000100",
			4998 => "0000001100111101011001",
			4999 => "0000000100111101011001",
			5000 => "0011001010000000000100",
			5001 => "0000000100111101011001",
			5002 => "1111111100111101011001",
			5003 => "0001101101111100001000",
			5004 => "0001110100010100000100",
			5005 => "0000001100111101011001",
			5006 => "0000000100111101011001",
			5007 => "0001101101111100000100",
			5008 => "0000000100111101011001",
			5009 => "0000000100111101011001",
			5010 => "0001111100001000100000",
			5011 => "0001101100011000010000",
			5012 => "0011000111111000001000",
			5013 => "0000011110100000000100",
			5014 => "0000001100111101011001",
			5015 => "0000001100111101011001",
			5016 => "0011000111111000000100",
			5017 => "0000000100111101011001",
			5018 => "0000001100111101011001",
			5019 => "0010101010110000001000",
			5020 => "0001011100101100000100",
			5021 => "1111111100111101011001",
			5022 => "0000000100111101011001",
			5023 => "0000100010011100000100",
			5024 => "1111111100111101011001",
			5025 => "0000001100111101011001",
			5026 => "0010101001000100000100",
			5027 => "0000000100111101011001",
			5028 => "0001000011001100000100",
			5029 => "1111111100111101011001",
			5030 => "0000000100111101011001",
			5031 => "0011000100010100101100",
			5032 => "0001011110001100011100",
			5033 => "0010010110101000010000",
			5034 => "0001010110000100001000",
			5035 => "0001011101100000000100",
			5036 => "0000000100111101011001",
			5037 => "1111111100111101011001",
			5038 => "0000100010011100000100",
			5039 => "0000001100111101011001",
			5040 => "0000000100111101011001",
			5041 => "0001001000011100000100",
			5042 => "0000000100111101011001",
			5043 => "0010110000101000000100",
			5044 => "0000000100111101011001",
			5045 => "1111111100111101011001",
			5046 => "0010111000111100001000",
			5047 => "0010110100000000000100",
			5048 => "0000000100111101011001",
			5049 => "0000010100111101011001",
			5050 => "0010001011010100000100",
			5051 => "0000000100111101011001",
			5052 => "1111111100111101011001",
			5053 => "0011000100010100010100",
			5054 => "0011010101101100000100",
			5055 => "0000001100111101011001",
			5056 => "0010110000101000001000",
			5057 => "0010110000101000000100",
			5058 => "0000000100111101011001",
			5059 => "1111111100111101011001",
			5060 => "0000011100110100000100",
			5061 => "0000001100111101011001",
			5062 => "0000000100111101011001",
			5063 => "0010010110101000010000",
			5064 => "0011100000101000001000",
			5065 => "0010010110101000000100",
			5066 => "0000000100111101011001",
			5067 => "0000000100111101011001",
			5068 => "0010111011000100000100",
			5069 => "0000001100111101011001",
			5070 => "0000000100111101011001",
			5071 => "0011101011000100001000",
			5072 => "0001111100001000000100",
			5073 => "0000001100111101011001",
			5074 => "0000000100111101011001",
			5075 => "0011000100010100000100",
			5076 => "0000001100111101011001",
			5077 => "0000000100111101011001",
			5078 => "0011101100001010111100",
			5079 => "0011110010001001101000",
			5080 => "0001000000010100111000",
			5081 => "0000110100010100011000",
			5082 => "0010001100000100001000",
			5083 => "0010110100010100000100",
			5084 => "1111111101001000111101",
			5085 => "0000001101001000111101",
			5086 => "0010000111000100001000",
			5087 => "0001110100010100000100",
			5088 => "0000001101001000111101",
			5089 => "0000000101001000111101",
			5090 => "0010110100010100000100",
			5091 => "0000001101001000111101",
			5092 => "1111111101001000111101",
			5093 => "0011011110001100010000",
			5094 => "0000111101100000001000",
			5095 => "0000101110101000000100",
			5096 => "0000000101001000111101",
			5097 => "0000000101001000111101",
			5098 => "0010010110101000000100",
			5099 => "1111111101001000111101",
			5100 => "0000000101001000111101",
			5101 => "0001100100110100001000",
			5102 => "0001000001011100000100",
			5103 => "1111111101001000111101",
			5104 => "0000001101001000111101",
			5105 => "0001111100001000000100",
			5106 => "1111111101001000111101",
			5107 => "0000000101001000111101",
			5108 => "0000001011000100011100",
			5109 => "0011011110001100010000",
			5110 => "0010010110101000001000",
			5111 => "0000111000111000000100",
			5112 => "0000000101001000111101",
			5113 => "1111111101001000111101",
			5114 => "0011000100010100000100",
			5115 => "0000000101001000111101",
			5116 => "0000001101001000111101",
			5117 => "0000000111111000000100",
			5118 => "0000000101001000111101",
			5119 => "0011100111111000000100",
			5120 => "1111110101001000111101",
			5121 => "0000000101001000111101",
			5122 => "0001000010100100001000",
			5123 => "0011111011011100000100",
			5124 => "0000001101001000111101",
			5125 => "0000000101001000111101",
			5126 => "0011101110111100001000",
			5127 => "0001110111111000000100",
			5128 => "1111111101001000111101",
			5129 => "0000000101001000111101",
			5130 => "1111111101001000111101",
			5131 => "0011100000101000111000",
			5132 => "0011101011000100100000",
			5133 => "0001111011000100010000",
			5134 => "0000011110100000001000",
			5135 => "0010010010001100000100",
			5136 => "0000000101001000111101",
			5137 => "0000000101001000111101",
			5138 => "0000110011011100000100",
			5139 => "0000001101001000111101",
			5140 => "1111111101001000111101",
			5141 => "0010110100000000001000",
			5142 => "0011101011000100000100",
			5143 => "0000001101001000111101",
			5144 => "0000000101001000111101",
			5145 => "0001101100011000000100",
			5146 => "0000001101001000111101",
			5147 => "1111111101001000111101",
			5148 => "0001100100110100001100",
			5149 => "0010001011010100000100",
			5150 => "1111111101001000111101",
			5151 => "0000110101101100000100",
			5152 => "0000000101001000111101",
			5153 => "0000001101001000111101",
			5154 => "0010111000111100001000",
			5155 => "0001001111100000000100",
			5156 => "1111111101001000111101",
			5157 => "0000000101001000111101",
			5158 => "0000000101001000111101",
			5159 => "0000011110100000000100",
			5160 => "1111111101001000111101",
			5161 => "0000110101101100001100",
			5162 => "0010111100001000001000",
			5163 => "0000000100010100000100",
			5164 => "0000001101001000111101",
			5165 => "0000000101001000111101",
			5166 => "0000000101001000111101",
			5167 => "0011011100101100000100",
			5168 => "1111111101001000111101",
			5169 => "0011110100010000000100",
			5170 => "0000000101001000111101",
			5171 => "0000001101001000111101",
			5172 => "0010010111100101011000",
			5173 => "0011111011110100100000",
			5174 => "0000100111111100011100",
			5175 => "0011110110110100001100",
			5176 => "0010010110101000001000",
			5177 => "0000000001010100000100",
			5178 => "0000000101001000111101",
			5179 => "0000000101001000111101",
			5180 => "1111111101001000111101",
			5181 => "0010001001101000001000",
			5182 => "0011110010001000000100",
			5183 => "1111111101001000111101",
			5184 => "0000001101001000111101",
			5185 => "0000110101101100000100",
			5186 => "0000000101001000111101",
			5187 => "1111111101001000111101",
			5188 => "1111111101001000111101",
			5189 => "0001101100011000011100",
			5190 => "0001100001111000001100",
			5191 => "0000000011111100001000",
			5192 => "0000111101111000000100",
			5193 => "0000000101001000111101",
			5194 => "1111111101001000111101",
			5195 => "1111101101001000111101",
			5196 => "0010001011010100001000",
			5197 => "0000110000001100000100",
			5198 => "0000001101001000111101",
			5199 => "1111111101001000111101",
			5200 => "0001001101001000000100",
			5201 => "0000000101001000111101",
			5202 => "0000000101001000111101",
			5203 => "0000000100010100001100",
			5204 => "0000111100101100000100",
			5205 => "0000000101001000111101",
			5206 => "0001000000010100000100",
			5207 => "1111111101001000111101",
			5208 => "1111111101001000111101",
			5209 => "0010010110101000001000",
			5210 => "0010110000101000000100",
			5211 => "0000001101001000111101",
			5212 => "1111111101001000111101",
			5213 => "0011000000101000000100",
			5214 => "0000001101001000111101",
			5215 => "0000000101001000111101",
			5216 => "0000111110001100101100",
			5217 => "0010011101101000011100",
			5218 => "0010111100001000001100",
			5219 => "0001101101111100000100",
			5220 => "0000001101001000111101",
			5221 => "0011110101110100000100",
			5222 => "0000000101001000111101",
			5223 => "0000001101001000111101",
			5224 => "0000011100110100001000",
			5225 => "0010110100000000000100",
			5226 => "0000000101001000111101",
			5227 => "0000001101001000111101",
			5228 => "0001100100110100000100",
			5229 => "1111111101001000111101",
			5230 => "0000000101001000111101",
			5231 => "0011011101111000000100",
			5232 => "0000010101001000111101",
			5233 => "0011101000111000001000",
			5234 => "0000001111000100000100",
			5235 => "0000000101001000111101",
			5236 => "0000001101001000111101",
			5237 => "0000000101001000111101",
			5238 => "0000011100110100011000",
			5239 => "0001001010110100001100",
			5240 => "0011010000001100001000",
			5241 => "0011111010010100000100",
			5242 => "0000000101001000111101",
			5243 => "0000001101001000111101",
			5244 => "1111111101001000111101",
			5245 => "0011110010110100001000",
			5246 => "0001111100001000000100",
			5247 => "0000010101001000111101",
			5248 => "0000001101001000111101",
			5249 => "0000000101001000111101",
			5250 => "0010010111100100001100",
			5251 => "0000011100110100000100",
			5252 => "1111111101001000111101",
			5253 => "0000100010000100000100",
			5254 => "0000000101001000111101",
			5255 => "0000001101001000111101",
			5256 => "0010111100001000001000",
			5257 => "0001111100001000000100",
			5258 => "1111111101001000111101",
			5259 => "0000000101001000111101",
			5260 => "0010111000111100000100",
			5261 => "0000000101001000111101",
			5262 => "0000000101001000111101",
			5263 => "0011110000110111011000",
			5264 => "0000111001110001110100",
			5265 => "0010011001111000111100",
			5266 => "0010110000101000011100",
			5267 => "0000111000111000010000",
			5268 => "0010110100010100001000",
			5269 => "0011110110110100000100",
			5270 => "0000000101010100011011",
			5271 => "0000000101010100011011",
			5272 => "0011110000011100000100",
			5273 => "0000000101010100011011",
			5274 => "0000001101010100011011",
			5275 => "0011000000110000000100",
			5276 => "0000001101010100011011",
			5277 => "0001101101111100000100",
			5278 => "1111111101010100011011",
			5279 => "0000000101010100011011",
			5280 => "0011010110000100010000",
			5281 => "0010101100011100001000",
			5282 => "0011101010000000000100",
			5283 => "0000000101010100011011",
			5284 => "1111111101010100011011",
			5285 => "0010011001111000000100",
			5286 => "0000000101010100011011",
			5287 => "1111111101010100011011",
			5288 => "0011110111010000001000",
			5289 => "0010101100000100000100",
			5290 => "0000001101010100011011",
			5291 => "0000000101010100011011",
			5292 => "0000111100001000000100",
			5293 => "0000000101010100011011",
			5294 => "1111111101010100011011",
			5295 => "0011000111111000011000",
			5296 => "0000000000111000001100",
			5297 => "0001110000101000001000",
			5298 => "0010101001000100000100",
			5299 => "0000000101010100011011",
			5300 => "1111111101010100011011",
			5301 => "0000001101010100011011",
			5302 => "0011011100110000000100",
			5303 => "0000000101010100011011",
			5304 => "0011110000011100000100",
			5305 => "0000001101010100011011",
			5306 => "0000001101010100011011",
			5307 => "0010011001111000010000",
			5308 => "0001001001001100001000",
			5309 => "0001100111101000000100",
			5310 => "0000000101010100011011",
			5311 => "0000001101010100011011",
			5312 => "0001110100010100000100",
			5313 => "1111111101010100011011",
			5314 => "0000000101010100011011",
			5315 => "0001010110000100001000",
			5316 => "0000001110111100000100",
			5317 => "0000000101010100011011",
			5318 => "0000000101010100011011",
			5319 => "0001111100001000000100",
			5320 => "0000001101010100011011",
			5321 => "0000000101010100011011",
			5322 => "0001110100010100101000",
			5323 => "0011110111110000011000",
			5324 => "0010101001000100001100",
			5325 => "0000000010111100001000",
			5326 => "0011101000111100000100",
			5327 => "1111111101010100011011",
			5328 => "0000000101010100011011",
			5329 => "0000001101010100011011",
			5330 => "0011100100010100000100",
			5331 => "1111111101010100011011",
			5332 => "0000111101100000000100",
			5333 => "0000000101010100011011",
			5334 => "1111111101010100011011",
			5335 => "0001001000001000000100",
			5336 => "0000001101010100011011",
			5337 => "0000111101100000000100",
			5338 => "0000001101010100011011",
			5339 => "0010111011000100000100",
			5340 => "0000000101010100011011",
			5341 => "1111111101010100011011",
			5342 => "0010010110101000100000",
			5343 => "0010111011000100010000",
			5344 => "0011000100010100001000",
			5345 => "0010100110011000000100",
			5346 => "0000001101010100011011",
			5347 => "0000000101010100011011",
			5348 => "0000000000110000000100",
			5349 => "0000000101010100011011",
			5350 => "0000001101010100011011",
			5351 => "0001111011000100001000",
			5352 => "0011110101110100000100",
			5353 => "1111111101010100011011",
			5354 => "0000000101010100011011",
			5355 => "0010110100000000000100",
			5356 => "0000000101010100011011",
			5357 => "1111111101010100011011",
			5358 => "0001110000101000001100",
			5359 => "0011000000101000001000",
			5360 => "0000000010011000000100",
			5361 => "0000000101010100011011",
			5362 => "0000000101010100011011",
			5363 => "1111111101010100011011",
			5364 => "0001111100001000001000",
			5365 => "0011100011011100000100",
			5366 => "1111111101010100011011",
			5367 => "0000000101010100011011",
			5368 => "0001111000111000000100",
			5369 => "0000000101010100011011",
			5370 => "0000000101010100011011",
			5371 => "0011100100001001010100",
			5372 => "0000000000111000100100",
			5373 => "0011000100000000100000",
			5374 => "0011101101111000010000",
			5375 => "0001010000001100001000",
			5376 => "0001100100110100000100",
			5377 => "0000000101010100011011",
			5378 => "0000010101010100011011",
			5379 => "0001111100001000000100",
			5380 => "1111111101010100011011",
			5381 => "0000000101010100011011",
			5382 => "0010101001000100001000",
			5383 => "0011010001111100000100",
			5384 => "0000001101010100011011",
			5385 => "0000000101010100011011",
			5386 => "0011110110100000000100",
			5387 => "1111111101010100011011",
			5388 => "0000000101010100011011",
			5389 => "0000001101010100011011",
			5390 => "0001001101001000010000",
			5391 => "0010000111000100001100",
			5392 => "0000110001111100001000",
			5393 => "0011111110101100000100",
			5394 => "1111111101010100011011",
			5395 => "0000000101010100011011",
			5396 => "1111111101010100011011",
			5397 => "0000000101010100011011",
			5398 => "0010011101101000010000",
			5399 => "0011000100000000001000",
			5400 => "0011111101000100000100",
			5401 => "0000000101010100011011",
			5402 => "0000000101010100011011",
			5403 => "0001000100001100000100",
			5404 => "1111111101010100011011",
			5405 => "0000000101010100011011",
			5406 => "0001011010111100001000",
			5407 => "0010110011011100000100",
			5408 => "0000000101010100011011",
			5409 => "0000001101010100011011",
			5410 => "0000111010111000000100",
			5411 => "1111110101010100011011",
			5412 => "0000000101010100011011",
			5413 => "0011100001111100100000",
			5414 => "0011000100000000010100",
			5415 => "0001011010111100010000",
			5416 => "0000111110110000001000",
			5417 => "0000110111001000000100",
			5418 => "0000000101010100011011",
			5419 => "0000001101010100011011",
			5420 => "0010000111000100000100",
			5421 => "0000000101010100011011",
			5422 => "1111111101010100011011",
			5423 => "0000001101010100011011",
			5424 => "0010011111001100000100",
			5425 => "1111111101010100011011",
			5426 => "0010110000001100000100",
			5427 => "0000000101010100011011",
			5428 => "0000000101010100011011",
			5429 => "0001110000101000000100",
			5430 => "1111111101010100011011",
			5431 => "0001011100101000010000",
			5432 => "0001000011001100001000",
			5433 => "0001001000110100000100",
			5434 => "0000001101010100011011",
			5435 => "1111111101010100011011",
			5436 => "0000110100011000000100",
			5437 => "0000000101010100011011",
			5438 => "0000001101010100011011",
			5439 => "0011010111001000001000",
			5440 => "0011110101001000000100",
			5441 => "1111111101010100011011",
			5442 => "0000001101010100011011",
			5443 => "0010111101100000000100",
			5444 => "0000000101010100011011",
			5445 => "0000000101010100011011",
			5446 => "0001111110001101011000",
			5447 => "0001000110110000111100",
			5448 => "0000110010111100001000",
			5449 => "0011010100000000000100",
			5450 => "0000000101011001001101",
			5451 => "0000001101011001001101",
			5452 => "0010011100110100010100",
			5453 => "0000110000111000001000",
			5454 => "0001110111111000000100",
			5455 => "0000000101011001001101",
			5456 => "0000001101011001001101",
			5457 => "0011110110100100000100",
			5458 => "1111110101011001001101",
			5459 => "0001001001001100000100",
			5460 => "0000000101011001001101",
			5461 => "1111111101011001001101",
			5462 => "0000110100010100010000",
			5463 => "0011110001101000001000",
			5464 => "0000010110000000000100",
			5465 => "0000000101011001001101",
			5466 => "0000000101011001001101",
			5467 => "0010001000101100000100",
			5468 => "0000001101011001001101",
			5469 => "0000000101011001001101",
			5470 => "0010010010001100001000",
			5471 => "0000111100001000000100",
			5472 => "0000000101011001001101",
			5473 => "1111111101011001001101",
			5474 => "0000111001110000000100",
			5475 => "0000000101011001001101",
			5476 => "0000000101011001001101",
			5477 => "0001101100011000001000",
			5478 => "0011010110000100000100",
			5479 => "1111111101011001001101",
			5480 => "0000000101011001001101",
			5481 => "0001110100010100000100",
			5482 => "0000001101011001001101",
			5483 => "0011100000110000000100",
			5484 => "1111111101011001001101",
			5485 => "0001101011001100001000",
			5486 => "0010001101010000000100",
			5487 => "0000000101011001001101",
			5488 => "0000001101011001001101",
			5489 => "1111111101011001001101",
			5490 => "0010001001101000010000",
			5491 => "0010010100110100001100",
			5492 => "0010010001111000000100",
			5493 => "1111111101011001001101",
			5494 => "0011110110100000000100",
			5495 => "1111111101011001001101",
			5496 => "0000001101011001001101",
			5497 => "1111111101011001001101",
			5498 => "0001000011111000101000",
			5499 => "0010100001010100011000",
			5500 => "0001001011001000010000",
			5501 => "0011101100111000001000",
			5502 => "0010111010011100000100",
			5503 => "0000000101011001001101",
			5504 => "0000001101011001001101",
			5505 => "0010111110101100000100",
			5506 => "1111111101011001001101",
			5507 => "0000000101011001001101",
			5508 => "0010100101000100000100",
			5509 => "1111111101011001001101",
			5510 => "0000000101011001001101",
			5511 => "0011110000010100001000",
			5512 => "0000001011000100000100",
			5513 => "0000001101011001001101",
			5514 => "0000001101011001001101",
			5515 => "0001111001010100000100",
			5516 => "1111111101011001001101",
			5517 => "0000001101011001001101",
			5518 => "0001000000000000001000",
			5519 => "0000001010111100000100",
			5520 => "1111111101011001001101",
			5521 => "0000001101011001001101",
			5522 => "1111111101011001001101",
			5523 => "0001111101111001100000",
			5524 => "0000010000011000100000",
			5525 => "0000011100100000000100",
			5526 => "1111111101011110001001",
			5527 => "0000110000111000001100",
			5528 => "0010111110111100000100",
			5529 => "1111111101011110001001",
			5530 => "0000011100100000000100",
			5531 => "0000000101011110001001",
			5532 => "0000001101011110001001",
			5533 => "0010101100011100001100",
			5534 => "0010000010101000001000",
			5535 => "0001110100010100000100",
			5536 => "1111111101011110001001",
			5537 => "0000000101011110001001",
			5538 => "0000000101011110001001",
			5539 => "1111111101011110001001",
			5540 => "0000000100010100100100",
			5541 => "0000000110001000000100",
			5542 => "1111111101011110001001",
			5543 => "0001101101111100010000",
			5544 => "0011010100001000001000",
			5545 => "0000111100101100000100",
			5546 => "0000001101011110001001",
			5547 => "0000000101011110001001",
			5548 => "0010110101101100000100",
			5549 => "0000001101011110001001",
			5550 => "0000000101011110001001",
			5551 => "0001000110001100001000",
			5552 => "0011001001110000000100",
			5553 => "0000000101011110001001",
			5554 => "0000001101011110001001",
			5555 => "0001111100001000000100",
			5556 => "0000000101011110001001",
			5557 => "0000000101011110001001",
			5558 => "0001000100111000011000",
			5559 => "0001000011010100001100",
			5560 => "0010011011101000001000",
			5561 => "0011111001010100000100",
			5562 => "0000001101011110001001",
			5563 => "0000000101011110001001",
			5564 => "0000001101011110001001",
			5565 => "0001110111111000000100",
			5566 => "0000000101011110001001",
			5567 => "0001000000101100000100",
			5568 => "0000001101011110001001",
			5569 => "0000000101011110001001",
			5570 => "1111111101011110001001",
			5571 => "0010001001101000001100",
			5572 => "0000011011101000001000",
			5573 => "0000011011101000000100",
			5574 => "1111111101011110001001",
			5575 => "0000010101011110001001",
			5576 => "1111111101011110001001",
			5577 => "0001000010010000101000",
			5578 => "0010000110001000010100",
			5579 => "0000011110010100001000",
			5580 => "0001001110111000000100",
			5581 => "0000010101011110001001",
			5582 => "1111111101011110001001",
			5583 => "0011000001011000001000",
			5584 => "0010001001101000000100",
			5585 => "0000000101011110001001",
			5586 => "1111111101011110001001",
			5587 => "0000001101011110001001",
			5588 => "0011111111100000010000",
			5589 => "0011001000000000001000",
			5590 => "0010011010011000000100",
			5591 => "0000001101011110001001",
			5592 => "0000000101011110001001",
			5593 => "0001000011110100000100",
			5594 => "0000010101011110001001",
			5595 => "0000000101011110001001",
			5596 => "1111111101011110001001",
			5597 => "0001000000000000001000",
			5598 => "0001001010101000000100",
			5599 => "1111111101011110001001",
			5600 => "0000000101011110001001",
			5601 => "1111111101011110001001",
			5602 => "0001111101111001100000",
			5603 => "0001000110110001000100",
			5604 => "0001100001000100001000",
			5605 => "0001100001000100000100",
			5606 => "1111111101100010111101",
			5607 => "0000000101100010111101",
			5608 => "0011100110000100100000",
			5609 => "0010011101101000010000",
			5610 => "0001001110111000001000",
			5611 => "0001101101111100000100",
			5612 => "0000001101100010111101",
			5613 => "0000000101100010111101",
			5614 => "0010010110101000000100",
			5615 => "0000001101100010111101",
			5616 => "0000001101100010111101",
			5617 => "0001010000001100001000",
			5618 => "0001000010111000000100",
			5619 => "0000011101100010111101",
			5620 => "0000001101100010111101",
			5621 => "0001000011110000000100",
			5622 => "0000001101100010111101",
			5623 => "0000001101100010111101",
			5624 => "0011001000111100010000",
			5625 => "0001101011001100001000",
			5626 => "0001110100000000000100",
			5627 => "0000000101100010111101",
			5628 => "0000000101100010111101",
			5629 => "0001111101100000000100",
			5630 => "1111111101100010111101",
			5631 => "0000000101100010111101",
			5632 => "0010010100110100001000",
			5633 => "0001101010011000000100",
			5634 => "0000000101100010111101",
			5635 => "0000001101100010111101",
			5636 => "1111111101100010111101",
			5637 => "0001101100011000001000",
			5638 => "0010111100001000000100",
			5639 => "1111111101100010111101",
			5640 => "1111111101100010111101",
			5641 => "0001110100010100000100",
			5642 => "0000001101100010111101",
			5643 => "0001000001001100000100",
			5644 => "0000000101100010111101",
			5645 => "0010010010001100001000",
			5646 => "0010010000011000000100",
			5647 => "1111111101100010111101",
			5648 => "0000000101100010111101",
			5649 => "1111111101100010111101",
			5650 => "0010001001101000001100",
			5651 => "0011000110000100001000",
			5652 => "0001110100001000000100",
			5653 => "1111111101100010111101",
			5654 => "0000001101100010111101",
			5655 => "1111111101100010111101",
			5656 => "0001000010010000101100",
			5657 => "0010001111001000011000",
			5658 => "0011111000000100001100",
			5659 => "0001000100001100001000",
			5660 => "0010010111101100000100",
			5661 => "0000010101100010111101",
			5662 => "0000000101100010111101",
			5663 => "1111111101100010111101",
			5664 => "0010001001101000000100",
			5665 => "0000000101100010111101",
			5666 => "0001110111110000000100",
			5667 => "1111111101100010111101",
			5668 => "0000000101100010111101",
			5669 => "0011000110000100000100",
			5670 => "1111111101100010111101",
			5671 => "0011110000010100001000",
			5672 => "0011011100000000000100",
			5673 => "0000001101100010111101",
			5674 => "0000010101100010111101",
			5675 => "0001100100101100000100",
			5676 => "1111111101100010111101",
			5677 => "0000001101100010111101",
			5678 => "1111111101100010111101",
			5679 => "0001000011011001110100",
			5680 => "0000001100001001001100",
			5681 => "0001001011101100011100",
			5682 => "0010000110011100011000",
			5683 => "0001000000010000001100",
			5684 => "0000111010111000001000",
			5685 => "0000011100110100000100",
			5686 => "1111111101101001100001",
			5687 => "0000001101101001100001",
			5688 => "1111111101101001100001",
			5689 => "0000010110101000001000",
			5690 => "0001111100001000000100",
			5691 => "0000000101101001100001",
			5692 => "0000001101101001100001",
			5693 => "1111111101101001100001",
			5694 => "1111111101101001100001",
			5695 => "0010000101000100010000",
			5696 => "0010110001111100001100",
			5697 => "0011010001111100001000",
			5698 => "0000110000001100000100",
			5699 => "0000001101101001100001",
			5700 => "1111111101101001100001",
			5701 => "0000001101101001100001",
			5702 => "1111111101101001100001",
			5703 => "0000101110101000010000",
			5704 => "0001000100001100001000",
			5705 => "0000011100110100000100",
			5706 => "0000000101101001100001",
			5707 => "1111111101101001100001",
			5708 => "0000110000111000000100",
			5709 => "0000001101101001100001",
			5710 => "1111111101101001100001",
			5711 => "0000010110000000001000",
			5712 => "0000111011000100000100",
			5713 => "0000000101101001100001",
			5714 => "1111111101101001100001",
			5715 => "0000111100001000000100",
			5716 => "0000000101101001100001",
			5717 => "0000000101101001100001",
			5718 => "0011100000101000011100",
			5719 => "0010110111111000001100",
			5720 => "0001011000111100001000",
			5721 => "0001011000111100000100",
			5722 => "0000001101101001100001",
			5723 => "0000000101101001100001",
			5724 => "1111111101101001100001",
			5725 => "0010001000110000001100",
			5726 => "0001110000101000000100",
			5727 => "0000001101101001100001",
			5728 => "0011100000111000000100",
			5729 => "0000000101101001100001",
			5730 => "0000001101101001100001",
			5731 => "0000000101101001100001",
			5732 => "0011100100000000000100",
			5733 => "1111110101101001100001",
			5734 => "0000010010001100000100",
			5735 => "0000001101101001100001",
			5736 => "0000000101101001100001",
			5737 => "0011111001010100110000",
			5738 => "0000011110100000100100",
			5739 => "0001110111111000010000",
			5740 => "0011100111000100001000",
			5741 => "0001110111111000000100",
			5742 => "1111111101101001100001",
			5743 => "0000000101101001100001",
			5744 => "0010111110111100000100",
			5745 => "1111111101101001100001",
			5746 => "1111110101101001100001",
			5747 => "0001001101110100000100",
			5748 => "0000001101101001100001",
			5749 => "0000101001010000001000",
			5750 => "0011101011010100000100",
			5751 => "1111111101101001100001",
			5752 => "0000000101101001100001",
			5753 => "0000100010011100000100",
			5754 => "1111110101101001100001",
			5755 => "0000000101101001100001",
			5756 => "0011000000101000000100",
			5757 => "1111101101101001100001",
			5758 => "0000111100101100000100",
			5759 => "0000001101101001100001",
			5760 => "0000000101101001100001",
			5761 => "0001111101111000011000",
			5762 => "0000101100010000001000",
			5763 => "0000111101111000000100",
			5764 => "0000001101101001100001",
			5765 => "1111111101101001100001",
			5766 => "0000001100001000000100",
			5767 => "0000000101101001100001",
			5768 => "0001000001001100001000",
			5769 => "0001111001110000000100",
			5770 => "0000001101101001100001",
			5771 => "0000001101101001100001",
			5772 => "0000000101101001100001",
			5773 => "0010001010101100000100",
			5774 => "1111111101101001100001",
			5775 => "0011001001110100001100",
			5776 => "0001010110110100001000",
			5777 => "0011100001111100000100",
			5778 => "0000000101101001100001",
			5779 => "1111111101101001100001",
			5780 => "0000001101101001100001",
			5781 => "0011101011111000000100",
			5782 => "0000000101101001100001",
			5783 => "1111111101101001100001",
			5784 => "0001111101111001100000",
			5785 => "0001000110110001001000",
			5786 => "0001100001000100001000",
			5787 => "0001100001000100000100",
			5788 => "1111111101101110011101",
			5789 => "0000000101101110011101",
			5790 => "0011101000111100100000",
			5791 => "0001111011000100010000",
			5792 => "0000111100001000001000",
			5793 => "0011000000110000000100",
			5794 => "0000000101101110011101",
			5795 => "0000001101101110011101",
			5796 => "0010010010001100000100",
			5797 => "1111111101101110011101",
			5798 => "0000000101101110011101",
			5799 => "0000101001011100001000",
			5800 => "0001100001111000000100",
			5801 => "0000001101101110011101",
			5802 => "0000001101101110011101",
			5803 => "0000000000111000000100",
			5804 => "0000010101101110011101",
			5805 => "0000001101101110011101",
			5806 => "0001000010111000010000",
			5807 => "0011001000111100001000",
			5808 => "0010100110011000000100",
			5809 => "0000000101101110011101",
			5810 => "0000000101101110011101",
			5811 => "0010011101111100000100",
			5812 => "0000001101101110011101",
			5813 => "1111111101101110011101",
			5814 => "0001101001100100001000",
			5815 => "0010011101101000000100",
			5816 => "0000000101101110011101",
			5817 => "0000001101101110011101",
			5818 => "0011001000111000000100",
			5819 => "1111111101101110011101",
			5820 => "0000001101101110011101",
			5821 => "0001101100011000000100",
			5822 => "1111111101101110011101",
			5823 => "0001110100010100000100",
			5824 => "0000001101101110011101",
			5825 => "0001000001001100000100",
			5826 => "0000000101101110011101",
			5827 => "0010010010001100001000",
			5828 => "0010010000011000000100",
			5829 => "1111111101101110011101",
			5830 => "0000000101101110011101",
			5831 => "1111111101101110011101",
			5832 => "0010001001101000001100",
			5833 => "0011000110000100001000",
			5834 => "0001110100001000000100",
			5835 => "1111111101101110011101",
			5836 => "0000001101101110011101",
			5837 => "1111111101101110011101",
			5838 => "0001000010010000110000",
			5839 => "0010001111001000011000",
			5840 => "0011111000000100001100",
			5841 => "0001000100001100001000",
			5842 => "0001000011001100000100",
			5843 => "0000000101101110011101",
			5844 => "0000010101101110011101",
			5845 => "1111111101101110011101",
			5846 => "0010001001101000000100",
			5847 => "0000000101101110011101",
			5848 => "0001110111110000000100",
			5849 => "1111111101101110011101",
			5850 => "0000000101101110011101",
			5851 => "0010001010101100010000",
			5852 => "0001000011011000001000",
			5853 => "0001001001001100000100",
			5854 => "0000000101101110011101",
			5855 => "0000001101101110011101",
			5856 => "0000000000110000000100",
			5857 => "0000000101101110011101",
			5858 => "1111111101101110011101",
			5859 => "0000010000111100000100",
			5860 => "0000001101101110011101",
			5861 => "0000010101101110011101",
			5862 => "1111111101101110011101",
			5863 => "0010110000001101101100",
			5864 => "0000010000011000011000",
			5865 => "0001101101111100001100",
			5866 => "0001001011100000001000",
			5867 => "0001000011010100000100",
			5868 => "1111111101110100011001",
			5869 => "0000000101110100011001",
			5870 => "1111111101110100011001",
			5871 => "0011010011011100001000",
			5872 => "0000111000110000000100",
			5873 => "0000001101110100011001",
			5874 => "0000000101110100011001",
			5875 => "1111111101110100011001",
			5876 => "0011101100001000100100",
			5877 => "0001100001000100000100",
			5878 => "1111111101110100011001",
			5879 => "0011011100101100010000",
			5880 => "0000111001110000001000",
			5881 => "0010110111111000000100",
			5882 => "0000001101110100011001",
			5883 => "0000001101110100011001",
			5884 => "0000001011000100000100",
			5885 => "0000000101110100011001",
			5886 => "0000001101110100011001",
			5887 => "0001100001111000001000",
			5888 => "0011100111111000000100",
			5889 => "0000001101110100011001",
			5890 => "0000010101110100011001",
			5891 => "0011110100000100000100",
			5892 => "0000000101110100011001",
			5893 => "0000001101110100011001",
			5894 => "0001001010110100010100",
			5895 => "0001101011111100000100",
			5896 => "1111111101110100011001",
			5897 => "0001101101111100001000",
			5898 => "0011110110110100000100",
			5899 => "0000000101110100011001",
			5900 => "0000001101110100011001",
			5901 => "0000001010000000000100",
			5902 => "0000000101110100011001",
			5903 => "0000010101110100011001",
			5904 => "0001101001100100010000",
			5905 => "0010111100001000001000",
			5906 => "0001011101100000000100",
			5907 => "1111111101110100011001",
			5908 => "0000000101110100011001",
			5909 => "0001000100001100000100",
			5910 => "0000001101110100011001",
			5911 => "0000001101110100011001",
			5912 => "0011110010000100001000",
			5913 => "0011111100100100000100",
			5914 => "0000000101110100011001",
			5915 => "1111111101110100011001",
			5916 => "0000001101110100011001",
			5917 => "0011001110001100101100",
			5918 => "0011110101110000010000",
			5919 => "0001011000000000000100",
			5920 => "0000000101110100011001",
			5921 => "0011111110000100000100",
			5922 => "1111111101110100011001",
			5923 => "0010110100001000000100",
			5924 => "0000001101110100011001",
			5925 => "1111111101110100011001",
			5926 => "0010010100110100010100",
			5927 => "0001000001001100010000",
			5928 => "0011110010000100001000",
			5929 => "0011010111010000000100",
			5930 => "0000001101110100011001",
			5931 => "0000000101110100011001",
			5932 => "0000000000111000000100",
			5933 => "0000010101110100011001",
			5934 => "0000001101110100011001",
			5935 => "1111111101110100011001",
			5936 => "0000000111111000000100",
			5937 => "1111111101110100011001",
			5938 => "0000000101110100011001",
			5939 => "0010001001101000000100",
			5940 => "1111111101110100011001",
			5941 => "0001000110110000100000",
			5942 => "0011101101101100010000",
			5943 => "0001000011101100001000",
			5944 => "0010010100101100000100",
			5945 => "0000010101110100011001",
			5946 => "0000000101110100011001",
			5947 => "0010100110011100000100",
			5948 => "1111111101110100011001",
			5949 => "0000010101110100011001",
			5950 => "0001100100101100001000",
			5951 => "0011001011011100000100",
			5952 => "1111111101110100011001",
			5953 => "0000001101110100011001",
			5954 => "0010000001110100000100",
			5955 => "0000000101110100011001",
			5956 => "0000001101110100011001",
			5957 => "1111111101110100011001",
			5958 => "0001111110001110000000",
			5959 => "0001000110110001100000",
			5960 => "0000110100010100100000",
			5961 => "0011000000110000010000",
			5962 => "0000100110100000000100",
			5963 => "0000000101111010101101",
			5964 => "0011110100000100001000",
			5965 => "0001011000111100000100",
			5966 => "0000001101111010101101",
			5967 => "1111111101111010101101",
			5968 => "0000001101111010101101",
			5969 => "0010100111110100000100",
			5970 => "1111111101111010101101",
			5971 => "0011110111010000001000",
			5972 => "0000101001010000000100",
			5973 => "0000000101111010101101",
			5974 => "1111111101111010101101",
			5975 => "0000001101111010101101",
			5976 => "0010010010001100100000",
			5977 => "0000111100001000010000",
			5978 => "0010111110111100001000",
			5979 => "0000111011000100000100",
			5980 => "0000001101111010101101",
			5981 => "1111111101111010101101",
			5982 => "0000101111010000000100",
			5983 => "0000000101111010101101",
			5984 => "0000000101111010101101",
			5985 => "0011110101100100001000",
			5986 => "0001010011011100000100",
			5987 => "1111110101111010101101",
			5988 => "1111111101111010101101",
			5989 => "0010010010001100000100",
			5990 => "1111111101111010101101",
			5991 => "0000000101111010101101",
			5992 => "0000111001110000010000",
			5993 => "0011110101100100001000",
			5994 => "0010101001000100000100",
			5995 => "0000000101111010101101",
			5996 => "0000000101111010101101",
			5997 => "0010011001111000000100",
			5998 => "0000000101111010101101",
			5999 => "0000001101111010101101",
			6000 => "0011011100101100001000",
			6001 => "0010010110101000000100",
			6002 => "0000000101111010101101",
			6003 => "0000000101111010101101",
			6004 => "0011001010000000000100",
			6005 => "0000001101111010101101",
			6006 => "0000000101111010101101",
			6007 => "0001101100011000001000",
			6008 => "0011010110000100000100",
			6009 => "1111111101111010101101",
			6010 => "0000000101111010101101",
			6011 => "0001110100010100000100",
			6012 => "0000001101111010101101",
			6013 => "0010100001110000001000",
			6014 => "0011000011011100000100",
			6015 => "0000000101111010101101",
			6016 => "0000000101111010101101",
			6017 => "0011000000101000000100",
			6018 => "1111111101111010101101",
			6019 => "0000111110001100000100",
			6020 => "0000000101111010101101",
			6021 => "1111111101111010101101",
			6022 => "0010001001101000010000",
			6023 => "0000011011101000001100",
			6024 => "0010010001111000000100",
			6025 => "1111111101111010101101",
			6026 => "0000100111100000000100",
			6027 => "1111111101111010101101",
			6028 => "0000001101111010101101",
			6029 => "1111111101111010101101",
			6030 => "0001000011111000101100",
			6031 => "0011000110000100010000",
			6032 => "0001000000101100001000",
			6033 => "0010100110011000000100",
			6034 => "0000000101111010101101",
			6035 => "1111111101111010101101",
			6036 => "0000011101011100000100",
			6037 => "1111111101111010101101",
			6038 => "0000000101111010101101",
			6039 => "0000011011101000001100",
			6040 => "0001011001010100001000",
			6041 => "0010111110110000000100",
			6042 => "0000001101111010101101",
			6043 => "0000010101111010101101",
			6044 => "1111111101111010101101",
			6045 => "0011000001011000001000",
			6046 => "0010010111101100000100",
			6047 => "0000000101111010101101",
			6048 => "0000000101111010101101",
			6049 => "0000010100110100000100",
			6050 => "0000000101111010101101",
			6051 => "0000001101111010101101",
			6052 => "0001000000000000001100",
			6053 => "0011000000001100001000",
			6054 => "0010001101010000000100",
			6055 => "0000000101111010101101",
			6056 => "0000001101111010101101",
			6057 => "1111111101111010101101",
			6058 => "1111111101111010101101",
			6059 => "0000110000110001001000",
			6060 => "0011100001110100111100",
			6061 => "0000110011111100100100",
			6062 => "0000100000110100001000",
			6063 => "0011110101101100000100",
			6064 => "0000000110000001100001",
			6065 => "0000001110000001100001",
			6066 => "0011111010111000001100",
			6067 => "0001101100011000001000",
			6068 => "0011111010111000000100",
			6069 => "1111111110000001100001",
			6070 => "0000000110000001100001",
			6071 => "0000000110000001100001",
			6072 => "0011000111111000001000",
			6073 => "0000000100000000000100",
			6074 => "0000000110000001100001",
			6075 => "0000000110000001100001",
			6076 => "0001001110011000000100",
			6077 => "0000001110000001100001",
			6078 => "0000000110000001100001",
			6079 => "0011011000111100001000",
			6080 => "0010111010000000000100",
			6081 => "1111111110000001100001",
			6082 => "1111101110000001100001",
			6083 => "0010110100010100001000",
			6084 => "0001111010000000000100",
			6085 => "0000000110000001100001",
			6086 => "1111111110000001100001",
			6087 => "0001001010101000000100",
			6088 => "0000001110000001100001",
			6089 => "0000000110000001100001",
			6090 => "0001101110010100000100",
			6091 => "1111111110000001100001",
			6092 => "0000101001010000000100",
			6093 => "0000001110000001100001",
			6094 => "0000000110000001100001",
			6095 => "0011110110100100111000",
			6096 => "0001100001111000011000",
			6097 => "0011011100110000001000",
			6098 => "0000110111111000000100",
			6099 => "0000000110000001100001",
			6100 => "1111111110000001100001",
			6101 => "0001111011000100001000",
			6102 => "0010011001111000000100",
			6103 => "0000001110000001100001",
			6104 => "1111111110000001100001",
			6105 => "0000000110001000000100",
			6106 => "0000000110000001100001",
			6107 => "0000001110000001100001",
			6108 => "0010110111111000000100",
			6109 => "0000000110000001100001",
			6110 => "0000001011000100001100",
			6111 => "0001000000010100001000",
			6112 => "0000101110101100000100",
			6113 => "1111111110000001100001",
			6114 => "0000000110000001100001",
			6115 => "1111110110000001100001",
			6116 => "0011110110100100001000",
			6117 => "0000000110000100000100",
			6118 => "0000001110000001100001",
			6119 => "0000000110000001100001",
			6120 => "0001100100110100000100",
			6121 => "0000000110000001100001",
			6122 => "1111111110000001100001",
			6123 => "0000111011000100100000",
			6124 => "0010001001101000001000",
			6125 => "0000110100010100000100",
			6126 => "1111110110000001100001",
			6127 => "0000000110000001100001",
			6128 => "0001000000010100001000",
			6129 => "0011000100010100000100",
			6130 => "0000001110000001100001",
			6131 => "0000000110000001100001",
			6132 => "0000000100010100001000",
			6133 => "0011111010001100000100",
			6134 => "1111111110000001100001",
			6135 => "0000000110000001100001",
			6136 => "0001110111111000000100",
			6137 => "0000000110000001100001",
			6138 => "0000000110000001100001",
			6139 => "0010011001111000011100",
			6140 => "0000101110000100001100",
			6141 => "0011100010011000000100",
			6142 => "0000000110000001100001",
			6143 => "0001001101001000000100",
			6144 => "0000000110000001100001",
			6145 => "1111111110000001100001",
			6146 => "0000111100001000001000",
			6147 => "0000100010011100000100",
			6148 => "0000001110000001100001",
			6149 => "0000000110000001100001",
			6150 => "0011110101100100000100",
			6151 => "1111111110000001100001",
			6152 => "0000000110000001100001",
			6153 => "0011101101111000010000",
			6154 => "0011110010110100001000",
			6155 => "0011000000110000000100",
			6156 => "1111111110000001100001",
			6157 => "0000000110000001100001",
			6158 => "0010100110011000000100",
			6159 => "0000001110000001100001",
			6160 => "0000000110000001100001",
			6161 => "0001111000111000001000",
			6162 => "0001110100000000000100",
			6163 => "0000000110000001100001",
			6164 => "0000000110000001100001",
			6165 => "0011110111110000000100",
			6166 => "0000001110000001100001",
			6167 => "0000000110000001100001",
			6168 => "0001011000000010001000",
			6169 => "0000010000011000010100",
			6170 => "0001101101111100001000",
			6171 => "0000100101110100000100",
			6172 => "0000000110001000101101",
			6173 => "1111111110001000101101",
			6174 => "0000011100100000000100",
			6175 => "1111111110001000101101",
			6176 => "0001110111111000000100",
			6177 => "0000000110001000101101",
			6178 => "0000010110001000101101",
			6179 => "0011101101100000110100",
			6180 => "0000001010000000011100",
			6181 => "0011100111111000001100",
			6182 => "0001100001000100000100",
			6183 => "1111111110001000101101",
			6184 => "0010100001010000000100",
			6185 => "0000010110001000101101",
			6186 => "0000000110001000101101",
			6187 => "0001111011000100001000",
			6188 => "0001100100110100000100",
			6189 => "0000001110001000101101",
			6190 => "0000000110001000101101",
			6191 => "0000100101110000000100",
			6192 => "0000001110001000101101",
			6193 => "0000001110001000101101",
			6194 => "0011000000110000001000",
			6195 => "0000100001000000000100",
			6196 => "0000001110001000101101",
			6197 => "1111111110001000101101",
			6198 => "0001010110000100001000",
			6199 => "0011100100010100000100",
			6200 => "0000010110001000101101",
			6201 => "0000001110001000101101",
			6202 => "0010110101101100000100",
			6203 => "0000010110001000101101",
			6204 => "1111111110001000101101",
			6205 => "0000000000110000100000",
			6206 => "0000101010001000010000",
			6207 => "0001110100000000001000",
			6208 => "0011101100101000000100",
			6209 => "0000000110001000101101",
			6210 => "1111111110001000101101",
			6211 => "0000100010110100000100",
			6212 => "1111111110001000101101",
			6213 => "0000000110001000101101",
			6214 => "0001100100110100001000",
			6215 => "0001011101111000000100",
			6216 => "0000000110001000101101",
			6217 => "0000011110001000101101",
			6218 => "0011000100000000000100",
			6219 => "0000000110001000101101",
			6220 => "0000001110001000101101",
			6221 => "0001101001100100010000",
			6222 => "0011000100000000001000",
			6223 => "0000000111111000000100",
			6224 => "0000001110001000101101",
			6225 => "0000001110001000101101",
			6226 => "0000011001111000000100",
			6227 => "0000010110001000101101",
			6228 => "0000010110001000101101",
			6229 => "0001111101100000001000",
			6230 => "0000101000001100000100",
			6231 => "1111111110001000101101",
			6232 => "0000000110001000101101",
			6233 => "0001101111000000000100",
			6234 => "0000010110001000101101",
			6235 => "0000000110001000101101",
			6236 => "0001111101111000111000",
			6237 => "0011100001101000010100",
			6238 => "0001011000000000001000",
			6239 => "0000111110110000000100",
			6240 => "1111111110001000101101",
			6241 => "0000001110001000101101",
			6242 => "0000100010000000000100",
			6243 => "1111111110001000101101",
			6244 => "0000001000111100000100",
			6245 => "0000001110001000101101",
			6246 => "1111111110001000101101",
			6247 => "0010010001111000011000",
			6248 => "0001111101100000001100",
			6249 => "0001101011001100000100",
			6250 => "0000001110001000101101",
			6251 => "0000010111100100000100",
			6252 => "0000001110001000101101",
			6253 => "1111111110001000101101",
			6254 => "0000001010101100000100",
			6255 => "1111111110001000101101",
			6256 => "0010000010101000000100",
			6257 => "0000010110001000101101",
			6258 => "0000000110001000101101",
			6259 => "0000000111111000001000",
			6260 => "0011001110001100000100",
			6261 => "1111111110001000101101",
			6262 => "0000001110001000101101",
			6263 => "0000001110001000101101",
			6264 => "0010011000010100100000",
			6265 => "0010001001101000001100",
			6266 => "0011000110000100001000",
			6267 => "0011000110000100000100",
			6268 => "1111111110001000101101",
			6269 => "0000000110001000101101",
			6270 => "1111111110001000101101",
			6271 => "0000001000111100010000",
			6272 => "0010001111001000001000",
			6273 => "0010011010011000000100",
			6274 => "0000010110001000101101",
			6275 => "1111111110001000101101",
			6276 => "0000101110111000000100",
			6277 => "0000001110001000101101",
			6278 => "0000000110001000101101",
			6279 => "1111111110001000101101",
			6280 => "0001110101110100000100",
			6281 => "1111111110001000101101",
			6282 => "0000001110001000101101",
			6283 => "0001011000000010001100",
			6284 => "0000010000011000011100",
			6285 => "0000011100100000000100",
			6286 => "1111111110001111111001",
			6287 => "0011111000000000001100",
			6288 => "0001110111111000000100",
			6289 => "0000000110001111111001",
			6290 => "0000101101000100000100",
			6291 => "0000010110001111111001",
			6292 => "0000001110001111111001",
			6293 => "0000101001010000001000",
			6294 => "0000000111111000000100",
			6295 => "1111111110001111111001",
			6296 => "0000000110001111111001",
			6297 => "1111111110001111111001",
			6298 => "0001001001001100111100",
			6299 => "0000110101101100011100",
			6300 => "0000110100000000001100",
			6301 => "0010000101000100000100",
			6302 => "0000000110001111111001",
			6303 => "0010100001010000000100",
			6304 => "0000001110001111111001",
			6305 => "0000000110001111111001",
			6306 => "0010111100001000001000",
			6307 => "0011110111110000000100",
			6308 => "0000001110001111111001",
			6309 => "0000010110001111111001",
			6310 => "0010000001010100000100",
			6311 => "0000010110001111111001",
			6312 => "0000001110001111111001",
			6313 => "0001110100000000010000",
			6314 => "0000111101111000001000",
			6315 => "0011011100101000000100",
			6316 => "0000000110001111111001",
			6317 => "0000010110001111111001",
			6318 => "0010100001010000000100",
			6319 => "0000000110001111111001",
			6320 => "1111111110001111111001",
			6321 => "0000010110101000001000",
			6322 => "0001000000010000000100",
			6323 => "1111111110001111111001",
			6324 => "0000001110001111111001",
			6325 => "0000100111011000000100",
			6326 => "1111111110001111111001",
			6327 => "0000000110001111111001",
			6328 => "0000110001101000100000",
			6329 => "0001111100001000010000",
			6330 => "0000000100010100001000",
			6331 => "0000111000111100000100",
			6332 => "0000001110001111111001",
			6333 => "0000001110001111111001",
			6334 => "0001000000100000000100",
			6335 => "0000001110001111111001",
			6336 => "0000001110001111111001",
			6337 => "0001000110110000001000",
			6338 => "0001000100001100000100",
			6339 => "0000001110001111111001",
			6340 => "0000010110001111111001",
			6341 => "0000110111001000000100",
			6342 => "0000000110001111111001",
			6343 => "1111111110001111111001",
			6344 => "0011001001110000010000",
			6345 => "0010101100011100001000",
			6346 => "0001000100001100000100",
			6347 => "0000000110001111111001",
			6348 => "0000010110001111111001",
			6349 => "0011110011001000000100",
			6350 => "1111111110001111111001",
			6351 => "0000001110001111111001",
			6352 => "0000001110001111111001",
			6353 => "0001111101111000110000",
			6354 => "0011111101000100001000",
			6355 => "0011011000000000000100",
			6356 => "0000000110001111111001",
			6357 => "1111111110001111111001",
			6358 => "0000011011101000011100",
			6359 => "0010100101000100010000",
			6360 => "0011001000111000001000",
			6361 => "0010011011111100000100",
			6362 => "0000000110001111111001",
			6363 => "1111111110001111111001",
			6364 => "0001111101100000000100",
			6365 => "0000000110001111111001",
			6366 => "0000001110001111111001",
			6367 => "0011010001011000001000",
			6368 => "0011000110000100000100",
			6369 => "1111111110001111111001",
			6370 => "0000000110001111111001",
			6371 => "0000000110001111111001",
			6372 => "0011001100110000000100",
			6373 => "1111111110001111111001",
			6374 => "0011110010000000000100",
			6375 => "1111111110001111111001",
			6376 => "0000001110001111111001",
			6377 => "0010001001101000001100",
			6378 => "0001111100101000001000",
			6379 => "0011000110000100000100",
			6380 => "0000000110001111111001",
			6381 => "1111111110001111111001",
			6382 => "1111111110001111111001",
			6383 => "0001000010010000011000",
			6384 => "0010001111001000001100",
			6385 => "0010011010011000000100",
			6386 => "0000010110001111111001",
			6387 => "0011001011011100000100",
			6388 => "1111111110001111111001",
			6389 => "0000000110001111111001",
			6390 => "0010000111000000001000",
			6391 => "0001000001101100000100",
			6392 => "0000001110001111111001",
			6393 => "1111111110001111111001",
			6394 => "0000010110001111111001",
			6395 => "0000011001011000000100",
			6396 => "1111111110001111111001",
			6397 => "0000000110001111111001",
			6398 => "0001010011100010001000",
			6399 => "0000010000011000011100",
			6400 => "0001101101111100010000",
			6401 => "0010011110100000001000",
			6402 => "0000100101110100000100",
			6403 => "0000000110010111100101",
			6404 => "1111111110010111100101",
			6405 => "0000101010001000000100",
			6406 => "0000000110010111100101",
			6407 => "1111111110010111100101",
			6408 => "0011010011011100001000",
			6409 => "0001110111111000000100",
			6410 => "0000000110010111100101",
			6411 => "0000011110010111100101",
			6412 => "1111111110010111100101",
			6413 => "0011101000111000110100",
			6414 => "0011100111111000010100",
			6415 => "0001100001000100000100",
			6416 => "1111111110010111100101",
			6417 => "0001111011000100001000",
			6418 => "0000110000101000000100",
			6419 => "0000010110010111100101",
			6420 => "0000010110010111100101",
			6421 => "0001100001111000000100",
			6422 => "0000011110010111100101",
			6423 => "0000010110010111100101",
			6424 => "0000100100101000010000",
			6425 => "0011010000001100001000",
			6426 => "0010101001000100000100",
			6427 => "0000001110010111100101",
			6428 => "0000001110010111100101",
			6429 => "0011111010001100000100",
			6430 => "0000001110010111100101",
			6431 => "0000010110010111100101",
			6432 => "0001111011000100001000",
			6433 => "0010101100011100000100",
			6434 => "0000001110010111100101",
			6435 => "0000010110010111100101",
			6436 => "0011011010111100000100",
			6437 => "0000010110010111100101",
			6438 => "1111111110010111100101",
			6439 => "0000100111111100011100",
			6440 => "0010101010110000010000",
			6441 => "0001101101111100001000",
			6442 => "0001101110010100000100",
			6443 => "1111111110010111100101",
			6444 => "0000001110010111100101",
			6445 => "0001101010011000000100",
			6446 => "0000000110010111100101",
			6447 => "0000001110010111100101",
			6448 => "0010011101101000000100",
			6449 => "0000000110010111100101",
			6450 => "0000100100101000000100",
			6451 => "0000011110010111100101",
			6452 => "0000010110010111100101",
			6453 => "0001101001100100010000",
			6454 => "0011000100000000001000",
			6455 => "0011100110000100000100",
			6456 => "0000010110010111100101",
			6457 => "0000001110010111100101",
			6458 => "0010100110011000000100",
			6459 => "0000001110010111100101",
			6460 => "0000010110010111100101",
			6461 => "0001111101100000001000",
			6462 => "0000111001001000000100",
			6463 => "0000000110010111100101",
			6464 => "1111111110010111100101",
			6465 => "0000010110010111100101",
			6466 => "0001111101111001000100",
			6467 => "0011111110101100001100",
			6468 => "0011110100010000000100",
			6469 => "1111111110010111100101",
			6470 => "0011110001001000000100",
			6471 => "0000000110010111100101",
			6472 => "1111111110010111100101",
			6473 => "0001101011001100011000",
			6474 => "0011011111011100001100",
			6475 => "0010001000101100001000",
			6476 => "0001110101101100000100",
			6477 => "0000001110010111100101",
			6478 => "0000011110010111100101",
			6479 => "1111111110010111100101",
			6480 => "0011111100010100001000",
			6481 => "0001101011001100000100",
			6482 => "1111111110010111100101",
			6483 => "0000000110010111100101",
			6484 => "0000001110010111100101",
			6485 => "0001110101101100010000",
			6486 => "0000010110101000001000",
			6487 => "0011100110100100000100",
			6488 => "1111111110010111100101",
			6489 => "0000010110010111100101",
			6490 => "0000010111100100000100",
			6491 => "0000000110010111100101",
			6492 => "1111111110010111100101",
			6493 => "0000100000010000001000",
			6494 => "0000011101101000000100",
			6495 => "0000011110010111100101",
			6496 => "0000001110010111100101",
			6497 => "0011111001100000000100",
			6498 => "1111111110010111100101",
			6499 => "0000000110010111100101",
			6500 => "0010011000010100100100",
			6501 => "0010001001101000001100",
			6502 => "0011000110000100001000",
			6503 => "0000100111010100000100",
			6504 => "1111111110010111100101",
			6505 => "0000000110010111100101",
			6506 => "1111111110010111100101",
			6507 => "0010001101010000010000",
			6508 => "0010001111001000001000",
			6509 => "0010011010011000000100",
			6510 => "0000010110010111100101",
			6511 => "1111111110010111100101",
			6512 => "0000011001011000000100",
			6513 => "0000000110010111100101",
			6514 => "0000001110010111100101",
			6515 => "0010101100000100000100",
			6516 => "0000000110010111100101",
			6517 => "1111111110010111100101",
			6518 => "0001110101110100000100",
			6519 => "1111111110010111100101",
			6520 => "0000001110010111100101",
			6521 => "0001001011101100100000",
			6522 => "0010000110011100011100",
			6523 => "0001000000010000010100",
			6524 => "0011110100000100001100",
			6525 => "0011111001110100000100",
			6526 => "1111111110011101010001",
			6527 => "0001100001000100000100",
			6528 => "0000000110011101010001",
			6529 => "0000001110011101010001",
			6530 => "0001101110010100000100",
			6531 => "0000000110011101010001",
			6532 => "1111111110011101010001",
			6533 => "0001100001111000000100",
			6534 => "0000001110011101010001",
			6535 => "1111111110011101010001",
			6536 => "1111111110011101010001",
			6537 => "0010000101000100011000",
			6538 => "0010110001111100010100",
			6539 => "0011010001111100010000",
			6540 => "0000110000001100001100",
			6541 => "0011010110000100001000",
			6542 => "0011111010001100000100",
			6543 => "0000000110011101010001",
			6544 => "1111111110011101010001",
			6545 => "0000001110011101010001",
			6546 => "1111111110011101010001",
			6547 => "0000001110011101010001",
			6548 => "1111111110011101010001",
			6549 => "0000100111111101000000",
			6550 => "0000100111111100100000",
			6551 => "0000100100101000010000",
			6552 => "0001101101111100001000",
			6553 => "0011000100010100000100",
			6554 => "0000000110011101010001",
			6555 => "0000000110011101010001",
			6556 => "0011000111111000000100",
			6557 => "0000000110011101010001",
			6558 => "0000000110011101010001",
			6559 => "0011110110110100001000",
			6560 => "0001010110000100000100",
			6561 => "0000000110011101010001",
			6562 => "1111110110011101010001",
			6563 => "0001101100011000000100",
			6564 => "0000001110011101010001",
			6565 => "0000000110011101010001",
			6566 => "0000011100110100010000",
			6567 => "0001110100010100001000",
			6568 => "0001000011010100000100",
			6569 => "1111111110011101010001",
			6570 => "0000001110011101010001",
			6571 => "0010111100001000000100",
			6572 => "0000001110011101010001",
			6573 => "0000000110011101010001",
			6574 => "0010010111100100001000",
			6575 => "0001100100110100000100",
			6576 => "1111110110011101010001",
			6577 => "1111111110011101010001",
			6578 => "0010000110001000000100",
			6579 => "1111111110011101010001",
			6580 => "0000000110011101010001",
			6581 => "0001101100011000100000",
			6582 => "0001010000001100010000",
			6583 => "0000111001110000001000",
			6584 => "0000010110000000000100",
			6585 => "1111111110011101010001",
			6586 => "0000001110011101010001",
			6587 => "0001010011011100000100",
			6588 => "1111111110011101010001",
			6589 => "0000000110011101010001",
			6590 => "0001111001110000001000",
			6591 => "0010001001101000000100",
			6592 => "0000000110011101010001",
			6593 => "0000001110011101010001",
			6594 => "0000110111001000000100",
			6595 => "1111111110011101010001",
			6596 => "0000000110011101010001",
			6597 => "0010011101101000010000",
			6598 => "0001001111100000001000",
			6599 => "0010000010101000000100",
			6600 => "0000000110011101010001",
			6601 => "1111111110011101010001",
			6602 => "0010010110101000000100",
			6603 => "0000000110011101010001",
			6604 => "0000000110011101010001",
			6605 => "0001011010111100001000",
			6606 => "0001000011001100000100",
			6607 => "0000000110011101010001",
			6608 => "0000000110011101010001",
			6609 => "0000010010001100000100",
			6610 => "0000000110011101010001",
			6611 => "0000000110011101010001",
			6612 => "0011101000000010011000",
			6613 => "0010011111001101011000",
			6614 => "0010110101101100111100",
			6615 => "0011100100001000100000",
			6616 => "0010011011101000010000",
			6617 => "0010110101101100001000",
			6618 => "0010010111100100000100",
			6619 => "0000000110100101011101",
			6620 => "0000000110100101011101",
			6621 => "0001101100011000000100",
			6622 => "0000001110100101011101",
			6623 => "1111111110100101011101",
			6624 => "0001000011110000001000",
			6625 => "0000010010001100000100",
			6626 => "0000000110100101011101",
			6627 => "1111111110100101011101",
			6628 => "0011111101000100000100",
			6629 => "0000001110100101011101",
			6630 => "1111111110100101011101",
			6631 => "0011111101000100010000",
			6632 => "0001111000111000001000",
			6633 => "0000000010011000000100",
			6634 => "0000000110100101011101",
			6635 => "1111111110100101011101",
			6636 => "0010111101100000000100",
			6637 => "0000000110100101011101",
			6638 => "0000001110100101011101",
			6639 => "0011100100001000000100",
			6640 => "0000001110100101011101",
			6641 => "0000000000111000000100",
			6642 => "0000000110100101011101",
			6643 => "0000000110100101011101",
			6644 => "0001000100001100001100",
			6645 => "0001101100011000001000",
			6646 => "0011010100011000000100",
			6647 => "0000000110100101011101",
			6648 => "0000000110100101011101",
			6649 => "1111110110100101011101",
			6650 => "0001000011101100000100",
			6651 => "0000001110100101011101",
			6652 => "0011001000111000000100",
			6653 => "1111111110100101011101",
			6654 => "0000011100110100000100",
			6655 => "0000000110100101011101",
			6656 => "0000001110100101011101",
			6657 => "0000000000110000110000",
			6658 => "0001111000111000010100",
			6659 => "0010110011011100001000",
			6660 => "0000111001001000000100",
			6661 => "0000000110100101011101",
			6662 => "1111111110100101011101",
			6663 => "0000011001111000000100",
			6664 => "0000010110100101011101",
			6665 => "0000011001111000000100",
			6666 => "0000000110100101011101",
			6667 => "0000001110100101011101",
			6668 => "0010001011010100010000",
			6669 => "0000101001010000001000",
			6670 => "0011100100011000000100",
			6671 => "0000001110100101011101",
			6672 => "0000000110100101011101",
			6673 => "0011010011100000000100",
			6674 => "1111111110100101011101",
			6675 => "0000000110100101011101",
			6676 => "0001001010110100001000",
			6677 => "0001101101011000000100",
			6678 => "0000001110100101011101",
			6679 => "0000000110100101011101",
			6680 => "1111111110100101011101",
			6681 => "0011010110100100001100",
			6682 => "0001101001100100000100",
			6683 => "0000001110100101011101",
			6684 => "0001101111000000000100",
			6685 => "0000000110100101011101",
			6686 => "0000000110100101011101",
			6687 => "1111111110100101011101",
			6688 => "0011111110110100111100",
			6689 => "0011001000111100100000",
			6690 => "0010111000111000000100",
			6691 => "0000001110100101011101",
			6692 => "0000101100010100001100",
			6693 => "0001101010011000001000",
			6694 => "0011111101000100000100",
			6695 => "0000000110100101011101",
			6696 => "1111111110100101011101",
			6697 => "0000001110100101011101",
			6698 => "0001111001110000001000",
			6699 => "0011000000101000000100",
			6700 => "0000000110100101011101",
			6701 => "1111111110100101011101",
			6702 => "0010011001011000000100",
			6703 => "0000000110100101011101",
			6704 => "1111111110100101011101",
			6705 => "0000111010011100000100",
			6706 => "0000001110100101011101",
			6707 => "0011001000111100001000",
			6708 => "0011010110100100000100",
			6709 => "0000001110100101011101",
			6710 => "1111111110100101011101",
			6711 => "0011001000111000001000",
			6712 => "0011111110010000000100",
			6713 => "1111111110100101011101",
			6714 => "0000000110100101011101",
			6715 => "0000011001111000000100",
			6716 => "0000001110100101011101",
			6717 => "0000000110100101011101",
			6718 => "0000111100010100010100",
			6719 => "0010011100011000001100",
			6720 => "0001101000010000000100",
			6721 => "0000001110100101011101",
			6722 => "0010011110010100000100",
			6723 => "0000000110100101011101",
			6724 => "0000001110100101011101",
			6725 => "0001110011100000000100",
			6726 => "1111111110100101011101",
			6727 => "0000000110100101011101",
			6728 => "0001000011001100000100",
			6729 => "1111111110100101011101",
			6730 => "0000010101011100001100",
			6731 => "0010001000110000000100",
			6732 => "1111111110100101011101",
			6733 => "0000001000111000000100",
			6734 => "0000000110100101011101",
			6735 => "0000000110100101011101",
			6736 => "0010000001110100001000",
			6737 => "0011111011110000000100",
			6738 => "0000001110100101011101",
			6739 => "0000000110100101011101",
			6740 => "0000101101001000000100",
			6741 => "0000000110100101011101",
			6742 => "0000001110100101011101",
			6743 => "0001000000101110111000",
			6744 => "0001010100011001100100",
			6745 => "0010011111001100111100",
			6746 => "0000111011000000100000",
			6747 => "0010011101101000010000",
			6748 => "0011100110000100001000",
			6749 => "0010011101101000000100",
			6750 => "0000000110101101000001",
			6751 => "0000000110101101000001",
			6752 => "0000101001100000000100",
			6753 => "1111111110101101000001",
			6754 => "0000000110101101000001",
			6755 => "0011101101111000001000",
			6756 => "0010111001110000000100",
			6757 => "0000000110101101000001",
			6758 => "0000000110101101000001",
			6759 => "0001100100110100000100",
			6760 => "0000001110101101000001",
			6761 => "0000000110101101000001",
			6762 => "0001101010011000010000",
			6763 => "0001010100001000001000",
			6764 => "0010111001110000000100",
			6765 => "0000001110101101000001",
			6766 => "0000010110101101000001",
			6767 => "0001111000111000000100",
			6768 => "1111111110101101000001",
			6769 => "0000000110101101000001",
			6770 => "0000010010001100000100",
			6771 => "0000001110101101000001",
			6772 => "0011001000111000000100",
			6773 => "1111111110101101000001",
			6774 => "0000000110101101000001",
			6775 => "0011100100011000010100",
			6776 => "0011001100001000000100",
			6777 => "0000010110101101000001",
			6778 => "0010001001101000001000",
			6779 => "0010110101101100000100",
			6780 => "1111111110101101000001",
			6781 => "0000001110101101000001",
			6782 => "0011001000111000000100",
			6783 => "0000001110101101000001",
			6784 => "0000000110101101000001",
			6785 => "0011000000101000000100",
			6786 => "0000001110101101000001",
			6787 => "0011001000111100001000",
			6788 => "0001001001001100000100",
			6789 => "1111111110101101000001",
			6790 => "0000001110101101000001",
			6791 => "0001111001110000000100",
			6792 => "0000000110101101000001",
			6793 => "0000001110101101000001",
			6794 => "0010001001101000011000",
			6795 => "0010010100110100010100",
			6796 => "0010111100101100000100",
			6797 => "1111111110101101000001",
			6798 => "0011100001101000001000",
			6799 => "0001000110111000000100",
			6800 => "0000000110101101000001",
			6801 => "1111111110101101000001",
			6802 => "0010100110011000000100",
			6803 => "0000000110101101000001",
			6804 => "1111111110101101000001",
			6805 => "1111111110101101000001",
			6806 => "0011001100110000100000",
			6807 => "0001001000001000010000",
			6808 => "0010111110001100001000",
			6809 => "0000100111011000000100",
			6810 => "1111111110101101000001",
			6811 => "0000000110101101000001",
			6812 => "0000011101101000000100",
			6813 => "0000001110101101000001",
			6814 => "0000000110101101000001",
			6815 => "0011101001001000001000",
			6816 => "0010111110001100000100",
			6817 => "0000000110101101000001",
			6818 => "1111110110101101000001",
			6819 => "0011110100101000000100",
			6820 => "0000001110101101000001",
			6821 => "0000000110101101000001",
			6822 => "0001001110111000010000",
			6823 => "0001100101010000001000",
			6824 => "0001001101001000000100",
			6825 => "0000001110101101000001",
			6826 => "0000010110101101000001",
			6827 => "0010110110100000000100",
			6828 => "1111111110101101000001",
			6829 => "0000001110101101000001",
			6830 => "0010001111001000000100",
			6831 => "1111111110101101000001",
			6832 => "0011000110000100000100",
			6833 => "0000000110101101000001",
			6834 => "0000000110101101000001",
			6835 => "0010001101010000011100",
			6836 => "0000010110000000001100",
			6837 => "0001000110110000001000",
			6838 => "0010011110100000000100",
			6839 => "0000000110101101000001",
			6840 => "0000001110101101000001",
			6841 => "1111111110101101000001",
			6842 => "0011111001010100000100",
			6843 => "1111110110101101000001",
			6844 => "0001101011001100001000",
			6845 => "0010100101000100000100",
			6846 => "0000000110101101000001",
			6847 => "0000000110101101000001",
			6848 => "1111111110101101000001",
			6849 => "0001000101100000011100",
			6850 => "0011000111111000001000",
			6851 => "0011000111111000000100",
			6852 => "0000001110101101000001",
			6853 => "1111111110101101000001",
			6854 => "0010110000101000000100",
			6855 => "0000001110101101000001",
			6856 => "0000100010010100001000",
			6857 => "0000101100010000000100",
			6858 => "0000000110101101000001",
			6859 => "1111111110101101000001",
			6860 => "0001000011111000000100",
			6861 => "0000001110101101000001",
			6862 => "0000000110101101000001",
			6863 => "1111111110101101000001",
			6864 => "0010001011010110001000",
			6865 => "0000000011010001010100",
			6866 => "0001101010011000111000",
			6867 => "0000011001111000011100",
			6868 => "0001100100110100010000",
			6869 => "0010110011011100001000",
			6870 => "0000010010001100000100",
			6871 => "0000000110110101111101",
			6872 => "0000000110110101111101",
			6873 => "0000010010001100000100",
			6874 => "0000001110110101111101",
			6875 => "0000000110110101111101",
			6876 => "0000001101010000000100",
			6877 => "0000010110110101111101",
			6878 => "0000000011111100000100",
			6879 => "0000000110110101111101",
			6880 => "1111111110110101111101",
			6881 => "0001100100110100010000",
			6882 => "0000011001111000001000",
			6883 => "0001011010111100000100",
			6884 => "1111111110110101111101",
			6885 => "0000000110110101111101",
			6886 => "0010110101101100000100",
			6887 => "0000001110110101111101",
			6888 => "0000000110110101111101",
			6889 => "0001000011110000001000",
			6890 => "0001111101100000000100",
			6891 => "1111111110110101111101",
			6892 => "0000000110110101111101",
			6893 => "0000000110110101111101",
			6894 => "0010000001010100000100",
			6895 => "1111111110110101111101",
			6896 => "0011110110100000001000",
			6897 => "0001001000000100000100",
			6898 => "0000000110110101111101",
			6899 => "0000001110110101111101",
			6900 => "0010000001010100001000",
			6901 => "0000001000101100000100",
			6902 => "0000000110110101111101",
			6903 => "0000100110110101111101",
			6904 => "0011101000000000000100",
			6905 => "1111111110110101111101",
			6906 => "0000000110110101111101",
			6907 => "0001110111111000010100",
			6908 => "0000111100001000001000",
			6909 => "0010001001101000000100",
			6910 => "0000000110110101111101",
			6911 => "0000001110110101111101",
			6912 => "0001011001110000001000",
			6913 => "0011000000111000000100",
			6914 => "0000000110110101111101",
			6915 => "0000000110110101111101",
			6916 => "1111111110110101111101",
			6917 => "0000101111010000010000",
			6918 => "0010001001101000001000",
			6919 => "0001011101100000000100",
			6920 => "0000001110110101111101",
			6921 => "0000000110110101111101",
			6922 => "0011110001011000000100",
			6923 => "0000001110110101111101",
			6924 => "0000001110110101111101",
			6925 => "0000011100110100001100",
			6926 => "0010001001101000000100",
			6927 => "0000001110110101111101",
			6928 => "0001111100001000000100",
			6929 => "0000000110110101111101",
			6930 => "0000000110110101111101",
			6931 => "1111111110110101111101",
			6932 => "0000111011000101001100",
			6933 => "0001000100001100100000",
			6934 => "0010101010110000010100",
			6935 => "0011111011000000001000",
			6936 => "0011101010101100000100",
			6937 => "0000001110110101111101",
			6938 => "1111111110110101111101",
			6939 => "0001011000111100000100",
			6940 => "0000000110110101111101",
			6941 => "0010100110011000000100",
			6942 => "0000000110110101111101",
			6943 => "0000001110110101111101",
			6944 => "0011101111000100001000",
			6945 => "0001011001110000000100",
			6946 => "0000001110110101111101",
			6947 => "1111111110110101111101",
			6948 => "0000001110110101111101",
			6949 => "0000000100010100001100",
			6950 => "0010110100010100001000",
			6951 => "0000111110111100000100",
			6952 => "0000000110110101111101",
			6953 => "1111110110110101111101",
			6954 => "0000000110110101111101",
			6955 => "0000010110000000010000",
			6956 => "0011111110110000001000",
			6957 => "0001000110110000000100",
			6958 => "0000001110110101111101",
			6959 => "0000000110110101111101",
			6960 => "0011110000011100000100",
			6961 => "1111111110110101111101",
			6962 => "0000001110110101111101",
			6963 => "0001000000100000001000",
			6964 => "0001011001110000000100",
			6965 => "0000001110110101111101",
			6966 => "0000000110110101111101",
			6967 => "0010001101010000000100",
			6968 => "1111111110110101111101",
			6969 => "0000000110110101111101",
			6970 => "0011111000011000001100",
			6971 => "0011001011000100001000",
			6972 => "0011000111111000000100",
			6973 => "1111111110110101111101",
			6974 => "1111111110110101111101",
			6975 => "0000000110110101111101",
			6976 => "0000111100001000100000",
			6977 => "0000010110000000010000",
			6978 => "0001010011011100001000",
			6979 => "0001011000111100000100",
			6980 => "0000000110110101111101",
			6981 => "1111111110110101111101",
			6982 => "0010111011000000000100",
			6983 => "0000001110110101111101",
			6984 => "0000000110110101111101",
			6985 => "0000100111100000001000",
			6986 => "0011000111111000000100",
			6987 => "0000000110110101111101",
			6988 => "0000001110110101111101",
			6989 => "0000010110000000000100",
			6990 => "0000001110110101111101",
			6991 => "0000000110110101111101",
			6992 => "0011110110110100010000",
			6993 => "0011100111111000001000",
			6994 => "0000000011010000000100",
			6995 => "1111111110110101111101",
			6996 => "0000000110110101111101",
			6997 => "0011000000101000000100",
			6998 => "1111111110110101111101",
			6999 => "0000000110110101111101",
			7000 => "0011101100001000001000",
			7001 => "0001111011000100000100",
			7002 => "0000000110110101111101",
			7003 => "0000000110110101111101",
			7004 => "0011111011110100000100",
			7005 => "0000000110110101111101",
			7006 => "0000000110110101111101",
			7007 => "0001011010111110101100",
			7008 => "0011000000101001001100",
			7009 => "0011000100010100110000",
			7010 => "0010011011101000100000",
			7011 => "0001110100000000010000",
			7012 => "0001111100001000001000",
			7013 => "0001110000101000000100",
			7014 => "0000000110111110110001",
			7015 => "0000000110111110110001",
			7016 => "0011000100010100000100",
			7017 => "0000000110111110110001",
			7018 => "0000001110111110110001",
			7019 => "0001010100001000001000",
			7020 => "0001100100110100000100",
			7021 => "0000000110111110110001",
			7022 => "1111111110111110110001",
			7023 => "0000000000110000000100",
			7024 => "0000001110111110110001",
			7025 => "0000000110111110110001",
			7026 => "0001100100110100000100",
			7027 => "1111111110111110110001",
			7028 => "0011101010111100000100",
			7029 => "0000001110111110110001",
			7030 => "0011011010111100000100",
			7031 => "0000000110111110110001",
			7032 => "0000001110111110110001",
			7033 => "0001110000101000001100",
			7034 => "0000100111100000000100",
			7035 => "0000000110111110110001",
			7036 => "0001001001001100000100",
			7037 => "1111111110111110110001",
			7038 => "1111111110111110110001",
			7039 => "0011101100101100001100",
			7040 => "0011111010010100001000",
			7041 => "0000011100110100000100",
			7042 => "0000000110111110110001",
			7043 => "1111111110111110110001",
			7044 => "0000001110111110110001",
			7045 => "1111111110111110110001",
			7046 => "0011000000101000101000",
			7047 => "0001110100010100001000",
			7048 => "0001000101010100000100",
			7049 => "1111111110111110110001",
			7050 => "0000000110111110110001",
			7051 => "0010110100000000010000",
			7052 => "0010111100001000001000",
			7053 => "0001111011000100000100",
			7054 => "0000001110111110110001",
			7055 => "0000000110111110110001",
			7056 => "0000100011001000000100",
			7057 => "0000001110111110110001",
			7058 => "0000000110111110110001",
			7059 => "0010101001000100001000",
			7060 => "0001001000110100000100",
			7061 => "0000000110111110110001",
			7062 => "0000001110111110110001",
			7063 => "0000101110010000000100",
			7064 => "0000000110111110110001",
			7065 => "0000000110111110110001",
			7066 => "0011000000101000011000",
			7067 => "0010111100001000001000",
			7068 => "0001011100101100000100",
			7069 => "0000000110111110110001",
			7070 => "0000001110111110110001",
			7071 => "0001011100101000001000",
			7072 => "0000000111111000000100",
			7073 => "1111111110111110110001",
			7074 => "0000000110111110110001",
			7075 => "0001110100000000000100",
			7076 => "0000001110111110110001",
			7077 => "1111111110111110110001",
			7078 => "0011000100000000010000",
			7079 => "0001110100000000001000",
			7080 => "0001000110001100000100",
			7081 => "1111111110111110110001",
			7082 => "0000000110111110110001",
			7083 => "0010011011101000000100",
			7084 => "0000001110111110110001",
			7085 => "0000000110111110110001",
			7086 => "0001101100011000001000",
			7087 => "0011110010001000000100",
			7088 => "0000000110111110110001",
			7089 => "0000000110111110110001",
			7090 => "0010100110011000000100",
			7091 => "0000001110111110110001",
			7092 => "0000000110111110110001",
			7093 => "0001111000111000100000",
			7094 => "0011001000111100011100",
			7095 => "0001001110100100001000",
			7096 => "0000000111000000000100",
			7097 => "0000000110111110110001",
			7098 => "1111111110111110110001",
			7099 => "0010111101100000001000",
			7100 => "0010011111001100000100",
			7101 => "0000001110111110110001",
			7102 => "0000000110111110110001",
			7103 => "0010011101011100001000",
			7104 => "0010011011101000000100",
			7105 => "1111111110111110110001",
			7106 => "1111111110111110110001",
			7107 => "0000000110111110110001",
			7108 => "0000000110111110110001",
			7109 => "0011110001000000100000",
			7110 => "0011011101010100000100",
			7111 => "1111111110111110110001",
			7112 => "0001001111100000001100",
			7113 => "0011110001000000001000",
			7114 => "0001001001001100000100",
			7115 => "0000000110111110110001",
			7116 => "0000001110111110110001",
			7117 => "0000001110111110110001",
			7118 => "0010011011101000001000",
			7119 => "0001101101011000000100",
			7120 => "1111111110111110110001",
			7121 => "0000001110111110110001",
			7122 => "0001101011001100000100",
			7123 => "1111101110111110110001",
			7124 => "0000000110111110110001",
			7125 => "0011100100011000010100",
			7126 => "0001101011001100001100",
			7127 => "0010011101011100001000",
			7128 => "0010110110000100000100",
			7129 => "1111111110111110110001",
			7130 => "0000000110111110110001",
			7131 => "0000001110111110110001",
			7132 => "0001101001100100000100",
			7133 => "0000001110111110110001",
			7134 => "0000000110111110110001",
			7135 => "0000100110010000001100",
			7136 => "0011011011000000000100",
			7137 => "0000000110111110110001",
			7138 => "0001101011001100000100",
			7139 => "1111111110111110110001",
			7140 => "0000000110111110110001",
			7141 => "0001101010011000001000",
			7142 => "0011001000111100000100",
			7143 => "0000001110111110110001",
			7144 => "0000000110111110110001",
			7145 => "0001111001110000000100",
			7146 => "1111111110111110110001",
			7147 => "0000000110111110110001",
			7148 => "0011000100000010100000",
			7149 => "0001111001110001110000",
			7150 => "0001011010111100111100",
			7151 => "0011000100000000100000",
			7152 => "0000110011100000010000",
			7153 => "0000110100011000001000",
			7154 => "0011010111001000000100",
			7155 => "0000000111000111100101",
			7156 => "0000001111000111100101",
			7157 => "0010111001110000000100",
			7158 => "0000000111000111100101",
			7159 => "1111111111000111100101",
			7160 => "0011000000101000001000",
			7161 => "0010000111000100000100",
			7162 => "1111111111000111100101",
			7163 => "0000000111000111100101",
			7164 => "0001111100001000000100",
			7165 => "1111111111000111100101",
			7166 => "0000001111000111100101",
			7167 => "0001110100000000001100",
			7168 => "0001110100000000001000",
			7169 => "0010010111100100000100",
			7170 => "0000000111000111100101",
			7171 => "0000001111000111100101",
			7172 => "1111111111000111100101",
			7173 => "0010101100011100001000",
			7174 => "0001111000111000000100",
			7175 => "0000001111000111100101",
			7176 => "0000000111000111100101",
			7177 => "0000101001100000000100",
			7178 => "0000001111000111100101",
			7179 => "0000000111000111100101",
			7180 => "0010011101011100100000",
			7181 => "0010111101100000010000",
			7182 => "0011000100000000001000",
			7183 => "0001110100000000000100",
			7184 => "1111111111000111100101",
			7185 => "0000000111000111100101",
			7186 => "0001111000111000000100",
			7187 => "0000001111000111100101",
			7188 => "0000000111000111100101",
			7189 => "0001100100110100001000",
			7190 => "0001001000000100000100",
			7191 => "0000000111000111100101",
			7192 => "0000000111000111100101",
			7193 => "0001000100001100000100",
			7194 => "1111111111000111100101",
			7195 => "0000000111000111100101",
			7196 => "0011000000101000000100",
			7197 => "0000001111000111100101",
			7198 => "0011101000000000001000",
			7199 => "0000100010000000000100",
			7200 => "0000000111000111100101",
			7201 => "0000001111000111100101",
			7202 => "0000101110110100000100",
			7203 => "1111111111000111100101",
			7204 => "0000000111000111100101",
			7205 => "0010000001110100101000",
			7206 => "0001011010111000001100",
			7207 => "0000100101110000000100",
			7208 => "0000000111000111100101",
			7209 => "0010000111000100000100",
			7210 => "0000001111000111100101",
			7211 => "0000000111000111100101",
			7212 => "0011010110100100010000",
			7213 => "0001101101011000001000",
			7214 => "0000101100010100000100",
			7215 => "0000000111000111100101",
			7216 => "0000001111000111100101",
			7217 => "0001001110100100000100",
			7218 => "0000000111000111100101",
			7219 => "1111111111000111100101",
			7220 => "0010011011111100001000",
			7221 => "0000101100010000000100",
			7222 => "0000000111000111100101",
			7223 => "0000001111000111100101",
			7224 => "0000000111000111100101",
			7225 => "0010000010101000000100",
			7226 => "1111111111000111100101",
			7227 => "0000000111000111100101",
			7228 => "0011000100000000011100",
			7229 => "0001011010111000010100",
			7230 => "0010111000111000000100",
			7231 => "0000000111000111100101",
			7232 => "0010101100011100001100",
			7233 => "0000011001111000001000",
			7234 => "0000100100101000000100",
			7235 => "0000000111000111100101",
			7236 => "1111111111000111100101",
			7237 => "0000000111000111100101",
			7238 => "0000000111000111100101",
			7239 => "0011101000011000000100",
			7240 => "0000001111000111100101",
			7241 => "1111111111000111100101",
			7242 => "0011001000111100101000",
			7243 => "0011001000111100011000",
			7244 => "0001111001110000010000",
			7245 => "0011101101100000001000",
			7246 => "0000010010001100000100",
			7247 => "0000000111000111100101",
			7248 => "0000001111000111100101",
			7249 => "0011101100101100000100",
			7250 => "1111111111000111100101",
			7251 => "0000000111000111100101",
			7252 => "0010000111000100000100",
			7253 => "1111111111000111100101",
			7254 => "0000000111000111100101",
			7255 => "0000011001111000000100",
			7256 => "0000001111000111100101",
			7257 => "0011101001001000000100",
			7258 => "0000000111000111100101",
			7259 => "0010100001010000000100",
			7260 => "0000001111000111100101",
			7261 => "0000000111000111100101",
			7262 => "0001101010011000011100",
			7263 => "0001000000010100001100",
			7264 => "0010001111001000001000",
			7265 => "0011011110110000000100",
			7266 => "0000000111000111100101",
			7267 => "1111111111000111100101",
			7268 => "1111111111000111100101",
			7269 => "0011011011000000001000",
			7270 => "0000011110100000000100",
			7271 => "0000000111000111100101",
			7272 => "0000001111000111100101",
			7273 => "0001101010011000000100",
			7274 => "0000000111000111100101",
			7275 => "0000000111000111100101",
			7276 => "0000100100101000001100",
			7277 => "0011011001001000001000",
			7278 => "0010110000001100000100",
			7279 => "0000001111000111100101",
			7280 => "0000000111000111100101",
			7281 => "0000000111000111100101",
			7282 => "0010011101101000001000",
			7283 => "0001001101001100000100",
			7284 => "0000001111000111100101",
			7285 => "0000000111000111100101",
			7286 => "0011011010111000000100",
			7287 => "0000000111000111100101",
			7288 => "0000000111000111100101",
			7289 => "0010011001111001111000",
			7290 => "0011000100010100111100",
			7291 => "0011000100010100111000",
			7292 => "0001000001101100011100",
			7293 => "0011101111000100001100",
			7294 => "0010110100010100001000",
			7295 => "0011110111010000000100",
			7296 => "0000000111010001000001",
			7297 => "0000001111010001000001",
			7298 => "0000001111010001000001",
			7299 => "0011110000011100001000",
			7300 => "0000001110111100000100",
			7301 => "0000000111010001000001",
			7302 => "1111111111010001000001",
			7303 => "0011000111111000000100",
			7304 => "0000000111010001000001",
			7305 => "1111111111010001000001",
			7306 => "0010100001010100010000",
			7307 => "0000110010111100001000",
			7308 => "0000110010011000000100",
			7309 => "0000000111010001000001",
			7310 => "1111011111010001000001",
			7311 => "0000001100001000000100",
			7312 => "0000000111010001000001",
			7313 => "1111111111010001000001",
			7314 => "0010100001110000000100",
			7315 => "0000001111010001000001",
			7316 => "0011101011010100000100",
			7317 => "1111111111010001000001",
			7318 => "0000000111010001000001",
			7319 => "0000001111010001000001",
			7320 => "0000110100000000101100",
			7321 => "0000010110000000010100",
			7322 => "0011110101100100001100",
			7323 => "0000010000011000001000",
			7324 => "0011100010101000000100",
			7325 => "0000000111010001000001",
			7326 => "0000000111010001000001",
			7327 => "0000001111010001000001",
			7328 => "0011111011011100000100",
			7329 => "1111111111010001000001",
			7330 => "0000000111010001000001",
			7331 => "0011011100110000010000",
			7332 => "0010010010001100001000",
			7333 => "0011011101100000000100",
			7334 => "1111111111010001000001",
			7335 => "1111110111010001000001",
			7336 => "0010110100010100000100",
			7337 => "1111111111010001000001",
			7338 => "0000001111010001000001",
			7339 => "0001011100110000000100",
			7340 => "0000001111010001000001",
			7341 => "1111111111010001000001",
			7342 => "0011000100010100000100",
			7343 => "1111110111010001000001",
			7344 => "0011101110111100001000",
			7345 => "0011110110110100000100",
			7346 => "0000000111010001000001",
			7347 => "0000001111010001000001",
			7348 => "1111111111010001000001",
			7349 => "0000110101101101001000",
			7350 => "0000110101101100110100",
			7351 => "0000111100110000100000",
			7352 => "0010010111100100010000",
			7353 => "0000011100110100001000",
			7354 => "0001110111111000000100",
			7355 => "0000000111010001000001",
			7356 => "0000000111010001000001",
			7357 => "0001110000101000000100",
			7358 => "0000000111010001000001",
			7359 => "1111111111010001000001",
			7360 => "0000011100110100001000",
			7361 => "0001011101111000000100",
			7362 => "0000001111010001000001",
			7363 => "0000000111010001000001",
			7364 => "0010010111100100000100",
			7365 => "0000000111010001000001",
			7366 => "0000001111010001000001",
			7367 => "0001100100110100001100",
			7368 => "0011000100010100001000",
			7369 => "0011000100010100000100",
			7370 => "0000000111010001000001",
			7371 => "0000001111010001000001",
			7372 => "1111111111010001000001",
			7373 => "0011111011110100000100",
			7374 => "1111111111010001000001",
			7375 => "1111111111010001000001",
			7376 => "0010111100001000001100",
			7377 => "0001111011000100000100",
			7378 => "0000001111010001000001",
			7379 => "0011101011000100000100",
			7380 => "0000001111010001000001",
			7381 => "0000001111010001000001",
			7382 => "0011011110001100000100",
			7383 => "0000000111010001000001",
			7384 => "0000001111010001000001",
			7385 => "0010010110101000110000",
			7386 => "0011110101110100010100",
			7387 => "0011111011011100001000",
			7388 => "0001001000011100000100",
			7389 => "1111111111010001000001",
			7390 => "0000000111010001000001",
			7391 => "0001111100001000001000",
			7392 => "0010100001010000000100",
			7393 => "1111111111010001000001",
			7394 => "0000000111010001000001",
			7395 => "1111111111010001000001",
			7396 => "0001011100101100010000",
			7397 => "0011000111111000001000",
			7398 => "0000111100101100000100",
			7399 => "1111111111010001000001",
			7400 => "0000000111010001000001",
			7401 => "0011000100010100000100",
			7402 => "0000000111010001000001",
			7403 => "1111111111010001000001",
			7404 => "0010010110101000000100",
			7405 => "0000000111010001000001",
			7406 => "0011101000111000000100",
			7407 => "0000001111010001000001",
			7408 => "0000000111010001000001",
			7409 => "0011000000101000100000",
			7410 => "0011000000101000010000",
			7411 => "0011000000101000001000",
			7412 => "0010011111001100000100",
			7413 => "0000000111010001000001",
			7414 => "0000001111010001000001",
			7415 => "0001110100000000000100",
			7416 => "0000001111010001000001",
			7417 => "0000000111010001000001",
			7418 => "0011010001111100001000",
			7419 => "0001110100000000000100",
			7420 => "0000000111010001000001",
			7421 => "0000000111010001000001",
			7422 => "0001111000111000000100",
			7423 => "1111111111010001000001",
			7424 => "0000000111010001000001",
			7425 => "0001111100001000010000",
			7426 => "0001111100001000001000",
			7427 => "0010111100001000000100",
			7428 => "0000001111010001000001",
			7429 => "0000000111010001000001",
			7430 => "0011000000101000000100",
			7431 => "0000001111010001000001",
			7432 => "0000000111010001000001",
			7433 => "0010011101101000001000",
			7434 => "0000011100110100000100",
			7435 => "0000000111010001000001",
			7436 => "0000000111010001000001",
			7437 => "0000011100110100000100",
			7438 => "0000001111010001000001",
			7439 => "0000000111010001000001",
			7440 => "0011000111111011000000",
			7441 => "0010010110101001101100",
			7442 => "0000111001110000111100",
			7443 => "0010011001111000100000",
			7444 => "0000011110100000010000",
			7445 => "0001100111101000001000",
			7446 => "0010110100010100000100",
			7447 => "1111111111011011000101",
			7448 => "0000000111011011000101",
			7449 => "0000010110000000000100",
			7450 => "0000000111011011000101",
			7451 => "0000000111011011000101",
			7452 => "0010110100010100001000",
			7453 => "0001010011011100000100",
			7454 => "1111111111011011000101",
			7455 => "0000000111011011000101",
			7456 => "0001110100010100000100",
			7457 => "0000001111011011000101",
			7458 => "0000000111011011000101",
			7459 => "0001000011110000001100",
			7460 => "0011100000110000001000",
			7461 => "0000111100001000000100",
			7462 => "0000001111011011000101",
			7463 => "0000000111011011000101",
			7464 => "1111111111011011000101",
			7465 => "0010100001010000001000",
			7466 => "0010110100010100000100",
			7467 => "0000000111011011000101",
			7468 => "0000001111011011000101",
			7469 => "0000000100010100000100",
			7470 => "0000000111011011000101",
			7471 => "0000001111011011000101",
			7472 => "0000100101110000010100",
			7473 => "0001101101111100001100",
			7474 => "0000011110100000000100",
			7475 => "1111111111011011000101",
			7476 => "0000100101001000000100",
			7477 => "1111111111011011000101",
			7478 => "0000001111011011000101",
			7479 => "0001110100010100000100",
			7480 => "1111111111011011000101",
			7481 => "1111111111011011000101",
			7482 => "0010100001010000010000",
			7483 => "0000110101101100001000",
			7484 => "0001011101100000000100",
			7485 => "0000000111011011000101",
			7486 => "0000001111011011000101",
			7487 => "0001001001001100000100",
			7488 => "1111111111011011000101",
			7489 => "0000001111011011000101",
			7490 => "0010101100011100001000",
			7491 => "0011000111111000000100",
			7492 => "1111111111011011000101",
			7493 => "0000000111011011000101",
			7494 => "0000001111011011000101",
			7495 => "0001011100110000011000",
			7496 => "0010110000101000010000",
			7497 => "0011000111111000001100",
			7498 => "0011100000101000001000",
			7499 => "0000100010011100000100",
			7500 => "0000001111011011000101",
			7501 => "0000001111011011000101",
			7502 => "0000000111011011000101",
			7503 => "0000000111011011000101",
			7504 => "0010010110101000000100",
			7505 => "0000001111011011000101",
			7506 => "0000010111011011000101",
			7507 => "0010101001000100100000",
			7508 => "0001001000110100010000",
			7509 => "0010101000100100001000",
			7510 => "0001000010010100000100",
			7511 => "0000000111011011000101",
			7512 => "0000001111011011000101",
			7513 => "0011000111111000000100",
			7514 => "0000000111011011000101",
			7515 => "1111111111011011000101",
			7516 => "0000011100110100001000",
			7517 => "0000110110000100000100",
			7518 => "0000001111011011000101",
			7519 => "0000000111011011000101",
			7520 => "0001011110001100000100",
			7521 => "0000010111011011000101",
			7522 => "0000000111011011000101",
			7523 => "0011000111111000001100",
			7524 => "0001011100101100001000",
			7525 => "0010000110001000000100",
			7526 => "0000000111011011000101",
			7527 => "1111111111011011000101",
			7528 => "0000001111011011000101",
			7529 => "0000011100110100001000",
			7530 => "0010100110011000000100",
			7531 => "0000000111011011000101",
			7532 => "0000001111011011000101",
			7533 => "0011100000101000000100",
			7534 => "1111111111011011000101",
			7535 => "0000000111011011000101",
			7536 => "0011000100010100111100",
			7537 => "0001001000001000010100",
			7538 => "0000011100110100001100",
			7539 => "0001110100010100000100",
			7540 => "1111111111011011000101",
			7541 => "0001110000101000000100",
			7542 => "0000000111011011000101",
			7543 => "0000001111011011000101",
			7544 => "0011000111111000000100",
			7545 => "0000000111011011000101",
			7546 => "1111111111011011000101",
			7547 => "0000001011000100011000",
			7548 => "0011100100010100001100",
			7549 => "0000100110100000000100",
			7550 => "1111111111011011000101",
			7551 => "0010000111000100000100",
			7552 => "0000000111011011000101",
			7553 => "1111111111011011000101",
			7554 => "0000100011001000000100",
			7555 => "1111111111011011000101",
			7556 => "0011101001110000000100",
			7557 => "0000000111011011000101",
			7558 => "1111111111011011000101",
			7559 => "0010001010101100000100",
			7560 => "0000001111011011000101",
			7561 => "0000101100100100001000",
			7562 => "0010010000011000000100",
			7563 => "0000000111011011000101",
			7564 => "0000001111011011000101",
			7565 => "1111111111011011000101",
			7566 => "0001011001110000001000",
			7567 => "0000000110000100000100",
			7568 => "0000001111011011000101",
			7569 => "0000000111011011000101",
			7570 => "0001111000111000100000",
			7571 => "0001110100000000010000",
			7572 => "0001110100000000001000",
			7573 => "0001111100001000000100",
			7574 => "0000000111011011000101",
			7575 => "0000000111011011000101",
			7576 => "0001110100000000000100",
			7577 => "0000000111011011000101",
			7578 => "0000001111011011000101",
			7579 => "0010110011011100001000",
			7580 => "0000000011111100000100",
			7581 => "0000000111011011000101",
			7582 => "1111111111011011000101",
			7583 => "0001001001001100000100",
			7584 => "0000000111011011000101",
			7585 => "0000001111011011000101",
			7586 => "0000111000011000010000",
			7587 => "0001101100011000001000",
			7588 => "0010010111100100000100",
			7589 => "1111111111011011000101",
			7590 => "0000000111011011000101",
			7591 => "0001011000000000000100",
			7592 => "0000000111011011000101",
			7593 => "1111111111011011000101",
			7594 => "0001111101100000001000",
			7595 => "0000010110101000000100",
			7596 => "0000000111011011000101",
			7597 => "1111111111011011000101",
			7598 => "0011101110110000000100",
			7599 => "1111111111011011000101",
			7600 => "0000000111011011000101",
			7601 => "0010101010110010010000",
			7602 => "0010000111000101101100",
			7603 => "0000101110110100111000",
			7604 => "0010110111111000011000",
			7605 => "0010111110111100001100",
			7606 => "0010111110111100001000",
			7607 => "0010101001000100000100",
			7608 => "1111111111100101010001",
			7609 => "0000000111100101010001",
			7610 => "1111111111100101010001",
			7611 => "0010000001110000000100",
			7612 => "1111111111100101010001",
			7613 => "0000100101110000000100",
			7614 => "0000001111100101010001",
			7615 => "0000000111100101010001",
			7616 => "0010101001000100010000",
			7617 => "0010001011010100001000",
			7618 => "0000010110000000000100",
			7619 => "1111111111100101010001",
			7620 => "0000000111100101010001",
			7621 => "0010011101101000000100",
			7622 => "0000000111100101010001",
			7623 => "0000010111100101010001",
			7624 => "0000100111111100001000",
			7625 => "0000000010111100000100",
			7626 => "0000001111100101010001",
			7627 => "0000000111100101010001",
			7628 => "0010001111001000000100",
			7629 => "0000000111100101010001",
			7630 => "0000000111100101010001",
			7631 => "0010001001101000010100",
			7632 => "0010001001101000010000",
			7633 => "0010110100001000001000",
			7634 => "0000010010001100000100",
			7635 => "0000000111100101010001",
			7636 => "0000001111100101010001",
			7637 => "0001001100001100000100",
			7638 => "1111111111100101010001",
			7639 => "0000000111100101010001",
			7640 => "1111111111100101010001",
			7641 => "0010100110011000010000",
			7642 => "0010101001000100001000",
			7643 => "0010001001101000000100",
			7644 => "0000000111100101010001",
			7645 => "0000000111100101010001",
			7646 => "0010010111101000000100",
			7647 => "0000001111100101010001",
			7648 => "0000000111100101010001",
			7649 => "0010100001010000001000",
			7650 => "0001001000001000000100",
			7651 => "0000000111100101010001",
			7652 => "1111111111100101010001",
			7653 => "0000101100000000000100",
			7654 => "0000000111100101010001",
			7655 => "0000001111100101010001",
			7656 => "0001000000010100010000",
			7657 => "0010100001010000001000",
			7658 => "0011000111111000000100",
			7659 => "0000000111100101010001",
			7660 => "0000001111100101010001",
			7661 => "0000111000111100000100",
			7662 => "0000001111100101010001",
			7663 => "0000000111100101010001",
			7664 => "0000001110111100000100",
			7665 => "1111111111100101010001",
			7666 => "0010011001111000001100",
			7667 => "0001110100010100001000",
			7668 => "0010011100110100000100",
			7669 => "0000000111100101010001",
			7670 => "0000001111100101010001",
			7671 => "1111111111100101010001",
			7672 => "0000001111100101010001",
			7673 => "0001000000010101010000",
			7674 => "0000000111111000111100",
			7675 => "0010000111000100100000",
			7676 => "0010000111000100010000",
			7677 => "0001001001001100001000",
			7678 => "0001001010110100000100",
			7679 => "0000000111100101010001",
			7680 => "0000000111100101010001",
			7681 => "0001111100001000000100",
			7682 => "0000000111100101010001",
			7683 => "0000000111100101010001",
			7684 => "0000101100010100001000",
			7685 => "0001111011000100000100",
			7686 => "0000001111100101010001",
			7687 => "0000000111100101010001",
			7688 => "0001001010110100000100",
			7689 => "1111111111100101010001",
			7690 => "0000001111100101010001",
			7691 => "0001001010110100001100",
			7692 => "0011000000101000000100",
			7693 => "1111111111100101010001",
			7694 => "0000000000110000000100",
			7695 => "0000000111100101010001",
			7696 => "0000001111100101010001",
			7697 => "0001010101101100001000",
			7698 => "0010000111000100000100",
			7699 => "0000001111100101010001",
			7700 => "0000000111100101010001",
			7701 => "0010011011101000000100",
			7702 => "1111111111100101010001",
			7703 => "0000000111100101010001",
			7704 => "0000011110100000000100",
			7705 => "0000000111100101010001",
			7706 => "0001000000010100001100",
			7707 => "0011101110001100001000",
			7708 => "0010101100011100000100",
			7709 => "0000001111100101010001",
			7710 => "0000001111100101010001",
			7711 => "0000000111100101010001",
			7712 => "0000000111100101010001",
			7713 => "0010010110101000110000",
			7714 => "0000011100110100100000",
			7715 => "0000011110100000010000",
			7716 => "0000001011000100001000",
			7717 => "0001001111100000000100",
			7718 => "0000000111100101010001",
			7719 => "1111111111100101010001",
			7720 => "0001000010100100000100",
			7721 => "0000000111100101010001",
			7722 => "0000000111100101010001",
			7723 => "0001011100110000001000",
			7724 => "0001011100110000000100",
			7725 => "0000001111100101010001",
			7726 => "1111111111100101010001",
			7727 => "0011100000101000000100",
			7728 => "0000001111100101010001",
			7729 => "0000000111100101010001",
			7730 => "0010111000111100001100",
			7731 => "0011101000111000001000",
			7732 => "0011111001010100000100",
			7733 => "1111111111100101010001",
			7734 => "0000000111100101010001",
			7735 => "1111111111100101010001",
			7736 => "0000001111100101010001",
			7737 => "0011111110101100011100",
			7738 => "0011110001001000010000",
			7739 => "0001001011100000001000",
			7740 => "0011111001010100000100",
			7741 => "0000000111100101010001",
			7742 => "1111111111100101010001",
			7743 => "0011111010010100000100",
			7744 => "1111111111100101010001",
			7745 => "0000000111100101010001",
			7746 => "0010101010110000000100",
			7747 => "0000000111100101010001",
			7748 => "0010100101000100000100",
			7749 => "0000001111100101010001",
			7750 => "0000000111100101010001",
			7751 => "0000001110111100001100",
			7752 => "0010110011011100000100",
			7753 => "0000001111100101010001",
			7754 => "0011001000111000000100",
			7755 => "1111111111100101010001",
			7756 => "0000000111100101010001",
			7757 => "0001000100001100001000",
			7758 => "0001110100000000000100",
			7759 => "1111111111100101010001",
			7760 => "0000000111100101010001",
			7761 => "0010101100011100000100",
			7762 => "0000000111100101010001",
			7763 => "0000000111100101010001",
			7764 => "0010010110101011000100",
			7765 => "0000110011011101101100",
			7766 => "0011110110110101000000",
			7767 => "0011100011111100100000",
			7768 => "0000110000101000010000",
			7769 => "0000011110100000001000",
			7770 => "0010010010001100000100",
			7771 => "0000000111101111010101",
			7772 => "0000000111101111010101",
			7773 => "0001100111101000000100",
			7774 => "0000000111101111010101",
			7775 => "1111110111101111010101",
			7776 => "0011110001011000001000",
			7777 => "0010101100011100000100",
			7778 => "0000001111101111010101",
			7779 => "0000000111101111010101",
			7780 => "0001101101111100000100",
			7781 => "1111111111101111010101",
			7782 => "0000001111101111010101",
			7783 => "0010010010001100010000",
			7784 => "0000110000101000001000",
			7785 => "0010000001110100000100",
			7786 => "0000001111101111010101",
			7787 => "1111111111101111010101",
			7788 => "0011110101100100000100",
			7789 => "1111111111101111010101",
			7790 => "0000000111101111010101",
			7791 => "0011111010011100001000",
			7792 => "0001100111101000000100",
			7793 => "0000000111101111010101",
			7794 => "1111111111101111010101",
			7795 => "0001110111111000000100",
			7796 => "1111111111101111010101",
			7797 => "0000000111101111010101",
			7798 => "0010011001111000011000",
			7799 => "0000111000111000001100",
			7800 => "0001011101100000001000",
			7801 => "0000010110000000000100",
			7802 => "0000000111101111010101",
			7803 => "0000001111101111010101",
			7804 => "1111111111101111010101",
			7805 => "0011100000110000000100",
			7806 => "1111110111101111010101",
			7807 => "0011111011110100000100",
			7808 => "1111111111101111010101",
			7809 => "0000000111101111010101",
			7810 => "0001011001110000000100",
			7811 => "1111111111101111010101",
			7812 => "0001101101111100001000",
			7813 => "0010011001111000000100",
			7814 => "0000000111101111010101",
			7815 => "0000001111101111010101",
			7816 => "0011100100010100000100",
			7817 => "0000001111101111010101",
			7818 => "0000000111101111010101",
			7819 => "0000101010001000110000",
			7820 => "0010111011000100010100",
			7821 => "0000111101100000001000",
			7822 => "0000000000110000000100",
			7823 => "1111111111101111010101",
			7824 => "0000000111101111010101",
			7825 => "0001110100010100001000",
			7826 => "0011101011000100000100",
			7827 => "0000001111101111010101",
			7828 => "1111111111101111010101",
			7829 => "0000001111101111010101",
			7830 => "0001011100101100010000",
			7831 => "0001111011000100001000",
			7832 => "0001011100110000000100",
			7833 => "1111110111101111010101",
			7834 => "1111111111101111010101",
			7835 => "0001110000101000000100",
			7836 => "0000000111101111010101",
			7837 => "1111111111101111010101",
			7838 => "0010010110101000001000",
			7839 => "0011101011000100000100",
			7840 => "0000000111101111010101",
			7841 => "0000001111101111010101",
			7842 => "1111111111101111010101",
			7843 => "0011000111111000010000",
			7844 => "0000100011001000000100",
			7845 => "0000000111101111010101",
			7846 => "0000101100010100000100",
			7847 => "1111110111101111010101",
			7848 => "0011101100001000000100",
			7849 => "0000001111101111010101",
			7850 => "1111111111101111010101",
			7851 => "0000000000110000001000",
			7852 => "0010001001101000000100",
			7853 => "0000000111101111010101",
			7854 => "0000001111101111010101",
			7855 => "0010110000101000001000",
			7856 => "0001101101111100000100",
			7857 => "0000000111101111010101",
			7858 => "0000001111101111010101",
			7859 => "0001100100110100000100",
			7860 => "0000001111101111010101",
			7861 => "0000000111101111010101",
			7862 => "0000011110100000001100",
			7863 => "0010111100001000001000",
			7864 => "0000110110000100000100",
			7865 => "0000001111101111010101",
			7866 => "0000000111101111010101",
			7867 => "0000010111101111010101",
			7868 => "0011100100010100110100",
			7869 => "0010110000101000010100",
			7870 => "0000000010111100000100",
			7871 => "0000001111101111010101",
			7872 => "0000000000110000001000",
			7873 => "0000011110100000000100",
			7874 => "0000000111101111010101",
			7875 => "1111111111101111010101",
			7876 => "0011100111111000000100",
			7877 => "0000001111101111010101",
			7878 => "0000000111101111010101",
			7879 => "0011110001011000010000",
			7880 => "0000111001110000001000",
			7881 => "0000001101010000000100",
			7882 => "0000000111101111010101",
			7883 => "0000001111101111010101",
			7884 => "0010001111001000000100",
			7885 => "0000000111101111010101",
			7886 => "1111111111101111010101",
			7887 => "0000101110000100001000",
			7888 => "0011110101100100000100",
			7889 => "0000001111101111010101",
			7890 => "0000001111101111010101",
			7891 => "0000000000111000000100",
			7892 => "0000000111101111010101",
			7893 => "0000001111101111010101",
			7894 => "0000101110000100100000",
			7895 => "0001100001111000010000",
			7896 => "0011100100000000001000",
			7897 => "0010100111110100000100",
			7898 => "0000000111101111010101",
			7899 => "0000001111101111010101",
			7900 => "0010100011101000000100",
			7901 => "0000000111101111010101",
			7902 => "0000000111101111010101",
			7903 => "0001100100110100001000",
			7904 => "0000111010111100000100",
			7905 => "0000000111101111010101",
			7906 => "0000000111101111010101",
			7907 => "0000111101111000000100",
			7908 => "1111111111101111010101",
			7909 => "1111111111101111010101",
			7910 => "0001111100001000010000",
			7911 => "0001111100001000001000",
			7912 => "0000100111011000000100",
			7913 => "0000000111101111010101",
			7914 => "1111111111101111010101",
			7915 => "0001111100001000000100",
			7916 => "0000001111101111010101",
			7917 => "0000000111101111010101",
			7918 => "0010110100000000001000",
			7919 => "0001110100000000000100",
			7920 => "1111111111101111010101",
			7921 => "0000000111101111010101",
			7922 => "0010011101101000000100",
			7923 => "0000000111101111010101",
			7924 => "0000000111101111010101",
			7925 => "0011100101101111001100",
			7926 => "0011110101110101110000",
			7927 => "0000110110000101000000",
			7928 => "0010010111100100100000",
			7929 => "0000011100110100010000",
			7930 => "0010010110101000001000",
			7931 => "0000000011111100000100",
			7932 => "0000000111111010101011",
			7933 => "0000000111111010101011",
			7934 => "0001111011000100000100",
			7935 => "0000000111111010101011",
			7936 => "0000001111111010101011",
			7937 => "0000110011011100001000",
			7938 => "0000101101000100000100",
			7939 => "1111111111111010101011",
			7940 => "0000000111111010101011",
			7941 => "0001110000101000000100",
			7942 => "0000000111111010101011",
			7943 => "1111111111111010101011",
			7944 => "0011110100000100010000",
			7945 => "0011000000101000001000",
			7946 => "0011111010011100000100",
			7947 => "0000001111111010101011",
			7948 => "0000000111111010101011",
			7949 => "0001111100001000000100",
			7950 => "1111111111111010101011",
			7951 => "0000000111111010101011",
			7952 => "0011110100010000001000",
			7953 => "0000101100100100000100",
			7954 => "0000001111111010101011",
			7955 => "0000000111111010101011",
			7956 => "0000100101110000000100",
			7957 => "0000010111111010101011",
			7958 => "0000001111111010101011",
			7959 => "0011010001111100100000",
			7960 => "0011101000111100010000",
			7961 => "0000011100110100001000",
			7962 => "0000100010011100000100",
			7963 => "0000000111111010101011",
			7964 => "1111111111111010101011",
			7965 => "0011110101100100000100",
			7966 => "1111111111111010101011",
			7967 => "0000000111111010101011",
			7968 => "0011000000101000001000",
			7969 => "0000000010111100000100",
			7970 => "0000000111111010101011",
			7971 => "1111111111111010101011",
			7972 => "0011100011011100000100",
			7973 => "1111111111111010101011",
			7974 => "0000000111111010101011",
			7975 => "0001001101001000001100",
			7976 => "0001001110100100001000",
			7977 => "0001011010111100000100",
			7978 => "0000000111111010101011",
			7979 => "1111111111111010101011",
			7980 => "0000001111111010101011",
			7981 => "0000000111111010101011",
			7982 => "0000000000110000111000",
			7983 => "0011011100101100011100",
			7984 => "0001110100010100001100",
			7985 => "0001011100110000001000",
			7986 => "0011001110111100000100",
			7987 => "1111111111111010101011",
			7988 => "0000001111111010101011",
			7989 => "1111111111111010101011",
			7990 => "0001001000001000001000",
			7991 => "0001101101111100000100",
			7992 => "0000001111111010101011",
			7993 => "0000010111111010101011",
			7994 => "0001000011001100000100",
			7995 => "0000000111111010101011",
			7996 => "0000001111111010101011",
			7997 => "0010111100001000001100",
			7998 => "0000111101111000001000",
			7999 => "0011011110001100000100",
			8000 => "1111111111111010101011",
			8001 => "0000000111111010101011",
			8002 => "1111111111111010101011",
			8003 => "0000100010011100001000",
			8004 => "0010011101101000000100",
			8005 => "1111111111111010101011",
			8006 => "0000000111111010101011",
			8007 => "0001111000111000000100",
			8008 => "0000000111111010101011",
			8009 => "0000001111111010101011",
			8010 => "0010110101101100011100",
			8011 => "0010010111100100001100",
			8012 => "0000011100110100001000",
			8013 => "0001000101010100000100",
			8014 => "1111111111111010101011",
			8015 => "0000000111111010101011",
			8016 => "1111111111111010101011",
			8017 => "0001111011000100001000",
			8018 => "0011101101100000000100",
			8019 => "0000001111111010101011",
			8020 => "0000000111111010101011",
			8021 => "0000001010000000000100",
			8022 => "0000000111111010101011",
			8023 => "0000000111111010101011",
			8024 => "0001111101100000000100",
			8025 => "1111110111111010101011",
			8026 => "0000000111111010101011",
			8027 => "0010011101101000111000",
			8028 => "0011110111100000110000",
			8029 => "0001101100011000011100",
			8030 => "0011110010110100010000",
			8031 => "0001000010111000001000",
			8032 => "0000111101111000000100",
			8033 => "0000000111111010101011",
			8034 => "1111111111111010101011",
			8035 => "0011100110000100000100",
			8036 => "0000001111111010101011",
			8037 => "1111111111111010101011",
			8038 => "0011011100101000001000",
			8039 => "0000000011010000000100",
			8040 => "0000001111111010101011",
			8041 => "0000000111111010101011",
			8042 => "0000001111111010101011",
			8043 => "0001001111100000001100",
			8044 => "0000101110010000000100",
			8045 => "0000000111111010101011",
			8046 => "0001010000001100000100",
			8047 => "1111111111111010101011",
			8048 => "1111111111111010101011",
			8049 => "0011100110000100000100",
			8050 => "0000001111111010101011",
			8051 => "0000000111111010101011",
			8052 => "0000111010111000000100",
			8053 => "0000001111111010101011",
			8054 => "0000000111111010101011",
			8055 => "0000001111000100110100",
			8056 => "0000011001111000011100",
			8057 => "0001110100000000001100",
			8058 => "0000100100101000001000",
			8059 => "0001100100110100000100",
			8060 => "1111111111111010101011",
			8061 => "0000001111111010101011",
			8062 => "0000001111111010101011",
			8063 => "0001111000111000001000",
			8064 => "0001001011110000000100",
			8065 => "0000000111111010101011",
			8066 => "0000010111111010101011",
			8067 => "0001011010111100000100",
			8068 => "1111111111111010101011",
			8069 => "0000001111111010101011",
			8070 => "0010011111001100001000",
			8071 => "0000001000101100000100",
			8072 => "0000000111111010101011",
			8073 => "1111111111111010101011",
			8074 => "0010010100110100001000",
			8075 => "0001001000000100000100",
			8076 => "0000000111111010101011",
			8077 => "0000001111111010101011",
			8078 => "0001101001111100000100",
			8079 => "1111111111111010101011",
			8080 => "0000000111111010101011",
			8081 => "0001001100001100010100",
			8082 => "0011001001110000010000",
			8083 => "0001110100000000001000",
			8084 => "0011000100000000000100",
			8085 => "0000000111111010101011",
			8086 => "0000001111111010101011",
			8087 => "0011001000111100000100",
			8088 => "1111111111111010101011",
			8089 => "0000000111111010101011",
			8090 => "0000001111111010101011",
			8091 => "0010011011101000010000",
			8092 => "0000010010001100001000",
			8093 => "0001010001111100000100",
			8094 => "0000000111111010101011",
			8095 => "0000001111111010101011",
			8096 => "0011000000101000000100",
			8097 => "0000000111111010101011",
			8098 => "0000000111111010101011",
			8099 => "0000111000000000001000",
			8100 => "0001001111100000000100",
			8101 => "0000001111111010101011",
			8102 => "1111111111111010101011",
			8103 => "0001001000001000000100",
			8104 => "0000000111111010101011",
			8105 => "0000000111111010101011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2753, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5446, initial_addr_3'length));
	end generate gen_rom_7;

	gen_rom_8: if SELECT_ROM = 8 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0001011111010100000100",
			3 => "0000000000000000010101",
			4 => "1111111000000000010101",
			5 => "0001000101010100000100",
			6 => "0000000000000000101001",
			7 => "0001000001100100000100",
			8 => "0000000000000000101001",
			9 => "0000000000000000101001",
			10 => "0001000011010100000100",
			11 => "0000000000000000111101",
			12 => "0001000001100100000100",
			13 => "0000000000000000111101",
			14 => "0000000000000000111101",
			15 => "0010000110001000001000",
			16 => "0010000001010100000100",
			17 => "0000000000000001010001",
			18 => "0000000000000001010001",
			19 => "0000000000000001010001",
			20 => "0010110010011100001000",
			21 => "0010011001111100000100",
			22 => "0000000000000001100101",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0001110001001000001100",
			26 => "0001000100001100000100",
			27 => "0000000000000010000001",
			28 => "0001000001100100000100",
			29 => "0000000000000010000001",
			30 => "0000000000000010000001",
			31 => "0000000000000010000001",
			32 => "0001110001001000001100",
			33 => "0001000000010100000100",
			34 => "0000000000000010011101",
			35 => "0001000001100100000100",
			36 => "0000000000000010011101",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0010100110011000001100",
			40 => "0010101001000100000100",
			41 => "0000000000000011000001",
			42 => "0001101111000000000100",
			43 => "0000000000000011000001",
			44 => "0000000000000011000001",
			45 => "0010100110011100000100",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0000011100011000001100",
			49 => "0010100110011100001000",
			50 => "0010101000010100000100",
			51 => "0000000000000011100101",
			52 => "0000000000000011100101",
			53 => "0000000000000011100101",
			54 => "0010101010110000000100",
			55 => "0000000000000011100101",
			56 => "0000000000000011100101",
			57 => "0011001011011100001100",
			58 => "0010011001111100000100",
			59 => "0000000000000100001001",
			60 => "0010011000010100000100",
			61 => "0000000000000100001001",
			62 => "0000000000000100001001",
			63 => "0011001011011100000100",
			64 => "0000000000000100001001",
			65 => "0000000000000100001001",
			66 => "0010100110011000001100",
			67 => "0000000010101000000100",
			68 => "0000000000000100110101",
			69 => "0001101111000000000100",
			70 => "0000000000000100110101",
			71 => "0000000000000100110101",
			72 => "0001101000010000000100",
			73 => "0000000000000100110101",
			74 => "0000001000110000000100",
			75 => "0000000000000100110101",
			76 => "0000000000000100110101",
			77 => "0010001011010100001100",
			78 => "0001000011110000000100",
			79 => "0000000000000101100001",
			80 => "0001001111100000000100",
			81 => "0000000000000101100001",
			82 => "0000000000000101100001",
			83 => "0011100011010100001000",
			84 => "0001000000101100000100",
			85 => "0000000000000101100001",
			86 => "0000000000000101100001",
			87 => "0000000000000101100001",
			88 => "0001110001001000010000",
			89 => "0010011001111100000100",
			90 => "0000000000000110000101",
			91 => "0001000011110000000100",
			92 => "0000000000000110000101",
			93 => "0011001000000000000100",
			94 => "0000000000000110000101",
			95 => "0000000000000110000101",
			96 => "0000000000000110000101",
			97 => "0001010000010000010000",
			98 => "0001110001011000000100",
			99 => "0000000000000110101001",
			100 => "0001011110010000000100",
			101 => "0000000000000110101001",
			102 => "0010110001001000000100",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0011111110100100000100",
			107 => "0000000000000111001101",
			108 => "0000011111000000001100",
			109 => "0001100100111100000100",
			110 => "0000000000000111001101",
			111 => "0000110011101100000100",
			112 => "0000000000000111001101",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0011001011011100010000",
			116 => "0010011001111100000100",
			117 => "0000000000000111111001",
			118 => "0011001001110100000100",
			119 => "0000000000000111111001",
			120 => "0010011000010100000100",
			121 => "0000000000000111111001",
			122 => "0000000000000111111001",
			123 => "0011001011011100000100",
			124 => "0000000000000111111001",
			125 => "0000000000000111111001",
			126 => "0001110001001000010100",
			127 => "0001000000010100001000",
			128 => "0000011101011000000100",
			129 => "0000000000001000100101",
			130 => "0000000000001000100101",
			131 => "0010011001111100000100",
			132 => "0000000000001000100101",
			133 => "0011001001110100000100",
			134 => "0000000000001000100101",
			135 => "0000000000001000100101",
			136 => "0000000000001000100101",
			137 => "0001000000010100001100",
			138 => "0001001110100100000100",
			139 => "0000000000001001011001",
			140 => "0011111010110100000100",
			141 => "0000000000001001011001",
			142 => "0000000000001001011001",
			143 => "0001000001100100001100",
			144 => "0000101101101100000100",
			145 => "0000000000001001011001",
			146 => "0000101110100100000100",
			147 => "0000000000001001011001",
			148 => "0000000000001001011001",
			149 => "0000000000001001011001",
			150 => "0010110110100000010100",
			151 => "0001011001010100000100",
			152 => "0000000000001010001101",
			153 => "0010100101000100001100",
			154 => "0010101000010100000100",
			155 => "0000000000001010001101",
			156 => "0000110010111000000100",
			157 => "0000000000001010001101",
			158 => "0000000000001010001101",
			159 => "0000000000001010001101",
			160 => "0011011111010100000100",
			161 => "0000000000001010001101",
			162 => "0000000000001010001101",
			163 => "0010001111001000010100",
			164 => "0000100110111000000100",
			165 => "0000000000001011000001",
			166 => "0011001000000000000100",
			167 => "0000000000001011000001",
			168 => "0011001011011100001000",
			169 => "0000000001110100000100",
			170 => "0000000000001011000001",
			171 => "0000000000001011000001",
			172 => "0000000000001011000001",
			173 => "0000101110000000000100",
			174 => "0000000000001011000001",
			175 => "0000000000001011000001",
			176 => "0001110001001000010100",
			177 => "0011000100011000000100",
			178 => "0000000000001011101101",
			179 => "0001100100101100001100",
			180 => "0000101101101100000100",
			181 => "0000000000001011101101",
			182 => "0001101111000000000100",
			183 => "0000000000001011101101",
			184 => "0000000000001011101101",
			185 => "0000000000001011101101",
			186 => "0000000000001011101101",
			187 => "0001000000010100001100",
			188 => "0001100100111100000100",
			189 => "0000000000001100101001",
			190 => "0011111010110100000100",
			191 => "0000000000001100101001",
			192 => "0000000000001100101001",
			193 => "0001101001111100010000",
			194 => "0001011001010100000100",
			195 => "0000000000001100101001",
			196 => "0011011100010000001000",
			197 => "0001000001100100000100",
			198 => "0000000000001100101001",
			199 => "0000000000001100101001",
			200 => "0000000000001100101001",
			201 => "0000000000001100101001",
			202 => "0001111011110100010100",
			203 => "0010011001111100000100",
			204 => "0000000000001101100101",
			205 => "0000100110111000000100",
			206 => "0000000000001101100101",
			207 => "0010000111000100001000",
			208 => "0011001001110100000100",
			209 => "0000000000001101100101",
			210 => "0000000000001101100101",
			211 => "0000000000001101100101",
			212 => "0001101000010000000100",
			213 => "0000000000001101100101",
			214 => "0010111101000100000100",
			215 => "0000000000001101100101",
			216 => "0000000000001101100101",
			217 => "0001111000011000010100",
			218 => "0001111011000000000100",
			219 => "0000000000001110101001",
			220 => "0001001000001000000100",
			221 => "0000000000001110101001",
			222 => "0010100001010100001000",
			223 => "0011111000110100000100",
			224 => "0000001000001110101001",
			225 => "0000000000001110101001",
			226 => "0000000000001110101001",
			227 => "0010000110001000000100",
			228 => "0000000000001110101001",
			229 => "0011100011010100001000",
			230 => "0001101000010000000100",
			231 => "0000000000001110101001",
			232 => "0000000000001110101001",
			233 => "0000000000001110101001",
			234 => "0000101011110000010000",
			235 => "0000101101101100000100",
			236 => "0000000000001111101101",
			237 => "0001101000010000001000",
			238 => "0001101111000000000100",
			239 => "0000000000001111101101",
			240 => "0000000000001111101101",
			241 => "0000000000001111101101",
			242 => "0010000001010100000100",
			243 => "0000000000001111101101",
			244 => "0001100100111100000100",
			245 => "0000000000001111101101",
			246 => "0001001110100100000100",
			247 => "0000000000001111101101",
			248 => "0010101000010100000100",
			249 => "0000000000001111101101",
			250 => "0000000000001111101101",
			251 => "0010011010100000001100",
			252 => "0011111110100100001000",
			253 => "0001000111011100000100",
			254 => "0000000000010000111001",
			255 => "0000000000010000111001",
			256 => "0000000000010000111001",
			257 => "0011111100001100001100",
			258 => "0011000100000100001000",
			259 => "0001110111010000000100",
			260 => "0000000000010000111001",
			261 => "0000000000010000111001",
			262 => "0000000000010000111001",
			263 => "0001000000010100001100",
			264 => "0010011000100100001000",
			265 => "0001000011110000000100",
			266 => "0000000000010000111001",
			267 => "0000000000010000111001",
			268 => "0000000000010000111001",
			269 => "0000000000010000111001",
			270 => "0010100110011000010100",
			271 => "0010101000010100000100",
			272 => "0000000000010010001101",
			273 => "0000100110111000000100",
			274 => "0000000000010010001101",
			275 => "0001011100010000001000",
			276 => "0011001001110100000100",
			277 => "0000000000010010001101",
			278 => "0000001000010010001101",
			279 => "0000000000010010001101",
			280 => "0001001011001000001100",
			281 => "0010011000100100001000",
			282 => "0010001100000100000100",
			283 => "0000000000010010001101",
			284 => "0000000000010010001101",
			285 => "0000000000010010001101",
			286 => "0010100101000100001000",
			287 => "0010101100011100000100",
			288 => "0000000000010010001101",
			289 => "0000000000010010001101",
			290 => "0000000000010010001101",
			291 => "0001100101010000011000",
			292 => "0011011010000100010100",
			293 => "0001101111000000000100",
			294 => "0000000000010011001001",
			295 => "0011011110101100000100",
			296 => "0000000000010011001001",
			297 => "0010101000100100000100",
			298 => "0000000000010011001001",
			299 => "0001101000010000000100",
			300 => "0000000000010011001001",
			301 => "0000000000010011001001",
			302 => "0000000000010011001001",
			303 => "0010001001101000000100",
			304 => "0000000000010011001001",
			305 => "0000000000010011001001",
			306 => "0010000110001000011000",
			307 => "0001001110100100000100",
			308 => "0000000000010100000101",
			309 => "0011001001110100000100",
			310 => "0000000000010100000101",
			311 => "0001111011110100001100",
			312 => "0000011110010100000100",
			313 => "0000000000010100000101",
			314 => "0010000101000100000100",
			315 => "0000000000010100000101",
			316 => "0000000000010100000101",
			317 => "0000000000010100000101",
			318 => "0001001001000000000100",
			319 => "0000000000010100000101",
			320 => "0000000000010100000101",
			321 => "0001000000101100100000",
			322 => "0010010111101100001000",
			323 => "0001000111011100000100",
			324 => "0000000000010101011001",
			325 => "0000000000010101011001",
			326 => "0001101000010000001000",
			327 => "0010011010100100000100",
			328 => "0000000000010101011001",
			329 => "0000000000010101011001",
			330 => "0001000000010100001000",
			331 => "0010010011101000000100",
			332 => "0000000000010101011001",
			333 => "0000000000010101011001",
			334 => "0010011000010100000100",
			335 => "0000000000010101011001",
			336 => "0000000000010101011001",
			337 => "0010100101000100001000",
			338 => "0011000001111100000100",
			339 => "0000000000010101011001",
			340 => "0000001000010101011001",
			341 => "0000000000010101011001",
			342 => "0001000100001100011000",
			343 => "0000011101011000010100",
			344 => "0010000101000100000100",
			345 => "0000000000010110100101",
			346 => "0001011110110100001100",
			347 => "0000000001110100000100",
			348 => "0000000000010110100101",
			349 => "0010111101000100000100",
			350 => "0000000000010110100101",
			351 => "0000000000010110100101",
			352 => "0000000000010110100101",
			353 => "0000000000010110100101",
			354 => "0010000111000100001100",
			355 => "0000011011111100000100",
			356 => "0000000000010110100101",
			357 => "0000000010111100000100",
			358 => "0000000000010110100101",
			359 => "0000000000010110100101",
			360 => "0000000000010110100101",
			361 => "0001000000010100011000",
			362 => "0010110000110100010100",
			363 => "0001111011011100010000",
			364 => "0011001111011100001100",
			365 => "0000011011001100001000",
			366 => "0010000101000100000100",
			367 => "0000000000010111110001",
			368 => "0000000000010111110001",
			369 => "0000000000010111110001",
			370 => "0000000000010111110001",
			371 => "0000000000010111110001",
			372 => "0000000000010111110001",
			373 => "0010001111001000001100",
			374 => "0000011011111100000100",
			375 => "0000000000010111110001",
			376 => "0001110111110000000100",
			377 => "0000000000010111110001",
			378 => "0000000000010111110001",
			379 => "0000000000010111110001",
			380 => "0001011001100000011100",
			381 => "0011001001110100001000",
			382 => "0001000000101100000100",
			383 => "0000000000011001000101",
			384 => "0000000000011001000101",
			385 => "0010000111000100010000",
			386 => "0011101000011100001100",
			387 => "0001001110100100000100",
			388 => "0000000000011001000101",
			389 => "0010011001111100000100",
			390 => "0000000000011001000101",
			391 => "0000000000011001000101",
			392 => "0000000000011001000101",
			393 => "0000000000011001000101",
			394 => "0001101000010000000100",
			395 => "0000000000011001000101",
			396 => "0010110110100000000100",
			397 => "0000000000011001000101",
			398 => "0001110100010000000100",
			399 => "0000000000011001000101",
			400 => "0000000000011001000101",
			401 => "0001011110000100010000",
			402 => "0000011001011000000100",
			403 => "0000000000011010100001",
			404 => "0001001111100000000100",
			405 => "0000000000011010100001",
			406 => "0011001010111100000100",
			407 => "0000000000011010100001",
			408 => "0000001000011010100001",
			409 => "0000011010011000010000",
			410 => "0001111111011100000100",
			411 => "0000000000011010100001",
			412 => "0010101000010100000100",
			413 => "0000000000011010100001",
			414 => "0010000001010100000100",
			415 => "0000000000011010100001",
			416 => "0000000000011010100001",
			417 => "0010000001110100001100",
			418 => "0001110111010000000100",
			419 => "0000000000011010100001",
			420 => "0000001010101100000100",
			421 => "0000000000011010100001",
			422 => "0000000000011010100001",
			423 => "0000000000011010100001",
			424 => "0010011010100000001100",
			425 => "0011111110100100001000",
			426 => "0001000111011100000100",
			427 => "0000000000011011111101",
			428 => "0000000000011011111101",
			429 => "0000000000011011111101",
			430 => "0011101000011100010100",
			431 => "0011000100000100010000",
			432 => "0001101001111100001100",
			433 => "0001011001010000000100",
			434 => "0000000000011011111101",
			435 => "0010110100010000000100",
			436 => "0000000000011011111101",
			437 => "0000000000011011111101",
			438 => "0000000000011011111101",
			439 => "0000000000011011111101",
			440 => "0010011000100100001100",
			441 => "0011001001110100000100",
			442 => "0000000000011011111101",
			443 => "0001110111110000000100",
			444 => "0000000000011011111101",
			445 => "0000000000011011111101",
			446 => "0000000000011011111101",
			447 => "0000101011110000010100",
			448 => "0000101101101100000100",
			449 => "0000000000011101100001",
			450 => "0011001010111000000100",
			451 => "0000000000011101100001",
			452 => "0010011011001100000100",
			453 => "0000000000011101100001",
			454 => "0011110010010100000100",
			455 => "0000001000011101100001",
			456 => "0000000000011101100001",
			457 => "0011010110111100001100",
			458 => "0000011100011000000100",
			459 => "0000000000011101100001",
			460 => "0010001111001000000100",
			461 => "0000000000011101100001",
			462 => "0000000000011101100001",
			463 => "0010011000100100010000",
			464 => "0011001111011100000100",
			465 => "0000000000011101100001",
			466 => "0000111110100100000100",
			467 => "0000000000011101100001",
			468 => "0000011010011000000100",
			469 => "0000000000011101100001",
			470 => "0000000000011101100001",
			471 => "0000000000011101100001",
			472 => "0011011010000100100000",
			473 => "0011001001110100001000",
			474 => "0001000000101100000100",
			475 => "0000000000011110101101",
			476 => "0000000000011110101101",
			477 => "0001001110100100000100",
			478 => "0000000000011110101101",
			479 => "0010000111000100010000",
			480 => "0011101000011100001100",
			481 => "0011000001011000001000",
			482 => "0000011110010100000100",
			483 => "0000000000011110101101",
			484 => "0000000000011110101101",
			485 => "0000000000011110101101",
			486 => "0000000000011110101101",
			487 => "0000000000011110101101",
			488 => "0000011101011000000100",
			489 => "0000000000011110101101",
			490 => "0000000000011110101101",
			491 => "0011010110111100011100",
			492 => "0001111011000000000100",
			493 => "0000000000011111111001",
			494 => "0001100101010000010100",
			495 => "0010010011101000010000",
			496 => "0001101001100100000100",
			497 => "0000000000011111111001",
			498 => "0010011011001100000100",
			499 => "0000000000011111111001",
			500 => "0000101100111000000100",
			501 => "0000000000011111111001",
			502 => "0000000000011111111001",
			503 => "0000000000011111111001",
			504 => "0000000000011111111001",
			505 => "0000101000000100000100",
			506 => "0000000000011111111001",
			507 => "0001101000010000000100",
			508 => "0000000000011111111001",
			509 => "0000000000011111111001",
			510 => "0001000011011000100100",
			511 => "0010000110001000011000",
			512 => "0010010111101100000100",
			513 => "0000000000100001010101",
			514 => "0010110110100000010000",
			515 => "0011101000011100001100",
			516 => "0000110001011100000100",
			517 => "0000000000100001010101",
			518 => "0010110100010000000100",
			519 => "0000000000100001010101",
			520 => "0000000000100001010101",
			521 => "0000000000100001010101",
			522 => "0000000000100001010101",
			523 => "0001001001000000001000",
			524 => "0000111110111000000100",
			525 => "0000000000100001010101",
			526 => "0000000000100001010101",
			527 => "0000000000100001010101",
			528 => "0010001010101100001000",
			529 => "0001101000010000000100",
			530 => "0000000000100001010101",
			531 => "0000001000100001010101",
			532 => "0000000000100001010101",
			533 => "0011100110111000011100",
			534 => "0011001001110100000100",
			535 => "0000000000100010101001",
			536 => "0010000111000100010100",
			537 => "0000111011111000000100",
			538 => "0000000000100010101001",
			539 => "0011000111010000001100",
			540 => "0000100010010100000100",
			541 => "0000000000100010101001",
			542 => "0011011100010000000100",
			543 => "0000000000100010101001",
			544 => "0000000000100010101001",
			545 => "0000000000100010101001",
			546 => "0000000000100010101001",
			547 => "0001000110001100000100",
			548 => "0000000000100010101001",
			549 => "0010101000010100000100",
			550 => "0000000000100010101001",
			551 => "0011111000110100000100",
			552 => "0000000000100010101001",
			553 => "0000000000100010101001",
			554 => "0001000011011000101000",
			555 => "0000011010011000010100",
			556 => "0000110101000000010000",
			557 => "0010000101000100000100",
			558 => "0000000000100100001101",
			559 => "0001000011101100001000",
			560 => "0010010011101000000100",
			561 => "0000000000100100001101",
			562 => "0000000000100100001101",
			563 => "0000000000100100001101",
			564 => "0000000000100100001101",
			565 => "0011011010000100010000",
			566 => "0011111001001100001100",
			567 => "0001001110100100000100",
			568 => "0000000000100100001101",
			569 => "0001010101110000000100",
			570 => "0000000000100100001101",
			571 => "0000000000100100001101",
			572 => "0000000000100100001101",
			573 => "0000000000100100001101",
			574 => "0010100101000100001000",
			575 => "0000011001011000000100",
			576 => "0000000000100100001101",
			577 => "0000001000100100001101",
			578 => "0000000000100100001101",
			579 => "0000010100110100010100",
			580 => "0001000111011100000100",
			581 => "0000000000100110000001",
			582 => "0010000001110100001100",
			583 => "0000000000111000000100",
			584 => "0000000000100110000001",
			585 => "0000011001011000000100",
			586 => "0000000000100110000001",
			587 => "0000000000100110000001",
			588 => "0000000000100110000001",
			589 => "0000110110001100001100",
			590 => "0011000100000100001000",
			591 => "0001110111010000000100",
			592 => "0000000000100110000001",
			593 => "0000000000100110000001",
			594 => "0000000000100110000001",
			595 => "0011000111010000010000",
			596 => "0011110110001100000100",
			597 => "0000000000100110000001",
			598 => "0010101001000100000100",
			599 => "0000000000100110000001",
			600 => "0001110100010000000100",
			601 => "0000000000100110000001",
			602 => "0000000000100110000001",
			603 => "0000010100111100001000",
			604 => "0011000100000100000100",
			605 => "0000000000100110000001",
			606 => "0000000000100110000001",
			607 => "0000000000100110000001",
			608 => "0001000011011000101100",
			609 => "0000011010011000011000",
			610 => "0010111110101100010000",
			611 => "0010000101000100000100",
			612 => "0000000000100111101101",
			613 => "0001111011011100001000",
			614 => "0010001100000100000100",
			615 => "0000000000100111101101",
			616 => "0000000000100111101101",
			617 => "0000000000100111101101",
			618 => "0010001100000100000100",
			619 => "0000000000100111101101",
			620 => "0000000000100111101101",
			621 => "0011011010000100010000",
			622 => "0011101000001000001100",
			623 => "0001011110110100001000",
			624 => "0001110111010000000100",
			625 => "0000000000100111101101",
			626 => "0000000000100111101101",
			627 => "0000000000100111101101",
			628 => "0000000000100111101101",
			629 => "0000000000100111101101",
			630 => "0010100101000100001000",
			631 => "0000011001011000000100",
			632 => "0000000000100111101101",
			633 => "0000001000100111101101",
			634 => "0000000000100111101101",
			635 => "0010001100000100011100",
			636 => "0010111110101100010000",
			637 => "0000011010011000001100",
			638 => "0000001010101100000100",
			639 => "0000000000101001100001",
			640 => "0000001000110000000100",
			641 => "0000000000101001100001",
			642 => "0000000000101001100001",
			643 => "0000000000101001100001",
			644 => "0000011101011000001000",
			645 => "0010011010100100000100",
			646 => "0000000000101001100001",
			647 => "0000000000101001100001",
			648 => "0000000000101001100001",
			649 => "0001000000010100001000",
			650 => "0010011000100100000100",
			651 => "0000000000101001100001",
			652 => "0000000000101001100001",
			653 => "0000000111111000010100",
			654 => "0001100100101100010000",
			655 => "0000000010011000000100",
			656 => "0000000000101001100001",
			657 => "0001100100111100000100",
			658 => "0000000000101001100001",
			659 => "0001101001111100000100",
			660 => "0000000000101001100001",
			661 => "0000000000101001100001",
			662 => "0000000000101001100001",
			663 => "0000000000101001100001",
			664 => "0000001011000100101000",
			665 => "0001111011011100011000",
			666 => "0000011010011000010100",
			667 => "0010100001010000010000",
			668 => "0010000101000100000100",
			669 => "0000000000101010111101",
			670 => "0010111110101100001000",
			671 => "0000000001110100000100",
			672 => "0000000000101010111101",
			673 => "0000000000101010111101",
			674 => "0000000000101010111101",
			675 => "0000000000101010111101",
			676 => "0000000000101010111101",
			677 => "0001111011110100001100",
			678 => "0010000111000100001000",
			679 => "0001101111000000000100",
			680 => "0000000000101010111101",
			681 => "0000000000101010111101",
			682 => "0000000000101010111101",
			683 => "0000000000101010111101",
			684 => "0000000000101000000100",
			685 => "0000000000101010111101",
			686 => "0000000000101010111101",
			687 => "0000010100110100010100",
			688 => "0001000111011100000100",
			689 => "0000000000101100111001",
			690 => "0010000001110100001100",
			691 => "0000000000111000000100",
			692 => "0000000000101100111001",
			693 => "0000011001011000000100",
			694 => "0000000000101100111001",
			695 => "0000000000101100111001",
			696 => "0000000000101100111001",
			697 => "0011101000011100010100",
			698 => "0011000100000100010000",
			699 => "0001110111010000000100",
			700 => "0000000000101100111001",
			701 => "0010110110100000001000",
			702 => "0011001001110100000100",
			703 => "0000000000101100111001",
			704 => "0000000000101100111001",
			705 => "0000000000101100111001",
			706 => "0000000000101100111001",
			707 => "0011000100000100010000",
			708 => "0010010111110100001100",
			709 => "0010101001000100000100",
			710 => "0000000000101100111001",
			711 => "0000011011001100000100",
			712 => "0000000000101100111001",
			713 => "0000000000101100111001",
			714 => "0000000000101100111001",
			715 => "0000010100111100000100",
			716 => "0000000000101100111001",
			717 => "0000000000101100111001",
			718 => "0001000000101100110000",
			719 => "0001100101010000100100",
			720 => "0000101000110100010100",
			721 => "0001000111011100010000",
			722 => "0010000001010100000100",
			723 => "0000000000101110101101",
			724 => "0000011101011000001000",
			725 => "0011111000011100000100",
			726 => "0000000000101110101101",
			727 => "0000000000101110101101",
			728 => "0000000000101110101101",
			729 => "0000000000101110101101",
			730 => "0011011010000100001100",
			731 => "0000010111101000000100",
			732 => "0000000000101110101101",
			733 => "0011110011001100000100",
			734 => "0000000000101110101101",
			735 => "0000000000101110101101",
			736 => "0000000000101110101101",
			737 => "0010010111110100001000",
			738 => "0001000011101100000100",
			739 => "0000000000101110101101",
			740 => "0000000000101110101101",
			741 => "0000000000101110101101",
			742 => "0010100101000100001000",
			743 => "0000011001011000000100",
			744 => "0000000000101110101101",
			745 => "0000001000101110101101",
			746 => "0000000000101110101101",
			747 => "0011001001110100010000",
			748 => "0001010111111100001100",
			749 => "0010100110011100000100",
			750 => "1111111000110000111001",
			751 => "0010100110011100000100",
			752 => "0000000000110000111001",
			753 => "0000000000110000111001",
			754 => "0000000000110000111001",
			755 => "0010011010100100010100",
			756 => "0000101100001100001100",
			757 => "0000111000000100001000",
			758 => "0001100100111100000100",
			759 => "0000000000110000111001",
			760 => "0000000000110000111001",
			761 => "0000000000110000111001",
			762 => "0011011110110100000100",
			763 => "0000000000110000111001",
			764 => "0000000000110000111001",
			765 => "0011010110111100001100",
			766 => "0000110010111000001000",
			767 => "0000011100011000000100",
			768 => "0000000000110000111001",
			769 => "0000001000110000111001",
			770 => "0000000000110000111001",
			771 => "0001110100010000001100",
			772 => "0000111100001100000100",
			773 => "0000000000110000111001",
			774 => "0010000001010100000100",
			775 => "0000000000110000111001",
			776 => "0000000000110000111001",
			777 => "0001100100101100001000",
			778 => "0011101110000000000100",
			779 => "0000000000110000111001",
			780 => "0000001000110000111001",
			781 => "0000000000110000111001",
			782 => "0000100011000000001100",
			783 => "0000000001110100000100",
			784 => "0000000000110010110101",
			785 => "0001010111111100000100",
			786 => "0000000000110010110101",
			787 => "0000000000110010110101",
			788 => "0011100110111000011000",
			789 => "0011000001011000010100",
			790 => "0000000111111000010000",
			791 => "0000100010010100000100",
			792 => "0000000000110010110101",
			793 => "0000010101011100000100",
			794 => "0000000000110010110101",
			795 => "0011001010111000000100",
			796 => "0000000000110010110101",
			797 => "0000000000110010110101",
			798 => "0000000000110010110101",
			799 => "0000000000110010110101",
			800 => "0000011101011000010000",
			801 => "0010010011101000000100",
			802 => "0000000000110010110101",
			803 => "0011111000011100000100",
			804 => "0000000000110010110101",
			805 => "0000000111000000000100",
			806 => "0000000000110010110101",
			807 => "0000000000110010110101",
			808 => "0000000011010000001000",
			809 => "0000001010101100000100",
			810 => "0000000000110010110101",
			811 => "0000000000110010110101",
			812 => "0000000000110010110101",
			813 => "0000010101011100000100",
			814 => "1111111000110100100001",
			815 => "0001100101010000100100",
			816 => "0010010011101000011000",
			817 => "0010011010100100010000",
			818 => "0000000010011000001100",
			819 => "0001100100111100000100",
			820 => "0000000000110100100001",
			821 => "0000111000000100000100",
			822 => "0000000000110100100001",
			823 => "0000000000110100100001",
			824 => "0000000000110100100001",
			825 => "0001010010011100000100",
			826 => "0000000000110100100001",
			827 => "0000001000110100100001",
			828 => "0010101000010100001000",
			829 => "0000110101000000000100",
			830 => "0000000000110100100001",
			831 => "1111111000110100100001",
			832 => "0000000000110100100001",
			833 => "0001111111011100000100",
			834 => "0000000000110100100001",
			835 => "0000011101011000000100",
			836 => "0000000000110100100001",
			837 => "0010000111000100000100",
			838 => "0000000000110100100001",
			839 => "0000000000110100100001",
			840 => "0010011010100100100100",
			841 => "0010011010100100011100",
			842 => "0010010100111100000100",
			843 => "1111111000110110111101",
			844 => "0001111000011000001000",
			845 => "0010011000010000000100",
			846 => "0000000000110110111101",
			847 => "1111111000110110111101",
			848 => "0011101111101000001100",
			849 => "0001101000010000000100",
			850 => "1111111000110110111101",
			851 => "0001100101010000000100",
			852 => "0000010000110110111101",
			853 => "0000000000110110111101",
			854 => "1111111000110110111101",
			855 => "0001111111011100000100",
			856 => "1111111000110110111101",
			857 => "0000001000110110111101",
			858 => "0001110111010000010000",
			859 => "0001010111111100001100",
			860 => "0011001001110100000100",
			861 => "1111111000110110111101",
			862 => "0010110101110100000100",
			863 => "0000000000110110111101",
			864 => "1111111000110110111101",
			865 => "0000001000110110111101",
			866 => "0010000111000100011000",
			867 => "0010101010110000010000",
			868 => "0001110000011100001000",
			869 => "0000001000101100000100",
			870 => "0000001000110110111101",
			871 => "0000001000110110111101",
			872 => "0000000010011000000100",
			873 => "0000001000110110111101",
			874 => "0000010000110110111101",
			875 => "0000000011111100000100",
			876 => "0000000000110110111101",
			877 => "0000001000110110111101",
			878 => "1111111000110110111101",
			879 => "0010010100111100000100",
			880 => "1111111000111000110001",
			881 => "0001000011010100100100",
			882 => "0001100100111100001100",
			883 => "0010011010100100000100",
			884 => "0000000000111000110001",
			885 => "0010110100010000000100",
			886 => "0000000000111000110001",
			887 => "0000000000111000110001",
			888 => "0000011101011000010000",
			889 => "0001110111110000001100",
			890 => "0001000000010100001000",
			891 => "0010000101000100000100",
			892 => "0000000000111000110001",
			893 => "0000000000111000110001",
			894 => "0000000000111000110001",
			895 => "0000000000111000110001",
			896 => "0010001001101000000100",
			897 => "0000000000111000110001",
			898 => "0000000000111000110001",
			899 => "0010100101000100010000",
			900 => "0011011001100000000100",
			901 => "0000001000111000110001",
			902 => "0011011010000100000100",
			903 => "0000000000111000110001",
			904 => "0000011010011000000100",
			905 => "0000000000111000110001",
			906 => "0000000000111000110001",
			907 => "0000000000111000110001",
			908 => "0000011100011000101100",
			909 => "0010011010100000011000",
			910 => "0000011011111100000100",
			911 => "1111111000111011000101",
			912 => "0001110001101000000100",
			913 => "1111111000111011000101",
			914 => "0011011001010000000100",
			915 => "0000001000111011000101",
			916 => "0011101011101100001000",
			917 => "0011001001110100000100",
			918 => "1111111000111011000101",
			919 => "0000000000111011000101",
			920 => "1111111000111011000101",
			921 => "0001111111011100000100",
			922 => "1111111000111011000101",
			923 => "0011100010010100001000",
			924 => "0000010100110100000100",
			925 => "0000001000111011000101",
			926 => "0000001000111011000101",
			927 => "0001100101010000000100",
			928 => "0000000000111011000101",
			929 => "1111111000111011000101",
			930 => "0011010011001000000100",
			931 => "1111111000111011000101",
			932 => "0010000110001000010100",
			933 => "0001110111010000000100",
			934 => "0000000000111011000101",
			935 => "0011000101100100001100",
			936 => "0010111110101000001000",
			937 => "0010110000110100000100",
			938 => "0000001000111011000101",
			939 => "0000001000111011000101",
			940 => "0000000000111011000101",
			941 => "0000000000111011000101",
			942 => "0001000111011100000100",
			943 => "1111111000111011000101",
			944 => "0000000000111011000101",
			945 => "0010010100111100000100",
			946 => "1111111000111101001001",
			947 => "0011000001101000011100",
			948 => "0010100001010000001100",
			949 => "0001010111111100001000",
			950 => "0010000101000100000100",
			951 => "0000000000111101001001",
			952 => "0000000000111101001001",
			953 => "0000000000111101001001",
			954 => "0000100011110000001000",
			955 => "0001001111100000000100",
			956 => "0000000000111101001001",
			957 => "0000000000111101001001",
			958 => "0010001011010100000100",
			959 => "0000000000111101001001",
			960 => "0000000000111101001001",
			961 => "0001001100001100001000",
			962 => "0010011010100100000100",
			963 => "0000000000111101001001",
			964 => "0000001000111101001001",
			965 => "0000101000110100001100",
			966 => "0001111011011100000100",
			967 => "0000000000111101001001",
			968 => "0000011101011000000100",
			969 => "0000000000111101001001",
			970 => "0000000000111101001001",
			971 => "0010000111000100001100",
			972 => "0000001010101100000100",
			973 => "0000000000111101001001",
			974 => "0000010100110100000100",
			975 => "0000000000111101001001",
			976 => "0000000000111101001001",
			977 => "0000000000111101001001",
			978 => "0000011100011000110100",
			979 => "0010011010100100101100",
			980 => "0010011010100100100000",
			981 => "0000010101011100000100",
			982 => "1111111000111111100101",
			983 => "0011001001110100001100",
			984 => "0010011000010000000100",
			985 => "0000000000111111100101",
			986 => "0010011001111100000100",
			987 => "1111111000111111100101",
			988 => "1111111000111111100101",
			989 => "0011101011101100001000",
			990 => "0000101000000100000100",
			991 => "1111111000111111100101",
			992 => "0000010000111111100101",
			993 => "0010011010100000000100",
			994 => "1111111000111111100101",
			995 => "0000000000111111100101",
			996 => "0011000001101000001000",
			997 => "0001011001010000000100",
			998 => "1111111000111111100101",
			999 => "0000000000111111100101",
			1000 => "0000010000111111100101",
			1001 => "0001101000010000000100",
			1002 => "0000011000111111100101",
			1003 => "1111111000111111100101",
			1004 => "0001010111111100001000",
			1005 => "0001110111010000000100",
			1006 => "1111111000111111100101",
			1007 => "0000010000111111100101",
			1008 => "0010001111001000001100",
			1009 => "0010000110001000001000",
			1010 => "0010011010100100000100",
			1011 => "0000011000111111100101",
			1012 => "0000011000111111100101",
			1013 => "0000010000111111100101",
			1014 => "0001110101110100000100",
			1015 => "1111111000111111100101",
			1016 => "0000001000111111100101",
			1017 => "0000100011000000001000",
			1018 => "0011001001110100000100",
			1019 => "0000000001000001111001",
			1020 => "0000000001000001111001",
			1021 => "0001010110010000100100",
			1022 => "0000011100011000011000",
			1023 => "0001001001000000010000",
			1024 => "0011111000001000001100",
			1025 => "0000001010101100000100",
			1026 => "0000000001000001111001",
			1027 => "0011110010010100000100",
			1028 => "0000000001000001111001",
			1029 => "0000000001000001111001",
			1030 => "0000000001000001111001",
			1031 => "0000000111111000000100",
			1032 => "0000000001000001111001",
			1033 => "0000000001000001111001",
			1034 => "0011100011110000001000",
			1035 => "0011001001110100000100",
			1036 => "0000000001000001111001",
			1037 => "0000000001000001111001",
			1038 => "0000000001000001111001",
			1039 => "0011000111010000010100",
			1040 => "0010010011101000000100",
			1041 => "0000000001000001111001",
			1042 => "0000110101000000000100",
			1043 => "0000000001000001111001",
			1044 => "0001110101110100001000",
			1045 => "0011010110111100000100",
			1046 => "0000000001000001111001",
			1047 => "0000000001000001111001",
			1048 => "0000000001000001111001",
			1049 => "0001100100101100001000",
			1050 => "0011101110000000000100",
			1051 => "0000000001000001111001",
			1052 => "0000000001000001111001",
			1053 => "0000000001000001111001",
			1054 => "0010010100101100000100",
			1055 => "1111111001000011101101",
			1056 => "0001000011110000100000",
			1057 => "0001111011011100010100",
			1058 => "0000011010011000010000",
			1059 => "0001100100111100000100",
			1060 => "0000000001000011101101",
			1061 => "0010111110101100001000",
			1062 => "0010101000100100000100",
			1063 => "0000000001000011101101",
			1064 => "1111111001000011101101",
			1065 => "0000000001000011101101",
			1066 => "0000000001000011101101",
			1067 => "0011011111010100001000",
			1068 => "0000000111000000000100",
			1069 => "0000000001000011101101",
			1070 => "0000000001000011101101",
			1071 => "0000000001000011101101",
			1072 => "0001100100101100010100",
			1073 => "0011001011011100010000",
			1074 => "0011001001110100000100",
			1075 => "0000000001000011101101",
			1076 => "0011100110001100001000",
			1077 => "0001111000011000000100",
			1078 => "0000000001000011101101",
			1079 => "0000000001000011101101",
			1080 => "0000000001000011101101",
			1081 => "0000000001000011101101",
			1082 => "0000000001000011101101",
			1083 => "0000100011000000001100",
			1084 => "0010000101000100000100",
			1085 => "0000000001000101110001",
			1086 => "0011000001101000000100",
			1087 => "0000000001000101110001",
			1088 => "0000000001000101110001",
			1089 => "0001100100101100110100",
			1090 => "0000000111000000011000",
			1091 => "0010000001010100001000",
			1092 => "0010011010100100000100",
			1093 => "0000000001000101110001",
			1094 => "0000000001000101110001",
			1095 => "0010010011101000000100",
			1096 => "0000000001000101110001",
			1097 => "0000111110100100000100",
			1098 => "0000000001000101110001",
			1099 => "0010010011101000000100",
			1100 => "0000000001000101110001",
			1101 => "0000000001000101110001",
			1102 => "0010010010101100010100",
			1103 => "0001001001000000001100",
			1104 => "0011111000001000001000",
			1105 => "0011110010010100000100",
			1106 => "0000000001000101110001",
			1107 => "0000000001000101110001",
			1108 => "0000000001000101110001",
			1109 => "0001000000101100000100",
			1110 => "0000000001000101110001",
			1111 => "0000000001000101110001",
			1112 => "0011001000011000000100",
			1113 => "0000000001000101110001",
			1114 => "0000000001000101110001",
			1115 => "0000000001000101110001",
			1116 => "0010010111101100001000",
			1117 => "0001000000100000000100",
			1118 => "1111111001001000010101",
			1119 => "0000000001001000010101",
			1120 => "0011101000011100110100",
			1121 => "0001000110001100100000",
			1122 => "0001101000010000010000",
			1123 => "0001010111111100001000",
			1124 => "0001101111000000000100",
			1125 => "0000000001001000010101",
			1126 => "0000000001001000010101",
			1127 => "0001000110001100000100",
			1128 => "0000001001001000010101",
			1129 => "0000000001001000010101",
			1130 => "0001110100010000001100",
			1131 => "0001001100001100001000",
			1132 => "0011001010001100000100",
			1133 => "0000000001001000010101",
			1134 => "0000000001001000010101",
			1135 => "0000000001001000010101",
			1136 => "0000000001001000010101",
			1137 => "0001100101010000001100",
			1138 => "0010110100010000000100",
			1139 => "0000000001001000010101",
			1140 => "0011000001011000000100",
			1141 => "0000001001001000010101",
			1142 => "0000000001001000010101",
			1143 => "0011000111010000000100",
			1144 => "0000000001001000010101",
			1145 => "0000000001001000010101",
			1146 => "0010010111110100001100",
			1147 => "0001110100010000001000",
			1148 => "0011000111010000000100",
			1149 => "1111111001001000010101",
			1150 => "0000000001001000010101",
			1151 => "0000000001001000010101",
			1152 => "0001100100101100001000",
			1153 => "0011001111011100000100",
			1154 => "0000000001001000010101",
			1155 => "0000000001001000010101",
			1156 => "0000000001001000010101",
			1157 => "0010011010100100011100",
			1158 => "0000101101101100000100",
			1159 => "1111111001001011001001",
			1160 => "0011101111101000010100",
			1161 => "0011000100011000000100",
			1162 => "1111111001001011001001",
			1163 => "0001111001001000000100",
			1164 => "0000010001001011001001",
			1165 => "0010010101010000000100",
			1166 => "1111111001001011001001",
			1167 => "0001100101010000000100",
			1168 => "0000001001001011001001",
			1169 => "0000000001001011001001",
			1170 => "1111111001001011001001",
			1171 => "0001010111111100010100",
			1172 => "0001001000001000001000",
			1173 => "0010000101000100000100",
			1174 => "0000000001001011001001",
			1175 => "1111111001001011001001",
			1176 => "0001000011001100000100",
			1177 => "0000101001001011001001",
			1178 => "0011111100001100000100",
			1179 => "0000001001001011001001",
			1180 => "1111111001001011001001",
			1181 => "0001101001111100011100",
			1182 => "0010011010100100001000",
			1183 => "0010101001000100000100",
			1184 => "0000001001001011001001",
			1185 => "0000000001001011001001",
			1186 => "0011011010000100001100",
			1187 => "0011010110111100000100",
			1188 => "0000001001001011001001",
			1189 => "0001111011011100000100",
			1190 => "0000000001001011001001",
			1191 => "0000001001001011001001",
			1192 => "0000000111000000000100",
			1193 => "1111111001001011001001",
			1194 => "0000001001001011001001",
			1195 => "0001000000010100000100",
			1196 => "1111111001001011001001",
			1197 => "0010000111000100001000",
			1198 => "0011001111011100000100",
			1199 => "0000000001001011001001",
			1200 => "0000001001001011001001",
			1201 => "1111111001001011001001",
			1202 => "0011001011000000000100",
			1203 => "0000000001001101001101",
			1204 => "0001101001111100101100",
			1205 => "0001000011110000011100",
			1206 => "0010110000110100010000",
			1207 => "0001100100111100000100",
			1208 => "0000000001001101001101",
			1209 => "0000011010011000001000",
			1210 => "0001111011011100000100",
			1211 => "0000000001001101001101",
			1212 => "0000000001001101001101",
			1213 => "0000000001001101001101",
			1214 => "0010110110100000001000",
			1215 => "0000010100110100000100",
			1216 => "0000000001001101001101",
			1217 => "0000000001001101001101",
			1218 => "0000000001001101001101",
			1219 => "0010010100101100000100",
			1220 => "0000000001001101001101",
			1221 => "0000101101001000001000",
			1222 => "0001111000011000000100",
			1223 => "0000000001001101001101",
			1224 => "0000000001001101001101",
			1225 => "0000000001001101001101",
			1226 => "0011100011010100010000",
			1227 => "0000010100111100001100",
			1228 => "0000100110001100000100",
			1229 => "0000000001001101001101",
			1230 => "0010101010110000000100",
			1231 => "0000000001001101001101",
			1232 => "0000000001001101001101",
			1233 => "0000000001001101001101",
			1234 => "0000000001001101001101",
			1235 => "0000010111101000001000",
			1236 => "0001000000100000000100",
			1237 => "1111111001001111111001",
			1238 => "0000000001001111111001",
			1239 => "0000000111000000100100",
			1240 => "0011111000011100010100",
			1241 => "0001110001011000010000",
			1242 => "0010000101000100000100",
			1243 => "0000000001001111111001",
			1244 => "0001001110100100001000",
			1245 => "0010110000110100000100",
			1246 => "1111111001001111111001",
			1247 => "0000000001001111111001",
			1248 => "0000000001001111111001",
			1249 => "0000001001001111111001",
			1250 => "0000011010011000001000",
			1251 => "0001010010000000000100",
			1252 => "0000000001001111111001",
			1253 => "0000000001001111111001",
			1254 => "0011010110111100000100",
			1255 => "0000000001001111111001",
			1256 => "1111111001001111111001",
			1257 => "0001100101010000010000",
			1258 => "0010110100010000000100",
			1259 => "0000000001001111111001",
			1260 => "0001000011110000000100",
			1261 => "0000000001001111111001",
			1262 => "0001011100010000000100",
			1263 => "0000001001001111111001",
			1264 => "0000000001001111111001",
			1265 => "0001000000010100001100",
			1266 => "0010100110011000000100",
			1267 => "0000000001001111111001",
			1268 => "0000011001100100000100",
			1269 => "1111111001001111111001",
			1270 => "0000000001001111111001",
			1271 => "0000000011010000001000",
			1272 => "0010001011010100000100",
			1273 => "0000000001001111111001",
			1274 => "0000000001001111111001",
			1275 => "0001001011001000000100",
			1276 => "0000000001001111111001",
			1277 => "0000000001001111111001",
			1278 => "0011001011000000000100",
			1279 => "0000000001010001111101",
			1280 => "0011100110111000011000",
			1281 => "0000100010010100000100",
			1282 => "0000000001010001111101",
			1283 => "0010000111000100010000",
			1284 => "0000011011111100000100",
			1285 => "0000000001010001111101",
			1286 => "0011000111010000001000",
			1287 => "0010101000100100000100",
			1288 => "0000000001010001111101",
			1289 => "0000000001010001111101",
			1290 => "0000000001010001111101",
			1291 => "0000000001010001111101",
			1292 => "0011001010001100010100",
			1293 => "0010000001010100000100",
			1294 => "0000000001010001111101",
			1295 => "0010010111110100001100",
			1296 => "0001110101110100001000",
			1297 => "0000010100110100000100",
			1298 => "0000000001010001111101",
			1299 => "0000000001010001111101",
			1300 => "0000000001010001111101",
			1301 => "0000000001010001111101",
			1302 => "0010000110001000001100",
			1303 => "0001111011110100001000",
			1304 => "0000011100011000000100",
			1305 => "0000000001010001111101",
			1306 => "0000000001010001111101",
			1307 => "0000000001010001111101",
			1308 => "0000011001100100000100",
			1309 => "0000000001010001111101",
			1310 => "0000000001010001111101",
			1311 => "0000010100110100100000",
			1312 => "0001100100111100000100",
			1313 => "1111111001010101010001",
			1314 => "0011110110111000010000",
			1315 => "0001000111011100001000",
			1316 => "0011110110111000000100",
			1317 => "1111111001010101010001",
			1318 => "0000000001010101010001",
			1319 => "0000011101011100000100",
			1320 => "0000000001010101010001",
			1321 => "0000001001010101010001",
			1322 => "0001101000010000001000",
			1323 => "0000101000011100000100",
			1324 => "0000000001010101010001",
			1325 => "0000000001010101010001",
			1326 => "1111111001010101010001",
			1327 => "0000011100011000101000",
			1328 => "0001100100111100010100",
			1329 => "0000110001011100000100",
			1330 => "1111111001010101010001",
			1331 => "0001000011110000001100",
			1332 => "0001001110100100000100",
			1333 => "0000001001010101010001",
			1334 => "0001000101000000000100",
			1335 => "0000000001010101010001",
			1336 => "0000000001010101010001",
			1337 => "0000010001010101010001",
			1338 => "0001001110111000010000",
			1339 => "0011101000101000001000",
			1340 => "0010110010001000000100",
			1341 => "0000000001010101010001",
			1342 => "0000000001010101010001",
			1343 => "0001001000011100000100",
			1344 => "0000000001010101010001",
			1345 => "1111111001010101010001",
			1346 => "0000000001010101010001",
			1347 => "0010000110001000011100",
			1348 => "0011011010000100010100",
			1349 => "0001110111010000001100",
			1350 => "0011100110111000001000",
			1351 => "0000101011110000000100",
			1352 => "0000000001010101010001",
			1353 => "0000001001010101010001",
			1354 => "1111111001010101010001",
			1355 => "0001110111110000000100",
			1356 => "0000001001010101010001",
			1357 => "0000000001010101010001",
			1358 => "0011101110100100000100",
			1359 => "1111111001010101010001",
			1360 => "0000001001010101010001",
			1361 => "0001110101110100000100",
			1362 => "1111111001010101010001",
			1363 => "0000000001010101010001",
			1364 => "0010011010100000100100",
			1365 => "0001100100111100000100",
			1366 => "1111111001011000101101",
			1367 => "0011110010010100001100",
			1368 => "0010011011001100000100",
			1369 => "0000000001011000101101",
			1370 => "0001001010110100000100",
			1371 => "0000000001011000101101",
			1372 => "0000001001011000101101",
			1373 => "0000010111101000000100",
			1374 => "1111111001011000101101",
			1375 => "0000010001111000001000",
			1376 => "0001100101010000000100",
			1377 => "0000001001011000101101",
			1378 => "0000000001011000101101",
			1379 => "0001100101010000000100",
			1380 => "0000000001011000101101",
			1381 => "1111111001011000101101",
			1382 => "0000011100011000101000",
			1383 => "0000010100110100010100",
			1384 => "0001001000001000001000",
			1385 => "0001100100111100000100",
			1386 => "0000000001011000101101",
			1387 => "0000000001011000101101",
			1388 => "0001010011001000001000",
			1389 => "0010110100010000000100",
			1390 => "0000000001011000101101",
			1391 => "0000001001011000101101",
			1392 => "0000000001011000101101",
			1393 => "0010000101000100001000",
			1394 => "0000110001011100000100",
			1395 => "0000000001011000101101",
			1396 => "0000000001011000101101",
			1397 => "0000000010111100001000",
			1398 => "0010010010101100000100",
			1399 => "1111111001011000101101",
			1400 => "0000000001011000101101",
			1401 => "0000000001011000101101",
			1402 => "0001010111111100001000",
			1403 => "0011101101101100000100",
			1404 => "0000000001011000101101",
			1405 => "1111111001011000101101",
			1406 => "0011010110111100001000",
			1407 => "0011100011110000000100",
			1408 => "0000001001011000101101",
			1409 => "0000000001011000101101",
			1410 => "0001111011011100000100",
			1411 => "1111111001011000101101",
			1412 => "0000001010101100001000",
			1413 => "0010010011101000000100",
			1414 => "0000001001011000101101",
			1415 => "0000000001011000101101",
			1416 => "0010000111000100000100",
			1417 => "0000001001011000101101",
			1418 => "0000000001011000101101",
			1419 => "0000010001111000001100",
			1420 => "0000010101011100000100",
			1421 => "1111111001011011100001",
			1422 => "0001000111011100000100",
			1423 => "1111111001011011100001",
			1424 => "0000000001011011100001",
			1425 => "0000011101011000111100",
			1426 => "0011111000011100011100",
			1427 => "0011011010001000001000",
			1428 => "0010001011010100000100",
			1429 => "1111111001011011100001",
			1430 => "0000000001011011100001",
			1431 => "0011000001011000010000",
			1432 => "0011111111101000001000",
			1433 => "0011001001110100000100",
			1434 => "1111111001011011100001",
			1435 => "0000000001011011100001",
			1436 => "0011111000110100000100",
			1437 => "0000001001011011100001",
			1438 => "0000000001011011100001",
			1439 => "0000000001011011100001",
			1440 => "0001110110110100010100",
			1441 => "0001000100001100010000",
			1442 => "0011111000011100001000",
			1443 => "0000101000110100000100",
			1444 => "1111101001011011100001",
			1445 => "0000000001011011100001",
			1446 => "0010110010110100000100",
			1447 => "1111111001011011100001",
			1448 => "0000000001011011100001",
			1449 => "0000000001011011100001",
			1450 => "0001101001111100001000",
			1451 => "0000010100110100000100",
			1452 => "0000000001011011100001",
			1453 => "0000001001011011100001",
			1454 => "1111111001011011100001",
			1455 => "0010101000010100001000",
			1456 => "0000111110100100000100",
			1457 => "0000001001011011100001",
			1458 => "1111111001011011100001",
			1459 => "0001100100101100001000",
			1460 => "0010110001001000000100",
			1461 => "0000000001011011100001",
			1462 => "0000001001011011100001",
			1463 => "0000000001011011100001",
			1464 => "0010010100111100000100",
			1465 => "0000000001011101101101",
			1466 => "0001000011010100110000",
			1467 => "0001100100111100001100",
			1468 => "0010011010100100000100",
			1469 => "0000000001011101101101",
			1470 => "0010110100010000000100",
			1471 => "0000000001011101101101",
			1472 => "0000000001011101101101",
			1473 => "0000011100011000001000",
			1474 => "0011110010010100000100",
			1475 => "0000000001011101101101",
			1476 => "0000000001011101101101",
			1477 => "0010110110100000010000",
			1478 => "0010000101000100001000",
			1479 => "0001111011011100000100",
			1480 => "0000000001011101101101",
			1481 => "0000000001011101101101",
			1482 => "0000100011110000000100",
			1483 => "0000000001011101101101",
			1484 => "0000000001011101101101",
			1485 => "0010010011101000000100",
			1486 => "0000000001011101101101",
			1487 => "0011111000011100000100",
			1488 => "0000000001011101101101",
			1489 => "0000000001011101101101",
			1490 => "0010100101000100010000",
			1491 => "0011011001100000000100",
			1492 => "0000001001011101101101",
			1493 => "0011011010000100000100",
			1494 => "0000000001011101101101",
			1495 => "0010010011101000000100",
			1496 => "0000000001011101101101",
			1497 => "0000000001011101101101",
			1498 => "0000000001011101101101",
			1499 => "0011001010111000000100",
			1500 => "1111111001011111110001",
			1501 => "0001001011001000111000",
			1502 => "0001100101010000101000",
			1503 => "0001000011110000011000",
			1504 => "0010000001010100001100",
			1505 => "0010111011110100000100",
			1506 => "0000000001011111110001",
			1507 => "0001000110001100000100",
			1508 => "0000001001011111110001",
			1509 => "0000000001011111110001",
			1510 => "0000011101011000001000",
			1511 => "0011001010001100000100",
			1512 => "0000000001011111110001",
			1513 => "0000000001011111110001",
			1514 => "0000000001011111110001",
			1515 => "0011001000000000000100",
			1516 => "0000000001011111110001",
			1517 => "0011110011001100001000",
			1518 => "0000011011111100000100",
			1519 => "0000000001011111110001",
			1520 => "0000001001011111110001",
			1521 => "0000000001011111110001",
			1522 => "0000011101011000001000",
			1523 => "0001000011101100000100",
			1524 => "1111111001011111110001",
			1525 => "0000000001011111110001",
			1526 => "0010001111001000000100",
			1527 => "0000000001011111110001",
			1528 => "0000000001011111110001",
			1529 => "0010100101000100000100",
			1530 => "0000001001011111110001",
			1531 => "0000000001011111110001",
			1532 => "0000010100110101000000",
			1533 => "0000010100110100110000",
			1534 => "0000010101011100000100",
			1535 => "1111111001100010100101",
			1536 => "0011001001110100010100",
			1537 => "0000010101011100001000",
			1538 => "0001110110100100000100",
			1539 => "0000001001100010100101",
			1540 => "1111111001100010100101",
			1541 => "0011001000000000000100",
			1542 => "1111111001100010100101",
			1543 => "0000011110010100000100",
			1544 => "0000000001100010100101",
			1545 => "1111111001100010100101",
			1546 => "0001110111010000001100",
			1547 => "0001101000010000000100",
			1548 => "1111111001100010100101",
			1549 => "0000110110111000000100",
			1550 => "0000010001100010100101",
			1551 => "1111111001100010100101",
			1552 => "0011000001101000001000",
			1553 => "0000010111101000000100",
			1554 => "1111111001100010100101",
			1555 => "0000001001100010100101",
			1556 => "1111111001100010100101",
			1557 => "0001110111010000001000",
			1558 => "0011001001110100000100",
			1559 => "1111111001100010100101",
			1560 => "0000000001100010100101",
			1561 => "0000111110000000000100",
			1562 => "0000010001100010100101",
			1563 => "0000000001100010100101",
			1564 => "0011011100010100000100",
			1565 => "1111111001100010100101",
			1566 => "0001100100101100010100",
			1567 => "0001001001000000010000",
			1568 => "0010000110001000001100",
			1569 => "0001010111111100000100",
			1570 => "0000001001100010100101",
			1571 => "0000011100011000000100",
			1572 => "0000001001100010100101",
			1573 => "0000001001100010100101",
			1574 => "0000000001100010100101",
			1575 => "0000010001100010100101",
			1576 => "1111111001100010100101",
			1577 => "0000101101101100001000",
			1578 => "0000110001011100000100",
			1579 => "1111111001100101001001",
			1580 => "0000000001100101001001",
			1581 => "0011111000000100011000",
			1582 => "0011001010111000000100",
			1583 => "0000000001100101001001",
			1584 => "0011000001011000010000",
			1585 => "0010011011001100000100",
			1586 => "0000000001100101001001",
			1587 => "0001000110111000000100",
			1588 => "0000000001100101001001",
			1589 => "0001101111000000000100",
			1590 => "0000000001100101001001",
			1591 => "0000001001100101001001",
			1592 => "0000000001100101001001",
			1593 => "0000011101011000101000",
			1594 => "0010110110100000011100",
			1595 => "0001111011011100010000",
			1596 => "0001010011001000001000",
			1597 => "0001101001111100000100",
			1598 => "0000000001100101001001",
			1599 => "0000000001100101001001",
			1600 => "0000011101011000000100",
			1601 => "1111111001100101001001",
			1602 => "0000000001100101001001",
			1603 => "0000011100011000001000",
			1604 => "0011001111011100000100",
			1605 => "0000000001100101001001",
			1606 => "0000000001100101001001",
			1607 => "0000001001100101001001",
			1608 => "0010010011101000001000",
			1609 => "0001001101001000000100",
			1610 => "0000000001100101001001",
			1611 => "1111111001100101001001",
			1612 => "1111111001100101001001",
			1613 => "0010100110011100001000",
			1614 => "0001110000011100000100",
			1615 => "0000000001100101001001",
			1616 => "0000001001100101001001",
			1617 => "0000000001100101001001",
			1618 => "0000101100111000000100",
			1619 => "1111111001100111010101",
			1620 => "0001001011001000111000",
			1621 => "0001100101010000101100",
			1622 => "0001000011110000011100",
			1623 => "0000001010101100001100",
			1624 => "0001110111010000000100",
			1625 => "0000000001100111010101",
			1626 => "0000010100110100000100",
			1627 => "0000000001100111010101",
			1628 => "0000001001100111010101",
			1629 => "0001110110110100001000",
			1630 => "0000011101011000000100",
			1631 => "1111111001100111010101",
			1632 => "0000000001100111010101",
			1633 => "0001110101110100000100",
			1634 => "0000000001100111010101",
			1635 => "0000000001100111010101",
			1636 => "0011001000000000000100",
			1637 => "0000000001100111010101",
			1638 => "0011100110001100001000",
			1639 => "0000011011111100000100",
			1640 => "0000000001100111010101",
			1641 => "0000001001100111010101",
			1642 => "0000000001100111010101",
			1643 => "0000011101011000000100",
			1644 => "1111111001100111010101",
			1645 => "0010001111001000000100",
			1646 => "0000000001100111010101",
			1647 => "0000000001100111010101",
			1648 => "0010100101000100001000",
			1649 => "0001101000010000000100",
			1650 => "0000000001100111010101",
			1651 => "0000001001100111010101",
			1652 => "0000000001100111010101",
			1653 => "0010011010100000010000",
			1654 => "0010011001111100000100",
			1655 => "1111111001101010100001",
			1656 => "0001000010100100000100",
			1657 => "1111111001101010100001",
			1658 => "0001101001111100000100",
			1659 => "0000001001101010100001",
			1660 => "0000000001101010100001",
			1661 => "0001110001011000100100",
			1662 => "0011110010111000100000",
			1663 => "0001000010110000010000",
			1664 => "0010110000110100001100",
			1665 => "0010010011101000001000",
			1666 => "0001101111000000000100",
			1667 => "0000000001101010100001",
			1668 => "1111111001101010100001",
			1669 => "0000000001101010100001",
			1670 => "0000001001101010100001",
			1671 => "0001101001111100001100",
			1672 => "0010110100010000000100",
			1673 => "0000000001101010100001",
			1674 => "0000110110001100000100",
			1675 => "0000001001101010100001",
			1676 => "0000000001101010100001",
			1677 => "0000000001101010100001",
			1678 => "1111111001101010100001",
			1679 => "0001010110010000001100",
			1680 => "0010011010100100001000",
			1681 => "0010011010100100000100",
			1682 => "0000000001101010100001",
			1683 => "0000000001101010100001",
			1684 => "0000001001101010100001",
			1685 => "0001110110110100010000",
			1686 => "0001010110010000001000",
			1687 => "0010101000010100000100",
			1688 => "1111101001101010100001",
			1689 => "0000000001101010100001",
			1690 => "0001011110110100000100",
			1691 => "0000000001101010100001",
			1692 => "0000000001101010100001",
			1693 => "0010101010110000010000",
			1694 => "0000001010101100001000",
			1695 => "0000110101000000000100",
			1696 => "0000000001101010100001",
			1697 => "1111111001101010100001",
			1698 => "0010010010101100000100",
			1699 => "0000000001101010100001",
			1700 => "0000001001101010100001",
			1701 => "0010011000100100000100",
			1702 => "1111111001101010100001",
			1703 => "0000000001101010100001",
			1704 => "0010010100111100000100",
			1705 => "1111111001101100111101",
			1706 => "0011010110010000010100",
			1707 => "0001000111011100010000",
			1708 => "0010010111101100000100",
			1709 => "0000000001101100111101",
			1710 => "0011001001110100000100",
			1711 => "0000000001101100111101",
			1712 => "0011000110100100000100",
			1713 => "0000000001101100111101",
			1714 => "0000000001101100111101",
			1715 => "0000000001101100111101",
			1716 => "0010110000110100010000",
			1717 => "0000011010011000001100",
			1718 => "0001100100111100000100",
			1719 => "0000000001101100111101",
			1720 => "0011001111011100000100",
			1721 => "1111111001101100111101",
			1722 => "0000000001101100111101",
			1723 => "0000000001101100111101",
			1724 => "0011010111011000010000",
			1725 => "0000101101001000001100",
			1726 => "0000011101111100000100",
			1727 => "0000000001101100111101",
			1728 => "0011000001011000000100",
			1729 => "0000000001101100111101",
			1730 => "0000000001101100111101",
			1731 => "0000000001101100111101",
			1732 => "0010000110001000010000",
			1733 => "0000101000110100001000",
			1734 => "0000101000000100000100",
			1735 => "0000000001101100111101",
			1736 => "0000000001101100111101",
			1737 => "0000001010101100000100",
			1738 => "0000000001101100111101",
			1739 => "0000000001101100111101",
			1740 => "0000010100111100000100",
			1741 => "0000000001101100111101",
			1742 => "0000000001101100111101",
			1743 => "0011001011000000000100",
			1744 => "1111111001101111110001",
			1745 => "0010110110100000111000",
			1746 => "0010010010101100100100",
			1747 => "0011100110111000010100",
			1748 => "0010010101010000000100",
			1749 => "0000000001101111110001",
			1750 => "0001000010110000001000",
			1751 => "0001110111010000000100",
			1752 => "0000000001101111110001",
			1753 => "0000000001101111110001",
			1754 => "0001100101010000000100",
			1755 => "0000001001101111110001",
			1756 => "0000000001101111110001",
			1757 => "0001101000010000000100",
			1758 => "0000000001101111110001",
			1759 => "0001010110010000001000",
			1760 => "0001000100001100000100",
			1761 => "1111111001101111110001",
			1762 => "0000000001101111110001",
			1763 => "0000000001101111110001",
			1764 => "0011000001101000001100",
			1765 => "0011001001110100000100",
			1766 => "0000000001101111110001",
			1767 => "0001110001011000000100",
			1768 => "0000000001101111110001",
			1769 => "0000000001101111110001",
			1770 => "0010011000010100000100",
			1771 => "0000001001101111110001",
			1772 => "0000000001101111110001",
			1773 => "0010010011101000011000",
			1774 => "0010000001010100001000",
			1775 => "0010010011101000000100",
			1776 => "0000000001101111110001",
			1777 => "0000000001101111110001",
			1778 => "0011001111011100000100",
			1779 => "0000000001101111110001",
			1780 => "0001101000010000000100",
			1781 => "0000000001101111110001",
			1782 => "0011010111011000000100",
			1783 => "0000000001101111110001",
			1784 => "1111111001101111110001",
			1785 => "0010000111000100000100",
			1786 => "0000000001101111110001",
			1787 => "0000000001101111110001",
			1788 => "0000100011000000001000",
			1789 => "0011001001110100000100",
			1790 => "1111111001110010111101",
			1791 => "0000000001110010111101",
			1792 => "0000011101011001001000",
			1793 => "0011111000000100011100",
			1794 => "0010011010100100001100",
			1795 => "0001000011110100000100",
			1796 => "0000000001110010111101",
			1797 => "0010000001110100000100",
			1798 => "0000000001110010111101",
			1799 => "0000000001110010111101",
			1800 => "0011110010010100001000",
			1801 => "0011000001101000000100",
			1802 => "0000000001110010111101",
			1803 => "0000000001110010111101",
			1804 => "0011001001110100000100",
			1805 => "0000000001110010111101",
			1806 => "0000001001110010111101",
			1807 => "0000101000110100010000",
			1808 => "0001010110010000001100",
			1809 => "0000001010101100000100",
			1810 => "0000000001110010111101",
			1811 => "0011111000110100000100",
			1812 => "0000000001110010111101",
			1813 => "1111111001110010111101",
			1814 => "0000000001110010111101",
			1815 => "0010100110011000010000",
			1816 => "0010010011101000001000",
			1817 => "0010011010100000000100",
			1818 => "0000000001110010111101",
			1819 => "0000001001110010111101",
			1820 => "0010101000010100000100",
			1821 => "0000000001110010111101",
			1822 => "0000000001110010111101",
			1823 => "0011011100010000001000",
			1824 => "0000010100110100000100",
			1825 => "0000000001110010111101",
			1826 => "0000000001110010111101",
			1827 => "1111111001110010111101",
			1828 => "0011011010000100001100",
			1829 => "0001010111111100000100",
			1830 => "0000000001110010111101",
			1831 => "0011111001001100000100",
			1832 => "0000001001110010111101",
			1833 => "0000000001110010111101",
			1834 => "0010011000100100000100",
			1835 => "0000000001110010111101",
			1836 => "0010000001110100000100",
			1837 => "0000001001110010111101",
			1838 => "0000000001110010111101",
			1839 => "0000101101101100001000",
			1840 => "0010111010010100000100",
			1841 => "1111111001110110001001",
			1842 => "0000000001110110001001",
			1843 => "0000011100011000110100",
			1844 => "0001100101010000101000",
			1845 => "0001001000001000010100",
			1846 => "0010110000110100001100",
			1847 => "0001100100111100001000",
			1848 => "0001101111000000000100",
			1849 => "0000000001110110001001",
			1850 => "0000000001110110001001",
			1851 => "1111111001110110001001",
			1852 => "0000010100110100000100",
			1853 => "0000000001110110001001",
			1854 => "0000001001110110001001",
			1855 => "0010011011001100000100",
			1856 => "0000000001110110001001",
			1857 => "0001101000010000001000",
			1858 => "0001100100111100000100",
			1859 => "0000000001110110001001",
			1860 => "0000001001110110001001",
			1861 => "0000010111101000000100",
			1862 => "0000000001110110001001",
			1863 => "0000001001110110001001",
			1864 => "0001110111010000001000",
			1865 => "0001111111011100000100",
			1866 => "0000000001110110001001",
			1867 => "0000000001110110001001",
			1868 => "1111111001110110001001",
			1869 => "0001010111111100001100",
			1870 => "0000011010011000001000",
			1871 => "0001000011001100000100",
			1872 => "0000000001110110001001",
			1873 => "0000000001110110001001",
			1874 => "1111111001110110001001",
			1875 => "0011010110111100001100",
			1876 => "0000100010110000000100",
			1877 => "0000001001110110001001",
			1878 => "0001110101100100000100",
			1879 => "0000000001110110001001",
			1880 => "0000000001110110001001",
			1881 => "0001111011011100000100",
			1882 => "1111111001110110001001",
			1883 => "0000011101011000001000",
			1884 => "0000011101011000000100",
			1885 => "0000000001110110001001",
			1886 => "1111111001110110001001",
			1887 => "0010000111000100000100",
			1888 => "0000001001110110001001",
			1889 => "0000000001110110001001",
			1890 => "0000011001011000000100",
			1891 => "1111111001111000100101",
			1892 => "0000011101011001000100",
			1893 => "0000111110100100100100",
			1894 => "0000011100011000011100",
			1895 => "0001001001001100010000",
			1896 => "0011001000011000001000",
			1897 => "0001111011011100000100",
			1898 => "1111111001111000100101",
			1899 => "0000000001111000100101",
			1900 => "0010101001000100000100",
			1901 => "0000000001111000100101",
			1902 => "0000000001111000100101",
			1903 => "0001101001111100001000",
			1904 => "0000110010010100000100",
			1905 => "0000001001111000100101",
			1906 => "0000000001111000100101",
			1907 => "0000000001111000100101",
			1908 => "0001010101110000000100",
			1909 => "0000000001111000100101",
			1910 => "0000001001111000100101",
			1911 => "0001110110110100001100",
			1912 => "0000011010011000000100",
			1913 => "0000000001111000100101",
			1914 => "0000011101011000000100",
			1915 => "1111111001111000100101",
			1916 => "0000000001111000100101",
			1917 => "0010101001000100001000",
			1918 => "0000011101011000000100",
			1919 => "0000001001111000100101",
			1920 => "0000000001111000100101",
			1921 => "0010110010110100000100",
			1922 => "0000000001111000100101",
			1923 => "0011000111010000000100",
			1924 => "0000000001111000100101",
			1925 => "1111111001111000100101",
			1926 => "0010000111000100000100",
			1927 => "0000001001111000100101",
			1928 => "0000000001111000100101",
			1929 => "0000101101101100001000",
			1930 => "0010111010010100000100",
			1931 => "1111111001111011110011",
			1932 => "0000000001111011110011",
			1933 => "0000011010011001001100",
			1934 => "0011100110111000101100",
			1935 => "0001010111111100011000",
			1936 => "0000001111000100001100",
			1937 => "0011111000110100001000",
			1938 => "0010000101000100000100",
			1939 => "0000000001111011110011",
			1940 => "1111111001111011110011",
			1941 => "0000000001111011110011",
			1942 => "0011000100011000000100",
			1943 => "0000000001111011110011",
			1944 => "0010011011001100000100",
			1945 => "0000000001111011110011",
			1946 => "0000001001111011110011",
			1947 => "0010011010100100010000",
			1948 => "0010110000110100001000",
			1949 => "0011001000011000000100",
			1950 => "0000000001111011110011",
			1951 => "0000000001111011110011",
			1952 => "0000100110111000000100",
			1953 => "0000000001111011110011",
			1954 => "1111111001111011110011",
			1955 => "0000001001111011110011",
			1956 => "0001111011011100010100",
			1957 => "0001000100001100010000",
			1958 => "0010111110101100001000",
			1959 => "0011111000110100000100",
			1960 => "0000000001111011110011",
			1961 => "1111111001111011110011",
			1962 => "0000001000101100000100",
			1963 => "0000000001111011110011",
			1964 => "0000000001111011110011",
			1965 => "0000000001111011110011",
			1966 => "0010001100000100000100",
			1967 => "0000001001111011110011",
			1968 => "0010111110101100000100",
			1969 => "0000000001111011110011",
			1970 => "1111111001111011110011",
			1971 => "0011101000000100000100",
			1972 => "0000001001111011110011",
			1973 => "0000000111000000000100",
			1974 => "1111111001111011110011",
			1975 => "0010000111000100001000",
			1976 => "0011000001101000000100",
			1977 => "0000000001111011110011",
			1978 => "0000001001111011110011",
			1979 => "0000000001111011110011",
			1980 => "0000000001111011110101",
			1981 => "0010110010011100000100",
			1982 => "0000000001111100000001",
			1983 => "1111110001111100000001",
			1984 => "0001011111010100000100",
			1985 => "0000000001111100001101",
			1986 => "1111111001111100001101",
			1987 => "0001000101010100000100",
			1988 => "0000000001111100100001",
			1989 => "0001000001100100000100",
			1990 => "0000000001111100100001",
			1991 => "0000000001111100100001",
			1992 => "0011000111010000001000",
			1993 => "0011001010111000000100",
			1994 => "0000000001111100110101",
			1995 => "0000000001111100110101",
			1996 => "0000000001111100110101",
			1997 => "0001011111100100000100",
			1998 => "0000000001111101001001",
			1999 => "0011011000101000000100",
			2000 => "1111001001111101001001",
			2001 => "0000000001111101001001",
			2002 => "0001000111011100001000",
			2003 => "0010000110001000000100",
			2004 => "0000000001111101011101",
			2005 => "0000000001111101011101",
			2006 => "0000000001111101011101",
			2007 => "0011011100111000001100",
			2008 => "0001000000010100000100",
			2009 => "0000000001111101111001",
			2010 => "0001000001100100000100",
			2011 => "0000000001111101111001",
			2012 => "0000000001111101111001",
			2013 => "0000000001111101111001",
			2014 => "0001000101010100001000",
			2015 => "0001001110100100000100",
			2016 => "0000000001111110011101",
			2017 => "0000000001111110011101",
			2018 => "0001000001100100001000",
			2019 => "0001000011010100000100",
			2020 => "0000000001111110011101",
			2021 => "0000000001111110011101",
			2022 => "0000000001111110011101",
			2023 => "0010100110011000001100",
			2024 => "0010101000010100000100",
			2025 => "0000000001111111000001",
			2026 => "0001101111000000000100",
			2027 => "0000000001111111000001",
			2028 => "0000000001111111000001",
			2029 => "0001101000010000000100",
			2030 => "0000000001111111000001",
			2031 => "0000000001111111000001",
			2032 => "0000011100011000001100",
			2033 => "0010100110011100001000",
			2034 => "0010101000010100000100",
			2035 => "0000000001111111100101",
			2036 => "0000000001111111100101",
			2037 => "0000000001111111100101",
			2038 => "0010101010110000000100",
			2039 => "0000000001111111100101",
			2040 => "0000000001111111100101",
			2041 => "0011001011011100001100",
			2042 => "0001000100001100000100",
			2043 => "0000000010000000001001",
			2044 => "0001000001100100000100",
			2045 => "0000000010000000001001",
			2046 => "0000000010000000001001",
			2047 => "0001111011110100000100",
			2048 => "0000000010000000001001",
			2049 => "0000000010000000001001",
			2050 => "0010100110011000001100",
			2051 => "0010101000010100000100",
			2052 => "0000000010000000110101",
			2053 => "0001101111000000000100",
			2054 => "0000000010000000110101",
			2055 => "0000000010000000110101",
			2056 => "0001101000010000000100",
			2057 => "0000000010000000110101",
			2058 => "0000001000110000000100",
			2059 => "0000000010000000110101",
			2060 => "0000000010000000110101",
			2061 => "0010001011010100001100",
			2062 => "0000000111000000000100",
			2063 => "0000000010000001100001",
			2064 => "0000000011111100000100",
			2065 => "0000000010000001100001",
			2066 => "0000000010000001100001",
			2067 => "0000011001100100001000",
			2068 => "0000001011000100000100",
			2069 => "0000000010000001100001",
			2070 => "0000000010000001100001",
			2071 => "0000000010000001100001",
			2072 => "0001000111011100010000",
			2073 => "0010000110001000001100",
			2074 => "0001000101010100001000",
			2075 => "0001001110000000000100",
			2076 => "0000000010000010000101",
			2077 => "0000000010000010000101",
			2078 => "0000000010000010000101",
			2079 => "0000000010000010000101",
			2080 => "0000000010000010000101",
			2081 => "0001110001001000010000",
			2082 => "0001110001011000000100",
			2083 => "0000000010000010101001",
			2084 => "0010110000110100000100",
			2085 => "0000000010000010101001",
			2086 => "0011011001100000000100",
			2087 => "0000000010000010101001",
			2088 => "0000000010000010101001",
			2089 => "0000000010000010101001",
			2090 => "0000101000000100000100",
			2091 => "0000000010000011001101",
			2092 => "0000011111000000001100",
			2093 => "0001001001000000001000",
			2094 => "0010001001101000000100",
			2095 => "0000000010000011001101",
			2096 => "0000000010000011001101",
			2097 => "0000000010000011001101",
			2098 => "0000000010000011001101",
			2099 => "0010011010100100010000",
			2100 => "0001111000011000001000",
			2101 => "0011001010111000000100",
			2102 => "0000000010000100000001",
			2103 => "0000000010000100000001",
			2104 => "0001010001000000000100",
			2105 => "0000000010000100000001",
			2106 => "0000000010000100000001",
			2107 => "0011000001101000000100",
			2108 => "0000000010000100000001",
			2109 => "0001111011110100000100",
			2110 => "0000000010000100000001",
			2111 => "0000000010000100000001",
			2112 => "0001000100001100010000",
			2113 => "0001001100001100000100",
			2114 => "0000000010000100110101",
			2115 => "0000101000110100001000",
			2116 => "0010010011101000000100",
			2117 => "0000000010000100110101",
			2118 => "0000000010000100110101",
			2119 => "0000000010000100110101",
			2120 => "0010011001111100000100",
			2121 => "0000000010000100110101",
			2122 => "0001100100101100000100",
			2123 => "0000000010000100110101",
			2124 => "0000000010000100110101",
			2125 => "0011001011011100010100",
			2126 => "0000011100011000001000",
			2127 => "0011111111101000000100",
			2128 => "0000000010000101101001",
			2129 => "0000000010000101101001",
			2130 => "0001111011011100000100",
			2131 => "0000000010000101101001",
			2132 => "0000010100111100000100",
			2133 => "0000000010000101101001",
			2134 => "0000000010000101101001",
			2135 => "0010111111010000000100",
			2136 => "0000000010000101101001",
			2137 => "1111111010000101101001",
			2138 => "0011001011011100010100",
			2139 => "0010010010101100000100",
			2140 => "0000000010000110011101",
			2141 => "0001101000010000000100",
			2142 => "0000000010000110011101",
			2143 => "0010011001000100001000",
			2144 => "0001010101110000000100",
			2145 => "0000000010000110011101",
			2146 => "0000000010000110011101",
			2147 => "0000000010000110011101",
			2148 => "0010111111010000000100",
			2149 => "0000000010000110011101",
			2150 => "1111111010000110011101",
			2151 => "0010001111001000010100",
			2152 => "0011001001110100000100",
			2153 => "0000000010000111010001",
			2154 => "0000000010101000000100",
			2155 => "0000000010000111010001",
			2156 => "0011010111111100000100",
			2157 => "0000000010000111010001",
			2158 => "0011001011011100000100",
			2159 => "0000000010000111010001",
			2160 => "0000000010000111010001",
			2161 => "0000001011000100000100",
			2162 => "0000000010000111010001",
			2163 => "0000000010000111010001",
			2164 => "0001010000010000010100",
			2165 => "0010110000110100000100",
			2166 => "0000000010000111111101",
			2167 => "0001011110010000000100",
			2168 => "0000000010000111111101",
			2169 => "0011000001101000000100",
			2170 => "0000000010000111111101",
			2171 => "0011001011011100000100",
			2172 => "0000000010000111111101",
			2173 => "0000000010000111111101",
			2174 => "0000000010000111111101",
			2175 => "0001111011110100010100",
			2176 => "0010011001111100000100",
			2177 => "0000000010001000111001",
			2178 => "0000100110111000000100",
			2179 => "0000000010001000111001",
			2180 => "0010000111000100001000",
			2181 => "0001110001101000000100",
			2182 => "0000000010001000111001",
			2183 => "0000000010001000111001",
			2184 => "0000000010001000111001",
			2185 => "0001101000010000000100",
			2186 => "0000000010001000111001",
			2187 => "0010111101000100000100",
			2188 => "0000000010001000111001",
			2189 => "0000000010001000111001",
			2190 => "0001000000100000011000",
			2191 => "0000011101011000010000",
			2192 => "0000001010101100000100",
			2193 => "0000000010001001111101",
			2194 => "0001001001000000001000",
			2195 => "0010101000010100000100",
			2196 => "0000000010001001111101",
			2197 => "0000000010001001111101",
			2198 => "0000000010001001111101",
			2199 => "0001100100101100000100",
			2200 => "0000000010001001111101",
			2201 => "0000000010001001111101",
			2202 => "0010100101000100001000",
			2203 => "0000011001011000000100",
			2204 => "0000000010001001111101",
			2205 => "0000001010001001111101",
			2206 => "0000000010001001111101",
			2207 => "0001000000010100010100",
			2208 => "0001111011011100010000",
			2209 => "0011001111011100001100",
			2210 => "0000011011001100001000",
			2211 => "0010000101000100000100",
			2212 => "0000000010001011000001",
			2213 => "0000000010001011000001",
			2214 => "0000000010001011000001",
			2215 => "0000000010001011000001",
			2216 => "0000000010001011000001",
			2217 => "0010001111001000001100",
			2218 => "0000011011111100000100",
			2219 => "0000000010001011000001",
			2220 => "0000000010011000000100",
			2221 => "0000000010001011000001",
			2222 => "0000000010001011000001",
			2223 => "0000000010001011000001",
			2224 => "0001000000010100010100",
			2225 => "0000001010101100000100",
			2226 => "0000000010001100000101",
			2227 => "0010011000100100001100",
			2228 => "0001110111110000001000",
			2229 => "0010000001010100000100",
			2230 => "0000000010001100000101",
			2231 => "0000000010001100000101",
			2232 => "0000000010001100000101",
			2233 => "0000000010001100000101",
			2234 => "0010000111000100001100",
			2235 => "0000011011111100000100",
			2236 => "0000000010001100000101",
			2237 => "0000000010011000000100",
			2238 => "0000000010001100000101",
			2239 => "0000000010001100000101",
			2240 => "0000000010001100000101",
			2241 => "0001000000100000011100",
			2242 => "0000011101011000010000",
			2243 => "0010000101000100000100",
			2244 => "0000000010001101010001",
			2245 => "0001001001000000001000",
			2246 => "0000000001110100000100",
			2247 => "0000000010001101010001",
			2248 => "0000000010001101010001",
			2249 => "0000000010001101010001",
			2250 => "0010001111001000001000",
			2251 => "0011011110110100000100",
			2252 => "0000000010001101010001",
			2253 => "0000000010001101010001",
			2254 => "0000000010001101010001",
			2255 => "0010100101000100001000",
			2256 => "0000011001011000000100",
			2257 => "0000000010001101010001",
			2258 => "0000001010001101010001",
			2259 => "0000000010001101010001",
			2260 => "0001000000010100011100",
			2261 => "0010110000110100010000",
			2262 => "0000000001110100000100",
			2263 => "0000000010001110100101",
			2264 => "0010010011101000001000",
			2265 => "0001110110110100000100",
			2266 => "0000000010001110100101",
			2267 => "0000000010001110100101",
			2268 => "0000000010001110100101",
			2269 => "0010100001010000001000",
			2270 => "0001101111000000000100",
			2271 => "0000000010001110100101",
			2272 => "0000000010001110100101",
			2273 => "0000000010001110100101",
			2274 => "0010100101000100001100",
			2275 => "0010011011001100000100",
			2276 => "0000000010001110100101",
			2277 => "0001111111011100000100",
			2278 => "0000000010001110100101",
			2279 => "0000000010001110100101",
			2280 => "0000000010001110100101",
			2281 => "0011001011011100011000",
			2282 => "0010101000010100000100",
			2283 => "0000000010001111100001",
			2284 => "0010011011001100000100",
			2285 => "0000000010001111100001",
			2286 => "0010100101000100001100",
			2287 => "0010011000010100001000",
			2288 => "0011001010111000000100",
			2289 => "0000000010001111100001",
			2290 => "0000000010001111100001",
			2291 => "0000000010001111100001",
			2292 => "0000000010001111100001",
			2293 => "0010000110001000000100",
			2294 => "0000000010001111100001",
			2295 => "1111111010001111100001",
			2296 => "0001000011011000011100",
			2297 => "0010011010100100000100",
			2298 => "0000000010010000101101",
			2299 => "0000111110100100001100",
			2300 => "0010111101000100001000",
			2301 => "0011011100010100000100",
			2302 => "0000000010010000101101",
			2303 => "0000000010010000101101",
			2304 => "0000000010010000101101",
			2305 => "0010011000100100001000",
			2306 => "0010001001101000000100",
			2307 => "0000000010010000101101",
			2308 => "0000000010010000101101",
			2309 => "0000000010010000101101",
			2310 => "0010100101000100001000",
			2311 => "0001101000010000000100",
			2312 => "0000000010010000101101",
			2313 => "0000001010010000101101",
			2314 => "0000000010010000101101",
			2315 => "0001110001001000011000",
			2316 => "0011001000011000000100",
			2317 => "0000000010010001100001",
			2318 => "0001100100101100010000",
			2319 => "0011100001011100000100",
			2320 => "0000000010010001100001",
			2321 => "0000101000110100000100",
			2322 => "0000000010010001100001",
			2323 => "0010100101000100000100",
			2324 => "0000000010010001100001",
			2325 => "0000000010010001100001",
			2326 => "0000000010010001100001",
			2327 => "0000000010010001100001",
			2328 => "0011111111101000010000",
			2329 => "0000011001011000000100",
			2330 => "0000000010010010101101",
			2331 => "0000101100111000000100",
			2332 => "0000000010010010101101",
			2333 => "0000011010011000000100",
			2334 => "0000000010010010101101",
			2335 => "0000000010010010101101",
			2336 => "0010000001010100000100",
			2337 => "0000000010010010101101",
			2338 => "0000111011110000000100",
			2339 => "0000000010010010101101",
			2340 => "0001100100111100000100",
			2341 => "0000000010010010101101",
			2342 => "0001001110100100000100",
			2343 => "0000000010010010101101",
			2344 => "0010101000010100000100",
			2345 => "0000000010010010101101",
			2346 => "0000000010010010101101",
			2347 => "0010100110011000011000",
			2348 => "0010101000010100000100",
			2349 => "0000000010010100000001",
			2350 => "0011001001110100000100",
			2351 => "0000000010010100000001",
			2352 => "0001011100010000001100",
			2353 => "0001001000011100000100",
			2354 => "0000000010010100000001",
			2355 => "0000011110010100000100",
			2356 => "0000000010010100000001",
			2357 => "0000001010010100000001",
			2358 => "0000000010010100000001",
			2359 => "0001001011001000001000",
			2360 => "0010000110001000000100",
			2361 => "0000000010010100000001",
			2362 => "0000000010010100000001",
			2363 => "0010100101000100001000",
			2364 => "0010101100011100000100",
			2365 => "0000000010010100000001",
			2366 => "0000000010010100000001",
			2367 => "0000000010010100000001",
			2368 => "0001001001000000100000",
			2369 => "0010000001010100010000",
			2370 => "0010111011110100000100",
			2371 => "0000000010010101011101",
			2372 => "0000111100001100001000",
			2373 => "0000010100110100000100",
			2374 => "0000000010010101011101",
			2375 => "0000000010010101011101",
			2376 => "0000000010010101011101",
			2377 => "0000011101011000001100",
			2378 => "0001000011101100001000",
			2379 => "0000001010101100000100",
			2380 => "0000000010010101011101",
			2381 => "0000000010010101011101",
			2382 => "0000000010010101011101",
			2383 => "0000000010010101011101",
			2384 => "0010000001110100001100",
			2385 => "0000000011010000000100",
			2386 => "0000000010010101011101",
			2387 => "0000010101011100000100",
			2388 => "0000000010010101011101",
			2389 => "0000000010010101011101",
			2390 => "0000000010010101011101",
			2391 => "0001000000010100100000",
			2392 => "0010110000110100010100",
			2393 => "0010000101000100000100",
			2394 => "0000000010010110111001",
			2395 => "0000011010011000001100",
			2396 => "0001110110110100001000",
			2397 => "0010101000100100000100",
			2398 => "0000000010010110111001",
			2399 => "0000000010010110111001",
			2400 => "0000000010010110111001",
			2401 => "0000000010010110111001",
			2402 => "0010100001010000001000",
			2403 => "0001101111000000000100",
			2404 => "0000000010010110111001",
			2405 => "0000000010010110111001",
			2406 => "0000000010010110111001",
			2407 => "0010001111001000001100",
			2408 => "0011001000000000000100",
			2409 => "0000000010010110111001",
			2410 => "0000000010011000000100",
			2411 => "0000000010010110111001",
			2412 => "0000000010010110111001",
			2413 => "0000000010010110111001",
			2414 => "0010110101110100010100",
			2415 => "0011001010111000000100",
			2416 => "0000000010011000010101",
			2417 => "0000000010011000000100",
			2418 => "0000000010011000010101",
			2419 => "0001100101010000001000",
			2420 => "0010011011001100000100",
			2421 => "0000000010011000010101",
			2422 => "0000000010011000010101",
			2423 => "0000000010011000010101",
			2424 => "0000011010011000010100",
			2425 => "0010000101000100000100",
			2426 => "0000000010011000010101",
			2427 => "0000110101000000001100",
			2428 => "0010010011101000001000",
			2429 => "0001011001010000000100",
			2430 => "0000000010011000010101",
			2431 => "0000000010011000010101",
			2432 => "0000000010011000010101",
			2433 => "0000000010011000010101",
			2434 => "0010000111000100000100",
			2435 => "0000000010011000010101",
			2436 => "0000000010011000010101",
			2437 => "0001101001111100011100",
			2438 => "0010010100111100000100",
			2439 => "0000000010011001100001",
			2440 => "0011001011011100010100",
			2441 => "0001101000010000000100",
			2442 => "0000000010011001100001",
			2443 => "0000100011110000001100",
			2444 => "0011011010000100001000",
			2445 => "0001100101010000000100",
			2446 => "0000000010011001100001",
			2447 => "0000000010011001100001",
			2448 => "0000000010011001100001",
			2449 => "0000000010011001100001",
			2450 => "0000000010011001100001",
			2451 => "0010000110001000000100",
			2452 => "0000000010011001100001",
			2453 => "0011111000011100000100",
			2454 => "0000000010011001100001",
			2455 => "0000000010011001100001",
			2456 => "0010000110001000011100",
			2457 => "0011011010000100011000",
			2458 => "0000100010010100000100",
			2459 => "0000000010011010101101",
			2460 => "0011000100000100010000",
			2461 => "0010011001111100000100",
			2462 => "0000000010011010101101",
			2463 => "0011100010111000001000",
			2464 => "0011001001110100000100",
			2465 => "0000000010011010101101",
			2466 => "0000000010011010101101",
			2467 => "0000000010011010101101",
			2468 => "0000000010011010101101",
			2469 => "0000000010011010101101",
			2470 => "0000100110111000000100",
			2471 => "0000000010011010101101",
			2472 => "0011100011010100000100",
			2473 => "0000000010011010101101",
			2474 => "0000000010011010101101",
			2475 => "0010001100000100011100",
			2476 => "0010111110101100010000",
			2477 => "0000011010011000001100",
			2478 => "0000001010101100000100",
			2479 => "0000000010011100100001",
			2480 => "0000001000110000000100",
			2481 => "0000000010011100100001",
			2482 => "0000000010011100100001",
			2483 => "0000000010011100100001",
			2484 => "0000011101011000001000",
			2485 => "0010011010100100000100",
			2486 => "0000000010011100100001",
			2487 => "0000000010011100100001",
			2488 => "0000000010011100100001",
			2489 => "0001000000010100001100",
			2490 => "0010011000100100001000",
			2491 => "0010001001101000000100",
			2492 => "0000000010011100100001",
			2493 => "0000000010011100100001",
			2494 => "0000000010011100100001",
			2495 => "0010000001110100010000",
			2496 => "0001100100101100001100",
			2497 => "0010111111011100000100",
			2498 => "0000000010011100100001",
			2499 => "0000000010011000000100",
			2500 => "0000000010011100100001",
			2501 => "0000000010011100100001",
			2502 => "0000000010011100100001",
			2503 => "0000000010011100100001",
			2504 => "0011100110111100001100",
			2505 => "0000011001011000000100",
			2506 => "0000000010011101111101",
			2507 => "0001001111100000000100",
			2508 => "0000000010011101111101",
			2509 => "0000001010011101111101",
			2510 => "0001101000010000001100",
			2511 => "0001111111011100000100",
			2512 => "0000000010011101111101",
			2513 => "0010011010100000000100",
			2514 => "0000000010011101111101",
			2515 => "0000000010011101111101",
			2516 => "0011111110000000000100",
			2517 => "0000000010011101111101",
			2518 => "0000011101011000010000",
			2519 => "0011101000000100001100",
			2520 => "0010111011110100000100",
			2521 => "0000000010011101111101",
			2522 => "0010000001010100000100",
			2523 => "0000000010011101111101",
			2524 => "0000000010011101111101",
			2525 => "0000000010011101111101",
			2526 => "0000000010011101111101",
			2527 => "0011111111101000010000",
			2528 => "0011011110101100000100",
			2529 => "0000000010011111010001",
			2530 => "0000101101101100000100",
			2531 => "0000000010011111010001",
			2532 => "0001101111000000000100",
			2533 => "0000000010011111010001",
			2534 => "0000000010011111010001",
			2535 => "0010101000010100000100",
			2536 => "0000000010011111010001",
			2537 => "0011100011010100010100",
			2538 => "0010110101110100000100",
			2539 => "0000000010011111010001",
			2540 => "0001001110100100000100",
			2541 => "0000000010011111010001",
			2542 => "0000001010101100000100",
			2543 => "0000000010011111010001",
			2544 => "0000110011101100000100",
			2545 => "0000000010011111010001",
			2546 => "0000000010011111010001",
			2547 => "0000000010011111010001",
			2548 => "0011100110111100001100",
			2549 => "0000011001011000000100",
			2550 => "0000000010100000110101",
			2551 => "0001001111100000000100",
			2552 => "0000000010100000110101",
			2553 => "0000001010100000110101",
			2554 => "0010000111000100100000",
			2555 => "0000101000110100010000",
			2556 => "0000001010101100000100",
			2557 => "0000000010100000110101",
			2558 => "0011111000000100000100",
			2559 => "0000000010100000110101",
			2560 => "0001001110100100000100",
			2561 => "0000000010100000110101",
			2562 => "0000000010100000110101",
			2563 => "0011001001110100000100",
			2564 => "0000000010100000110101",
			2565 => "0001001100001100000100",
			2566 => "0000000010100000110101",
			2567 => "0011001011011100000100",
			2568 => "0000000010100000110101",
			2569 => "0000000010100000110101",
			2570 => "0010110010001000000100",
			2571 => "0000000010100000110101",
			2572 => "0000000010100000110101",
			2573 => "0000010100110100010100",
			2574 => "0001000111011100000100",
			2575 => "0000000010100010101001",
			2576 => "0010000001110100001100",
			2577 => "0000000000111000000100",
			2578 => "0000000010100010101001",
			2579 => "0000011001011000000100",
			2580 => "0000000010100010101001",
			2581 => "0000000010100010101001",
			2582 => "0000000010100010101001",
			2583 => "0000110110001100001100",
			2584 => "0011000100000100001000",
			2585 => "0001110111010000000100",
			2586 => "0000000010100010101001",
			2587 => "0000000010100010101001",
			2588 => "0000000010100010101001",
			2589 => "0011000111010000010000",
			2590 => "0011110110001100000100",
			2591 => "0000000010100010101001",
			2592 => "0010101001000100000100",
			2593 => "0000000010100010101001",
			2594 => "0000011011001100000100",
			2595 => "0000000010100010101001",
			2596 => "0000000010100010101001",
			2597 => "0000010100111100001000",
			2598 => "0010010010101100000100",
			2599 => "0000000010100010101001",
			2600 => "0000000010100010101001",
			2601 => "0000000010100010101001",
			2602 => "0001000011011000101000",
			2603 => "0000011010011000011000",
			2604 => "0001111011011100010100",
			2605 => "0001000000010100010000",
			2606 => "0010000101000100000100",
			2607 => "0000000010100100001101",
			2608 => "0010111110101100001000",
			2609 => "0010101000100100000100",
			2610 => "0000000010100100001101",
			2611 => "0000000010100100001101",
			2612 => "0000000010100100001101",
			2613 => "0000000010100100001101",
			2614 => "0000000010100100001101",
			2615 => "0001111011110100001100",
			2616 => "0001110111010000000100",
			2617 => "0000000010100100001101",
			2618 => "0010000110001000000100",
			2619 => "0000000010100100001101",
			2620 => "0000000010100100001101",
			2621 => "0000000010100100001101",
			2622 => "0010100101000100001000",
			2623 => "0001101000010000000100",
			2624 => "0000000010100100001101",
			2625 => "0000001010100100001101",
			2626 => "0000000010100100001101",
			2627 => "0011001001110100001000",
			2628 => "0010100110011100000100",
			2629 => "0000000010100101101001",
			2630 => "0000000010100101101001",
			2631 => "0011010111011000010000",
			2632 => "0001010101110000000100",
			2633 => "0000000010100101101001",
			2634 => "0011000001011000001000",
			2635 => "0000010111101000000100",
			2636 => "0000000010100101101001",
			2637 => "0000000010100101101001",
			2638 => "0000000010100101101001",
			2639 => "0001110100010000010100",
			2640 => "0000011010011000000100",
			2641 => "0000000010100101101001",
			2642 => "0011000111010000001100",
			2643 => "0001010110010000000100",
			2644 => "0000000010100101101001",
			2645 => "0011010110111100000100",
			2646 => "0000000010100101101001",
			2647 => "0000000010100101101001",
			2648 => "0000000010100101101001",
			2649 => "0000000010100101101001",
			2650 => "0001011110000100010000",
			2651 => "0011001010111000000100",
			2652 => "0000000010100111010101",
			2653 => "0001001111100000000100",
			2654 => "0000000010100111010101",
			2655 => "0010001101010000000100",
			2656 => "0000001010100111010101",
			2657 => "0000000010100111010101",
			2658 => "0000011010011000011000",
			2659 => "0001100100111100000100",
			2660 => "0000000010100111010101",
			2661 => "0001111111011100000100",
			2662 => "0000000010100111010101",
			2663 => "0010010011101000001100",
			2664 => "0001011110110100001000",
			2665 => "0010000101000100000100",
			2666 => "0000000010100111010101",
			2667 => "0000000010100111010101",
			2668 => "0000000010100111010101",
			2669 => "0000000010100111010101",
			2670 => "0001100100101100001100",
			2671 => "0001110111010000000100",
			2672 => "0000000010100111010101",
			2673 => "0010101000010100000100",
			2674 => "0000000010100111010101",
			2675 => "0000000010100111010101",
			2676 => "0000000010100111010101",
			2677 => "0000011100011000101100",
			2678 => "0010011010100100011100",
			2679 => "0000010101011100000100",
			2680 => "1111111010101001010001",
			2681 => "0001111000011000001000",
			2682 => "0010011000010000000100",
			2683 => "0000000010101001010001",
			2684 => "1111111010101001010001",
			2685 => "0011101111101000001100",
			2686 => "0001101000010000000100",
			2687 => "1111111010101001010001",
			2688 => "0011001000011000000100",
			2689 => "0000100010101001010001",
			2690 => "0000000010101001010001",
			2691 => "1111111010101001010001",
			2692 => "0001110111010000001000",
			2693 => "0011001001110100000100",
			2694 => "1111111010101001010001",
			2695 => "0000000010101001010001",
			2696 => "0001100101010000000100",
			2697 => "0000011010101001010001",
			2698 => "0000000010101001010001",
			2699 => "0010111011110100000100",
			2700 => "1111111010101001010001",
			2701 => "0010000111000100001100",
			2702 => "0001110111010000000100",
			2703 => "0000001010101001010001",
			2704 => "0011001011011100000100",
			2705 => "0000010010101001010001",
			2706 => "0000001010101001010001",
			2707 => "1111111010101001010001",
			2708 => "0000111111100100010000",
			2709 => "0010011011001100000100",
			2710 => "0000000010101011000101",
			2711 => "0001001111100000000100",
			2712 => "0000000010101011000101",
			2713 => "0011000001111100000100",
			2714 => "0000000010101011000101",
			2715 => "0000001010101011000101",
			2716 => "0001101000010000010100",
			2717 => "0011001001110100000100",
			2718 => "0000000010101011000101",
			2719 => "0011000100000100001100",
			2720 => "0010111011110100000100",
			2721 => "0000000010101011000101",
			2722 => "0010011010100100000100",
			2723 => "0000000010101011000101",
			2724 => "0000000010101011000101",
			2725 => "0000000010101011000101",
			2726 => "0011111110000000000100",
			2727 => "0000000010101011000101",
			2728 => "0010010111110100010000",
			2729 => "0010111011110100000100",
			2730 => "0000000010101011000101",
			2731 => "0010000001010100000100",
			2732 => "0000000010101011000101",
			2733 => "0001001110100100000100",
			2734 => "0000000010101011000101",
			2735 => "0000000010101011000101",
			2736 => "0000000010101011000101",
			2737 => "0011111111101000011000",
			2738 => "0000011001011000000100",
			2739 => "0000000010101100101001",
			2740 => "0000101101101100000100",
			2741 => "0000000010101100101001",
			2742 => "0001100101010000001100",
			2743 => "0001101111000000000100",
			2744 => "0000000010101100101001",
			2745 => "0010010010101100000100",
			2746 => "0000000010101100101001",
			2747 => "0000000010101100101001",
			2748 => "0000000010101100101001",
			2749 => "0010000001010100000100",
			2750 => "0000000010101100101001",
			2751 => "0011100011010100010100",
			2752 => "0010110101110100000100",
			2753 => "0000000010101100101001",
			2754 => "0010101000010100000100",
			2755 => "0000000010101100101001",
			2756 => "0001001000011100000100",
			2757 => "0000000010101100101001",
			2758 => "0000001010101100000100",
			2759 => "0000000010101100101001",
			2760 => "0000000010101100101001",
			2761 => "0000000010101100101001",
			2762 => "0011101101101100011000",
			2763 => "0011001010111000000100",
			2764 => "0000000010101110100101",
			2765 => "0001101001111100010000",
			2766 => "0000101101101100000100",
			2767 => "0000000010101110100101",
			2768 => "0001101001100100000100",
			2769 => "0000000010101110100101",
			2770 => "0011001000011000000100",
			2771 => "0000001010101110100101",
			2772 => "0000000010101110100101",
			2773 => "0000000010101110100101",
			2774 => "0000011010011000011000",
			2775 => "0000110101000000010100",
			2776 => "0010101000100100000100",
			2777 => "0000000010101110100101",
			2778 => "0010010011101000001100",
			2779 => "0010000101000100000100",
			2780 => "0000000010101110100101",
			2781 => "0001100100111100000100",
			2782 => "0000000010101110100101",
			2783 => "0000000010101110100101",
			2784 => "0000000010101110100101",
			2785 => "0000000010101110100101",
			2786 => "0010000111000100001100",
			2787 => "0000001010101100000100",
			2788 => "0000000010101110100101",
			2789 => "0010111010010100000100",
			2790 => "0000000010101110100101",
			2791 => "0000000010101110100101",
			2792 => "0000000010101110100101",
			2793 => "0000011100011000110100",
			2794 => "0010011010100100100100",
			2795 => "0000010101011100000100",
			2796 => "1111111010110000110001",
			2797 => "0011001001110100010000",
			2798 => "0010011000010000000100",
			2799 => "0000000010110000110001",
			2800 => "0011001000000000000100",
			2801 => "1111111010110000110001",
			2802 => "0011001000000000000100",
			2803 => "0000000010110000110001",
			2804 => "1111111010110000110001",
			2805 => "0011101111101000001100",
			2806 => "0010010100101100000100",
			2807 => "1111111010110000110001",
			2808 => "0000101000000100000100",
			2809 => "1111111010110000110001",
			2810 => "0000010010110000110001",
			2811 => "1111111010110000110001",
			2812 => "0010111011110100001000",
			2813 => "0011001001110100000100",
			2814 => "1111111010110000110001",
			2815 => "0000000010110000110001",
			2816 => "0001100101010000000100",
			2817 => "0000010010110000110001",
			2818 => "0000000010110000110001",
			2819 => "0010111011110100000100",
			2820 => "1111111010110000110001",
			2821 => "0010000111000100001100",
			2822 => "0011001001110100000100",
			2823 => "0000001010110000110001",
			2824 => "0011001011011100000100",
			2825 => "0000001010110000110001",
			2826 => "0000001010110000110001",
			2827 => "1111111010110000110001",
			2828 => "0010011010100000010000",
			2829 => "0000100110111000000100",
			2830 => "1111111010110011001101",
			2831 => "0000101110100100001000",
			2832 => "0001000100001100000100",
			2833 => "0000000010110011001101",
			2834 => "0000000010110011001101",
			2835 => "1111111010110011001101",
			2836 => "0001000011110000101000",
			2837 => "0010110000110100010000",
			2838 => "0010101000100100000100",
			2839 => "0000000010110011001101",
			2840 => "0000011010011000001000",
			2841 => "0000010100110100000100",
			2842 => "0000000010110011001101",
			2843 => "1111111010110011001101",
			2844 => "0000000010110011001101",
			2845 => "0000111110100100000100",
			2846 => "0000001010110011001101",
			2847 => "0011101110000000001000",
			2848 => "0011101110000000000100",
			2849 => "0000000010110011001101",
			2850 => "1111111010110011001101",
			2851 => "0001111011011100000100",
			2852 => "0000000010110011001101",
			2853 => "0001001100001100000100",
			2854 => "0000000010110011001101",
			2855 => "0000001010110011001101",
			2856 => "0010101010110000001100",
			2857 => "0010110100010000000100",
			2858 => "0000000010110011001101",
			2859 => "0010111100100100000100",
			2860 => "0000001010110011001101",
			2861 => "0000000010110011001101",
			2862 => "0001000011010100000100",
			2863 => "1111111010110011001101",
			2864 => "0010000111000100000100",
			2865 => "0000001010110011001101",
			2866 => "0000000010110011001101",
			2867 => "0010010100111100000100",
			2868 => "0000000010110101001001",
			2869 => "0011111100001100100000",
			2870 => "0010110110100000010100",
			2871 => "0001101001111100010000",
			2872 => "0010000001010100000100",
			2873 => "0000000010110101001001",
			2874 => "0000100010010100000100",
			2875 => "0000000010110101001001",
			2876 => "0011001010111000000100",
			2877 => "0000000010110101001001",
			2878 => "0000000010110101001001",
			2879 => "0000000010110101001001",
			2880 => "0001101000010000000100",
			2881 => "0000000010110101001001",
			2882 => "0010000001010100000100",
			2883 => "0000000010110101001001",
			2884 => "0000000010110101001001",
			2885 => "0010011000100100010000",
			2886 => "0001110111110000001100",
			2887 => "0011101000011100000100",
			2888 => "0000000010110101001001",
			2889 => "0001100100111100000100",
			2890 => "0000000010110101001001",
			2891 => "0000000010110101001001",
			2892 => "0000000010110101001001",
			2893 => "0001100100101100001000",
			2894 => "0011001010011100000100",
			2895 => "0000000010110101001001",
			2896 => "0000000010110101001001",
			2897 => "0000000010110101001001",
			2898 => "0010011010100100100000",
			2899 => "0001100100111100001000",
			2900 => "0010011010100100000100",
			2901 => "1111111010111000000101",
			2902 => "0000000010111000000101",
			2903 => "0011101111101000010100",
			2904 => "0001001110111000000100",
			2905 => "1111111010111000000101",
			2906 => "0001101000010000001000",
			2907 => "0011000100011000000100",
			2908 => "0000000010111000000101",
			2909 => "0000001010111000000101",
			2910 => "0010010111101100000100",
			2911 => "1111111010111000000101",
			2912 => "0000000010111000000101",
			2913 => "1111111010111000000101",
			2914 => "0010110001001000011100",
			2915 => "0001000011110000010000",
			2916 => "0001100100111100001000",
			2917 => "0001010101110000000100",
			2918 => "1111111010111000000101",
			2919 => "0000001010111000000101",
			2920 => "0000011010011000000100",
			2921 => "1111111010111000000101",
			2922 => "0000000010111000000101",
			2923 => "0011100110111000000100",
			2924 => "0000001010111000000101",
			2925 => "0010010011101000000100",
			2926 => "1111111010111000000101",
			2927 => "0000000010111000000101",
			2928 => "0010110110100000010000",
			2929 => "0001101001111100001100",
			2930 => "0011000100000100000100",
			2931 => "0000001010111000000101",
			2932 => "0011000100000100000100",
			2933 => "0000000010111000000101",
			2934 => "0000001010111000000101",
			2935 => "0000000010111000000101",
			2936 => "0000001010101100001000",
			2937 => "0011111000011100000100",
			2938 => "0000001010111000000101",
			2939 => "1111111010111000000101",
			2940 => "0011101011110000000100",
			2941 => "1111111010111000000101",
			2942 => "0001100100101100000100",
			2943 => "0000001010111000000101",
			2944 => "1111111010111000000101",
			2945 => "0010010100101100000100",
			2946 => "0000000010111010001001",
			2947 => "0011111110100100100000",
			2948 => "0000101011110000010000",
			2949 => "0001110001011000001100",
			2950 => "0010000101000100000100",
			2951 => "0000000010111010001001",
			2952 => "0000001111000100000100",
			2953 => "0000000010111010001001",
			2954 => "0000000010111010001001",
			2955 => "0000000010111010001001",
			2956 => "0001111011011100001100",
			2957 => "0001101001111100001000",
			2958 => "0011011010001000000100",
			2959 => "0000000010111010001001",
			2960 => "0000000010111010001001",
			2961 => "0000000010111010001001",
			2962 => "0000000010111010001001",
			2963 => "0001111011011100010000",
			2964 => "0010010111110100001100",
			2965 => "0001000100001100001000",
			2966 => "0000011011001100000100",
			2967 => "0000000010111010001001",
			2968 => "0000000010111010001001",
			2969 => "0000000010111010001001",
			2970 => "0000000010111010001001",
			2971 => "0010000111000100001100",
			2972 => "0001001100001100000100",
			2973 => "0000000010111010001001",
			2974 => "0000010100110100000100",
			2975 => "0000000010111010001001",
			2976 => "0000000010111010001001",
			2977 => "0000000010111010001001",
			2978 => "0010011010100000010100",
			2979 => "0001100100111100000100",
			2980 => "1111111010111100110101",
			2981 => "0011110110111000001100",
			2982 => "0011001010111000000100",
			2983 => "0000000010111100110101",
			2984 => "0001001001001100000100",
			2985 => "0000000010111100110101",
			2986 => "0000000010111100110101",
			2987 => "1111111010111100110101",
			2988 => "0001000011110000101000",
			2989 => "0010110000110100010000",
			2990 => "0001100100111100001000",
			2991 => "0001010101110000000100",
			2992 => "0000000010111100110101",
			2993 => "0000000010111100110101",
			2994 => "0000011010011000000100",
			2995 => "1111111010111100110101",
			2996 => "0000000010111100110101",
			2997 => "0011111000011100000100",
			2998 => "0000001010111100110101",
			2999 => "0010010011101000001000",
			3000 => "0011000100000100000100",
			3001 => "0000000010111100110101",
			3002 => "0000000010111100110101",
			3003 => "0010000001010100001000",
			3004 => "0011010110111100000100",
			3005 => "0000000010111100110101",
			3006 => "1111111010111100110101",
			3007 => "0000000010111100110101",
			3008 => "0001101001111100001100",
			3009 => "0010110100010000000100",
			3010 => "0000000010111100110101",
			3011 => "0011111010110100000100",
			3012 => "0000001010111100110101",
			3013 => "0000000010111100110101",
			3014 => "0010010011101000000100",
			3015 => "1111111010111100110101",
			3016 => "0001100100101100001000",
			3017 => "0011001000011000000100",
			3018 => "0000000010111100110101",
			3019 => "0000001010111100110101",
			3020 => "0000000010111100110101",
			3021 => "0000001011000101000000",
			3022 => "0001000111011100110000",
			3023 => "0001110001011000010000",
			3024 => "0010000101000100000100",
			3025 => "0000000010111111001001",
			3026 => "0010010111110100001000",
			3027 => "0011001111011100000100",
			3028 => "0000000010111111001001",
			3029 => "0000000010111111001001",
			3030 => "0000000010111111001001",
			3031 => "0011000111010000010000",
			3032 => "0010010000001000000100",
			3033 => "0000000010111111001001",
			3034 => "0001110101110100001000",
			3035 => "0001110101100100000100",
			3036 => "0000000010111111001001",
			3037 => "0000000010111111001001",
			3038 => "0000000010111111001001",
			3039 => "0010101001000100000100",
			3040 => "0000000010111111001001",
			3041 => "0001000011110000000100",
			3042 => "0000000010111111001001",
			3043 => "0000100101010100000100",
			3044 => "0000000010111111001001",
			3045 => "0000000010111111001001",
			3046 => "0010000001110100001100",
			3047 => "0000000011010000000100",
			3048 => "0000000010111111001001",
			3049 => "0010010100111100000100",
			3050 => "0000000010111111001001",
			3051 => "0000000010111111001001",
			3052 => "0000000010111111001001",
			3053 => "0000000000101000001000",
			3054 => "0001001001000000000100",
			3055 => "0000000010111111001001",
			3056 => "0000010010111111001001",
			3057 => "0000000010111111001001",
			3058 => "0000011100011000110100",
			3059 => "0010011010100100101100",
			3060 => "0010011010100100100000",
			3061 => "0000010101011100000100",
			3062 => "1111111011000001101101",
			3063 => "0011001001110100001100",
			3064 => "0010011000010000000100",
			3065 => "0000000011000001101101",
			3066 => "0010011001111100000100",
			3067 => "1111111011000001101101",
			3068 => "1111111011000001101101",
			3069 => "0011101011101100001000",
			3070 => "0010010100101100000100",
			3071 => "1111111011000001101101",
			3072 => "0000010011000001101101",
			3073 => "0010011010100000000100",
			3074 => "1111111011000001101101",
			3075 => "0000000011000001101101",
			3076 => "0011000001101000001000",
			3077 => "0001011001010000000100",
			3078 => "1111111011000001101101",
			3079 => "0000000011000001101101",
			3080 => "0000010011000001101101",
			3081 => "0001101000010000000100",
			3082 => "0000010011000001101101",
			3083 => "1111111011000001101101",
			3084 => "0011011100010100001000",
			3085 => "0001001101001000000100",
			3086 => "1111111011000001101101",
			3087 => "0000000011000001101101",
			3088 => "0010100110011100010000",
			3089 => "0011001001110100000100",
			3090 => "0000001011000001101101",
			3091 => "0001110111010000000100",
			3092 => "0000001011000001101101",
			3093 => "0011001011011100000100",
			3094 => "0000010011000001101101",
			3095 => "0000010011000001101101",
			3096 => "0001110101110100000100",
			3097 => "1111111011000001101101",
			3098 => "0000000011000001101101",
			3099 => "0000011100011000101100",
			3100 => "0000010101011100001100",
			3101 => "0000011001011000000100",
			3102 => "1111111011000100110001",
			3103 => "0000011001011000000100",
			3104 => "0000000011000100110001",
			3105 => "1111111011000100110001",
			3106 => "0001000100001100010100",
			3107 => "0001110000011100001000",
			3108 => "0001011110010000000100",
			3109 => "1111111011000100110001",
			3110 => "0000000011000100110001",
			3111 => "0001101000010000001000",
			3112 => "0000011101111100000100",
			3113 => "1111111011000100110001",
			3114 => "0000001011000100110001",
			3115 => "1111111011000100110001",
			3116 => "0000100110001100000100",
			3117 => "0000001011000100110001",
			3118 => "0001100101010000000100",
			3119 => "0000001011000100110001",
			3120 => "1111111011000100110001",
			3121 => "0011001001110100001100",
			3122 => "0001100101010000001000",
			3123 => "0011111011110000000100",
			3124 => "1111111011000100110001",
			3125 => "0000000011000100110001",
			3126 => "1111111011000100110001",
			3127 => "0001100100101100100100",
			3128 => "0010110001001000001100",
			3129 => "0011001000011000001000",
			3130 => "0010000001110000000100",
			3131 => "0000001011000100110001",
			3132 => "1111111011000100110001",
			3133 => "0000001011000100110001",
			3134 => "0001101001111100010000",
			3135 => "0011011010000100001000",
			3136 => "0010110000110100000100",
			3137 => "0000001011000100110001",
			3138 => "0000001011000100110001",
			3139 => "0011011010000100000100",
			3140 => "0000000011000100110001",
			3141 => "0000001011000100110001",
			3142 => "0000011011001100000100",
			3143 => "0000000011000100110001",
			3144 => "0000001011000100110001",
			3145 => "0000000000110000000100",
			3146 => "1111111011000100110001",
			3147 => "0000000011000100110001",
			3148 => "0001001001000000111100",
			3149 => "0010000110001000110100",
			3150 => "0001000011110000100000",
			3151 => "0010000001010100010000",
			3152 => "0001110111010000000100",
			3153 => "0000000011000111000101",
			3154 => "0000111100001100001000",
			3155 => "0000010100110100000100",
			3156 => "0000000011000111000101",
			3157 => "0000000011000111000101",
			3158 => "0000000011000111000101",
			3159 => "0011000111010000001100",
			3160 => "0001110101110100001000",
			3161 => "0010010011101000000100",
			3162 => "0000000011000111000101",
			3163 => "0000000011000111000101",
			3164 => "0000000011000111000101",
			3165 => "0000000011000111000101",
			3166 => "0011001001110100000100",
			3167 => "0000000011000111000101",
			3168 => "0011001011011100001100",
			3169 => "0011101101001000001000",
			3170 => "0000010111101000000100",
			3171 => "0000000011000111000101",
			3172 => "0000000011000111000101",
			3173 => "0000000011000111000101",
			3174 => "0000000011000111000101",
			3175 => "0000100101010100000100",
			3176 => "0000000011000111000101",
			3177 => "0000000011000111000101",
			3178 => "0010000001110100001100",
			3179 => "0000000011010000000100",
			3180 => "0000000011000111000101",
			3181 => "0000010101011100000100",
			3182 => "0000000011000111000101",
			3183 => "0000000011000111000101",
			3184 => "0000000011000111000101",
			3185 => "0000100010010100001100",
			3186 => "0010000101000100000100",
			3187 => "0000000011001001111001",
			3188 => "0001010111111100000100",
			3189 => "1111111011001001111001",
			3190 => "0000000011001001111001",
			3191 => "0011100110111000100000",
			3192 => "0000010111101000010000",
			3193 => "0000101110000000001100",
			3194 => "0001000111011100000100",
			3195 => "0000000011001001111001",
			3196 => "0001101111000000000100",
			3197 => "0000000011001001111001",
			3198 => "0000000011001001111001",
			3199 => "0000000011001001111001",
			3200 => "0011000111010000001100",
			3201 => "0011011001011100000100",
			3202 => "0000000011001001111001",
			3203 => "0011001001110100000100",
			3204 => "0000000011001001111001",
			3205 => "0000000011001001111001",
			3206 => "0000000011001001111001",
			3207 => "0001110110110100010100",
			3208 => "0000011101011000001100",
			3209 => "0010111110101100001000",
			3210 => "0000001010101100000100",
			3211 => "0000000011001001111001",
			3212 => "1111111011001001111001",
			3213 => "0000000011001001111001",
			3214 => "0010001011010100000100",
			3215 => "0000000011001001111001",
			3216 => "0000000011001001111001",
			3217 => "0000110011110000001100",
			3218 => "0001001110100100000100",
			3219 => "0000000011001001111001",
			3220 => "0000010100110100000100",
			3221 => "0000000011001001111001",
			3222 => "0000000011001001111001",
			3223 => "0000011001100100001100",
			3224 => "0010101001000100000100",
			3225 => "0000000011001001111001",
			3226 => "0011000111010000000100",
			3227 => "0000000011001001111001",
			3228 => "0000000011001001111001",
			3229 => "0000000011001001111001",
			3230 => "0000011100011000101000",
			3231 => "0000010101011100000100",
			3232 => "1111111011001100100101",
			3233 => "0001000100001100010100",
			3234 => "0001110000011100001000",
			3235 => "0001011110010000000100",
			3236 => "1111111011001100100101",
			3237 => "0000000011001100100101",
			3238 => "0010011010100000000100",
			3239 => "1111111011001100100101",
			3240 => "0001010011001000000100",
			3241 => "0000001011001100100101",
			3242 => "0000000011001100100101",
			3243 => "0001011100010100001100",
			3244 => "0010000001110100001000",
			3245 => "0010110101110100000100",
			3246 => "0000010011001100100101",
			3247 => "0000001011001100100101",
			3248 => "0000000011001100100101",
			3249 => "1111111011001100100101",
			3250 => "0011001001110100001100",
			3251 => "0010101001000100001000",
			3252 => "0001001100001100000100",
			3253 => "1111111011001100100101",
			3254 => "0000001011001100100101",
			3255 => "1111111011001100100101",
			3256 => "0010000001110100100000",
			3257 => "0000011100011000001100",
			3258 => "0010101000010100000100",
			3259 => "0000001011001100100101",
			3260 => "0011100110111000000100",
			3261 => "0000001011001100100101",
			3262 => "1111111011001100100101",
			3263 => "0011010110111100000100",
			3264 => "0000001011001100100101",
			3265 => "0000000111000000001000",
			3266 => "0011111000011100000100",
			3267 => "0000001011001100100101",
			3268 => "1111111011001100100101",
			3269 => "0010101010110000000100",
			3270 => "0000001011001100100101",
			3271 => "0000000011001100100101",
			3272 => "1111111011001100100101",
			3273 => "0000010101011100000100",
			3274 => "1111111011001110101001",
			3275 => "0000100011110000110100",
			3276 => "0001010110010000011100",
			3277 => "0010011010100100010100",
			3278 => "0001000100001100001100",
			3279 => "0010000001010100000100",
			3280 => "0000000011001110101001",
			3281 => "0001111011011100000100",
			3282 => "0000000011001110101001",
			3283 => "0000000011001110101001",
			3284 => "0001110111010000000100",
			3285 => "0000000011001110101001",
			3286 => "0000000011001110101001",
			3287 => "0011011100010100000100",
			3288 => "0000000011001110101001",
			3289 => "0000001011001110101001",
			3290 => "0011001010001100010000",
			3291 => "0010010011101000000100",
			3292 => "0000000011001110101001",
			3293 => "0010101000010100001000",
			3294 => "0011010110111100000100",
			3295 => "0000000011001110101001",
			3296 => "1111111011001110101001",
			3297 => "0000000011001110101001",
			3298 => "0000001000110000000100",
			3299 => "0000000011001110101001",
			3300 => "0000000011001110101001",
			3301 => "0010001100000100000100",
			3302 => "0000000011001110101001",
			3303 => "0000011011001100000100",
			3304 => "0000000011001110101001",
			3305 => "0000000011001110101001",
			3306 => "0000101100111000000100",
			3307 => "1111111011010000100101",
			3308 => "0001001011001000110000",
			3309 => "0010101100011100100100",
			3310 => "0000011101011000011100",
			3311 => "0000001010101100001100",
			3312 => "0001110111010000000100",
			3313 => "0000000011010000100101",
			3314 => "0000010100110100000100",
			3315 => "0000000011010000100101",
			3316 => "0000001011010000100101",
			3317 => "0001000011110000001000",
			3318 => "0001110110110100000100",
			3319 => "0000000011010000100101",
			3320 => "0000000011010000100101",
			3321 => "0010100110011000000100",
			3322 => "0000000011010000100101",
			3323 => "0000000011010000100101",
			3324 => "0011011001100000000100",
			3325 => "0000000011010000100101",
			3326 => "0000001011010000100101",
			3327 => "0000100010010100000100",
			3328 => "0000000011010000100101",
			3329 => "0010000110001000000100",
			3330 => "0000000011010000100101",
			3331 => "0000000011010000100101",
			3332 => "0010100101000100001000",
			3333 => "0000111110010000000100",
			3334 => "0000000011010000100101",
			3335 => "0000001011010000100101",
			3336 => "0000000011010000100101",
			3337 => "0010011010100100100100",
			3338 => "0001100100111100000100",
			3339 => "1111111011010100000001",
			3340 => "0001101000010000001100",
			3341 => "0001001110111000000100",
			3342 => "1111111011010100000001",
			3343 => "0011001010111000000100",
			3344 => "0000000011010100000001",
			3345 => "0000001011010100000001",
			3346 => "0010010100101100000100",
			3347 => "1111111011010100000001",
			3348 => "0001000011101100001100",
			3349 => "0010010111101100001000",
			3350 => "0010010111101100000100",
			3351 => "0000000011010100000001",
			3352 => "0000000011010100000001",
			3353 => "1111111011010100000001",
			3354 => "0000001011010100000001",
			3355 => "0010110000110100100100",
			3356 => "0011100110111000010100",
			3357 => "0001001000001000010000",
			3358 => "0001010111111100001000",
			3359 => "0001100100111100000100",
			3360 => "0000000011010100000001",
			3361 => "1111111011010100000001",
			3362 => "0010011010100100000100",
			3363 => "0000000011010100000001",
			3364 => "0000001011010100000001",
			3365 => "0000001011010100000001",
			3366 => "0011100110111000000100",
			3367 => "1111010011010100000001",
			3368 => "0011001000011000001000",
			3369 => "0010010011101000000100",
			3370 => "1111111011010100000001",
			3371 => "0000000011010100000001",
			3372 => "0000001011010100000001",
			3373 => "0011010110111100010000",
			3374 => "0011000001011000001000",
			3375 => "0011100011110000000100",
			3376 => "0000001011010100000001",
			3377 => "0000000011010100000001",
			3378 => "0010110110100000000100",
			3379 => "0000000011010100000001",
			3380 => "0000000011010100000001",
			3381 => "0001110110110100001000",
			3382 => "0010101000010100000100",
			3383 => "1111101011010100000001",
			3384 => "0000000011010100000001",
			3385 => "0001100100101100001100",
			3386 => "0011101000000100001000",
			3387 => "0001110101110100000100",
			3388 => "0000001011010100000001",
			3389 => "1111111011010100000001",
			3390 => "0000001011010100000001",
			3391 => "1111111011010100000001",
			3392 => "0011001000000000001100",
			3393 => "0000100110111000000100",
			3394 => "1111111011010110111101",
			3395 => "0000100110111000000100",
			3396 => "0000000011010110111101",
			3397 => "1111111011010110111101",
			3398 => "0000011101011001000000",
			3399 => "0000111110100100100100",
			3400 => "0010011001111100001100",
			3401 => "0011001000000000001000",
			3402 => "0000010101011100000100",
			3403 => "0000000011010110111101",
			3404 => "0000000011010110111101",
			3405 => "1111111011010110111101",
			3406 => "0001100100111100001000",
			3407 => "0011111000101000000100",
			3408 => "0000000011010110111101",
			3409 => "0000001011010110111101",
			3410 => "0001001010110100001000",
			3411 => "0000011100011000000100",
			3412 => "1111111011010110111101",
			3413 => "0000000011010110111101",
			3414 => "0001101001111100000100",
			3415 => "0000001011010110111101",
			3416 => "0000000011010110111101",
			3417 => "0001110110110100010000",
			3418 => "0010010010101100001000",
			3419 => "0001100101010000000100",
			3420 => "0000000011010110111101",
			3421 => "0000000011010110111101",
			3422 => "0010010011101000000100",
			3423 => "1111111011010110111101",
			3424 => "1111110011010110111101",
			3425 => "0010101010110000001000",
			3426 => "0000010100110100000100",
			3427 => "0000000011010110111101",
			3428 => "0000001011010110111101",
			3429 => "1111111011010110111101",
			3430 => "0010101000010100001000",
			3431 => "0010010011101000000100",
			3432 => "0000001011010110111101",
			3433 => "1111111011010110111101",
			3434 => "0001100100101100001000",
			3435 => "0011011110110100000100",
			3436 => "0000000011010110111101",
			3437 => "0000001011010110111101",
			3438 => "0000000011010110111101",
			3439 => "0010010100111100000100",
			3440 => "1111111011011001011001",
			3441 => "0001100101010000110000",
			3442 => "0001000011110000100000",
			3443 => "0001010111111100000100",
			3444 => "1111111011011001011001",
			3445 => "0011111000110100001100",
			3446 => "0000010100110100000100",
			3447 => "0000000011011001011001",
			3448 => "0010000001110000000100",
			3449 => "0000001011011001011001",
			3450 => "0000000011011001011001",
			3451 => "0010101000010100001000",
			3452 => "0001101000010000000100",
			3453 => "0000000011011001011001",
			3454 => "1111111011011001011001",
			3455 => "0001010011001000000100",
			3456 => "0000000011011001011001",
			3457 => "0000000011011001011001",
			3458 => "0000100010110000001000",
			3459 => "0000100110111000000100",
			3460 => "0000000011011001011001",
			3461 => "0000001011011001011001",
			3462 => "0000011011001100000100",
			3463 => "0000000011011001011001",
			3464 => "0000000011011001011001",
			3465 => "0001000100001100001100",
			3466 => "0010011000100100001000",
			3467 => "0010100110011000000100",
			3468 => "0000000011011001011001",
			3469 => "1111111011011001011001",
			3470 => "0000000011011001011001",
			3471 => "0010000111000100001000",
			3472 => "0000010100110100000100",
			3473 => "0000000011011001011001",
			3474 => "0000000011011001011001",
			3475 => "0001101001111100000100",
			3476 => "0000000011011001011001",
			3477 => "1111111011011001011001",
			3478 => "0011001010111000000100",
			3479 => "0000000011011011100101",
			3480 => "0001000011010100110000",
			3481 => "0001100100111100001100",
			3482 => "0000010100110100000100",
			3483 => "0000000011011011100101",
			3484 => "0010110100010000000100",
			3485 => "0000000011011011100101",
			3486 => "0000000011011011100101",
			3487 => "0000011100011000001000",
			3488 => "0011110010010100000100",
			3489 => "0000000011011011100101",
			3490 => "0000000011011011100101",
			3491 => "0010000001010100010000",
			3492 => "0010110110100000001000",
			3493 => "0010000101000100000100",
			3494 => "0000000011011011100101",
			3495 => "0000000011011011100101",
			3496 => "0010000001010100000100",
			3497 => "0000000011011011100101",
			3498 => "0000000011011011100101",
			3499 => "0000100010110000001000",
			3500 => "0001010111111100000100",
			3501 => "0000000011011011100101",
			3502 => "0000000011011011100101",
			3503 => "0000000011011011100101",
			3504 => "0010100101000100010000",
			3505 => "0000010101011100000100",
			3506 => "0000000011011011100101",
			3507 => "0011011001100000000100",
			3508 => "0000000011011011100101",
			3509 => "0011011010000100000100",
			3510 => "0000000011011011100101",
			3511 => "0000000011011011100101",
			3512 => "0000000011011011100101",
			3513 => "0010011010100100101000",
			3514 => "0000101101101100000100",
			3515 => "1111111011011110100001",
			3516 => "0001100101010000100000",
			3517 => "0001001110111000001100",
			3518 => "0011001000011000000100",
			3519 => "1111111011011110100001",
			3520 => "0001110001011000000100",
			3521 => "0000000011011110100001",
			3522 => "1111111011011110100001",
			3523 => "0010011011001100000100",
			3524 => "1111111011011110100001",
			3525 => "0000100101000000001000",
			3526 => "0001111011000000000100",
			3527 => "0000000011011110100001",
			3528 => "0000010011011110100001",
			3529 => "0000010111101000000100",
			3530 => "1111111011011110100001",
			3531 => "0000001011011110100001",
			3532 => "1111111011011110100001",
			3533 => "0011001001110100001000",
			3534 => "0001010111111100000100",
			3535 => "1111111011011110100001",
			3536 => "0000000011011110100001",
			3537 => "0010001001101000011100",
			3538 => "0011011010000100010100",
			3539 => "0010110001001000001000",
			3540 => "0000011100011000000100",
			3541 => "0000000011011110100001",
			3542 => "0000001011011110100001",
			3543 => "0011010110111100000100",
			3544 => "0000001011011110100001",
			3545 => "0010111110101100000100",
			3546 => "0000000011011110100001",
			3547 => "0000001011011110100001",
			3548 => "0001000010110000000100",
			3549 => "1111111011011110100001",
			3550 => "0000001011011110100001",
			3551 => "0001000000010100001000",
			3552 => "0000011011001100000100",
			3553 => "1111111011011110100001",
			3554 => "0000000011011110100001",
			3555 => "0010000111000100001000",
			3556 => "0010001011010100000100",
			3557 => "0000000011011110100001",
			3558 => "0000001011011110100001",
			3559 => "1111111011011110100001",
			3560 => "0010011010100100100100",
			3561 => "0000101101101100000100",
			3562 => "1111111011100001010101",
			3563 => "0001100101010000011100",
			3564 => "0001001110111000001100",
			3565 => "0011001000011000000100",
			3566 => "1111111011100001010101",
			3567 => "0001110001011000000100",
			3568 => "0000000011100001010101",
			3569 => "1111111011100001010101",
			3570 => "0010011011001100000100",
			3571 => "1111111011100001010101",
			3572 => "0000111100010100000100",
			3573 => "0000101011100001010101",
			3574 => "0000100011110000000100",
			3575 => "0000001011100001010101",
			3576 => "0000000011100001010101",
			3577 => "1111111011100001010101",
			3578 => "0001010111111100001000",
			3579 => "0011001001110100000100",
			3580 => "1111111011100001010101",
			3581 => "0000000011100001010101",
			3582 => "0001101001111100100100",
			3583 => "0011110010111000011100",
			3584 => "0010110110100000001100",
			3585 => "0001001110111000001000",
			3586 => "0010011010100100000100",
			3587 => "0000000011100001010101",
			3588 => "0000001011100001010101",
			3589 => "0000001011100001010101",
			3590 => "0000000111000000001000",
			3591 => "0010010011101000000100",
			3592 => "0000001011100001010101",
			3593 => "1111111011100001010101",
			3594 => "0011010111011000000100",
			3595 => "0000000011100001010101",
			3596 => "0000001011100001010101",
			3597 => "0001010110010000000100",
			3598 => "1111111011100001010101",
			3599 => "0000001011100001010101",
			3600 => "0000011001100100000100",
			3601 => "1111111011100001010101",
			3602 => "0001100100101100000100",
			3603 => "0000001011100001010101",
			3604 => "0000000011100001010101",
			3605 => "0011001000000000001100",
			3606 => "0001001100111100000100",
			3607 => "1111111011100100101001",
			3608 => "0001000000101100000100",
			3609 => "0000000011100100101001",
			3610 => "0000000011100100101001",
			3611 => "0010110110100000111100",
			3612 => "0011001000011000100100",
			3613 => "0001111111011100001100",
			3614 => "0001001000001000000100",
			3615 => "0000000011100100101001",
			3616 => "0011111000011100000100",
			3617 => "0000001011100100101001",
			3618 => "0000000011100100101001",
			3619 => "0001110101100100001100",
			3620 => "0011001000000000000100",
			3621 => "0000000011100100101001",
			3622 => "0010000101000100000100",
			3623 => "0000000011100100101001",
			3624 => "1111111011100100101001",
			3625 => "0010110001001000000100",
			3626 => "0000000011100100101001",
			3627 => "0001100101010000000100",
			3628 => "0000000011100100101001",
			3629 => "0000000011100100101001",
			3630 => "0010011010100100001000",
			3631 => "0011001000011000000100",
			3632 => "0000000011100100101001",
			3633 => "0000000011100100101001",
			3634 => "0011101000011100000100",
			3635 => "0000001011100100101001",
			3636 => "0000110110001100000100",
			3637 => "0000000011100100101001",
			3638 => "0011111010110100000100",
			3639 => "0000000011100100101001",
			3640 => "0000000011100100101001",
			3641 => "0011000111010000010000",
			3642 => "0000111100001100000100",
			3643 => "0000000011100100101001",
			3644 => "0010111101000100001000",
			3645 => "0000101100001100000100",
			3646 => "1111111011100100101001",
			3647 => "0000000011100100101001",
			3648 => "0000000011100100101001",
			3649 => "0011101110000000001000",
			3650 => "0001110100010000000100",
			3651 => "0000000011100100101001",
			3652 => "1111111011100100101001",
			3653 => "0001100100101100001000",
			3654 => "0010010010101100000100",
			3655 => "0000000011100100101001",
			3656 => "0000001011100100101001",
			3657 => "0000000011100100101001",
			3658 => "0000010100110100011100",
			3659 => "0001100100111100000100",
			3660 => "1111111011100111010101",
			3661 => "0000110010010100010000",
			3662 => "0001000100001100000100",
			3663 => "1111111011100111010101",
			3664 => "0001110111010000001000",
			3665 => "0011001010111000000100",
			3666 => "1111111011100111010101",
			3667 => "0000001011100111010101",
			3668 => "0000000011100111010101",
			3669 => "0001101000010000000100",
			3670 => "0000000011100111010101",
			3671 => "1111111011100111010101",
			3672 => "0011001001110100000100",
			3673 => "1111111011100111010101",
			3674 => "0001100100111100001000",
			3675 => "0000001000101100000100",
			3676 => "0000001011100111010101",
			3677 => "0000010011100111010101",
			3678 => "0000011010011000011000",
			3679 => "0001111011011100010000",
			3680 => "0001000011110000001000",
			3681 => "0010110000110100000100",
			3682 => "1111111011100111010101",
			3683 => "0000000011100111010101",
			3684 => "0011101000110100000100",
			3685 => "0000001011100111010101",
			3686 => "1111111011100111010101",
			3687 => "0001101000010000000100",
			3688 => "0000001011100111010101",
			3689 => "1111111011100111010101",
			3690 => "0010110110100000001100",
			3691 => "0011100010111000001000",
			3692 => "0011011001100000000100",
			3693 => "0000000011100111010101",
			3694 => "0000001011100111010101",
			3695 => "0000000011100111010101",
			3696 => "0010101000010100000100",
			3697 => "1111111011100111010101",
			3698 => "0001100100101100000100",
			3699 => "0000001011100111010101",
			3700 => "0000000011100111010101",
			3701 => "0000100011000000001000",
			3702 => "0001011110010000000100",
			3703 => "1111111011101010100001",
			3704 => "0000000011101010100001",
			3705 => "0000111100001100111000",
			3706 => "0000011100011000100100",
			3707 => "0011111011110000010100",
			3708 => "0001111111011100001100",
			3709 => "0001001000001000000100",
			3710 => "0000000011101010100001",
			3711 => "0000010101011100000100",
			3712 => "0000000011101010100001",
			3713 => "0000000011101010100001",
			3714 => "0001010111111100000100",
			3715 => "0000000011101010100001",
			3716 => "0000000011101010100001",
			3717 => "0000111000000100001100",
			3718 => "0001001011100000001000",
			3719 => "0000100110111000000100",
			3720 => "0000000011101010100001",
			3721 => "0000000011101010100001",
			3722 => "0000000011101010100001",
			3723 => "0000000011101010100001",
			3724 => "0001110101110100001100",
			3725 => "0011110110001100001000",
			3726 => "0011011100010100000100",
			3727 => "0000000011101010100001",
			3728 => "0000001011101010100001",
			3729 => "0000000011101010100001",
			3730 => "0001010010000000000100",
			3731 => "0000000011101010100001",
			3732 => "0000000011101010100001",
			3733 => "0000000111000000001100",
			3734 => "0010010010101100000100",
			3735 => "0000000011101010100001",
			3736 => "0011010110111100000100",
			3737 => "0000000011101010100001",
			3738 => "1111111011101010100001",
			3739 => "0001001001001100001000",
			3740 => "0000011100011000000100",
			3741 => "0000000011101010100001",
			3742 => "0000000011101010100001",
			3743 => "0010011000100100001000",
			3744 => "0011101110100100000100",
			3745 => "0000000011101010100001",
			3746 => "1111111011101010100001",
			3747 => "0010000111000100001000",
			3748 => "0011001111011100000100",
			3749 => "0000000011101010100001",
			3750 => "0000000011101010100001",
			3751 => "0000000011101010100001",
			3752 => "0011001000000000010000",
			3753 => "0001001100111100000100",
			3754 => "1111111011101101110101",
			3755 => "0001000000101100001000",
			3756 => "0001101001100100000100",
			3757 => "0000000011101101110101",
			3758 => "0000000011101101110101",
			3759 => "0000000011101101110101",
			3760 => "0010110110100001000000",
			3761 => "0011001000011000100100",
			3762 => "0000100010110000100000",
			3763 => "0001000011110000010000",
			3764 => "0001010111111100001000",
			3765 => "0001101111000000000100",
			3766 => "0000000011101101110101",
			3767 => "1111111011101101110101",
			3768 => "0010101001000100000100",
			3769 => "0000000011101101110101",
			3770 => "0000000011101101110101",
			3771 => "0001101000010000001000",
			3772 => "0000101100001100000100",
			3773 => "0000001011101101110101",
			3774 => "0000000011101101110101",
			3775 => "0000011101111100000100",
			3776 => "0000000011101101110101",
			3777 => "0000000011101101110101",
			3778 => "1111111011101101110101",
			3779 => "0000011101111100001000",
			3780 => "0011001000011000000100",
			3781 => "0000000011101101110101",
			3782 => "0000000011101101110101",
			3783 => "0011101000011100001000",
			3784 => "0011011111010100000100",
			3785 => "0000001011101101110101",
			3786 => "0000000011101101110101",
			3787 => "0000110110001100000100",
			3788 => "0000000011101101110101",
			3789 => "0011111010110100000100",
			3790 => "0000000011101101110101",
			3791 => "0000000011101101110101",
			3792 => "0000011101011000010000",
			3793 => "0001101000010000000100",
			3794 => "0000000011101101110101",
			3795 => "0011101110100100001000",
			3796 => "0001010010000100000100",
			3797 => "1111111011101101110101",
			3798 => "0000000011101101110101",
			3799 => "0000000011101101110101",
			3800 => "0001100100101100001000",
			3801 => "0011001010001100000100",
			3802 => "0000000011101101110101",
			3803 => "0000001011101101110101",
			3804 => "0000000011101101110101",
			3805 => "0010011010100000101000",
			3806 => "0001100100111100000100",
			3807 => "1111111011110001101001",
			3808 => "0011110110111000011000",
			3809 => "0011001010111000000100",
			3810 => "1111111011110001101001",
			3811 => "0011111111101000001000",
			3812 => "0010100110011000000100",
			3813 => "0000000011110001101001",
			3814 => "0000001011110001101001",
			3815 => "0011110110111000001000",
			3816 => "0001101000010000000100",
			3817 => "0000000011110001101001",
			3818 => "0000000011110001101001",
			3819 => "0000000011110001101001",
			3820 => "0011011100010100001000",
			3821 => "0011011010001000000100",
			3822 => "1111111011110001101001",
			3823 => "0000000011110001101001",
			3824 => "1111111011110001101001",
			3825 => "0000011100011000101100",
			3826 => "0011100010010100011000",
			3827 => "0000110001011100001000",
			3828 => "0010001001101000000100",
			3829 => "1111111011110001101001",
			3830 => "0000000011110001101001",
			3831 => "0001110100010000001100",
			3832 => "0000101011110000001000",
			3833 => "0001110111010000000100",
			3834 => "1111111011110001101001",
			3835 => "0000001011110001101001",
			3836 => "0000001011110001101001",
			3837 => "0000000011110001101001",
			3838 => "0010101000010100000100",
			3839 => "0000001011110001101001",
			3840 => "0010011010100100001100",
			3841 => "0010011010100100000100",
			3842 => "1111111011110001101001",
			3843 => "0000100110001100000100",
			3844 => "0000000011110001101001",
			3845 => "0000000011110001101001",
			3846 => "1111111011110001101001",
			3847 => "0010000110001000100000",
			3848 => "0011011010000100011000",
			3849 => "0001110111010000001100",
			3850 => "0011100110111000001000",
			3851 => "0000101011110000000100",
			3852 => "0000000011110001101001",
			3853 => "0000001011110001101001",
			3854 => "1111111011110001101001",
			3855 => "0001110111110000001000",
			3856 => "0011000100000100000100",
			3857 => "0000001011110001101001",
			3858 => "0000000011110001101001",
			3859 => "0000000011110001101001",
			3860 => "0000100101000000000100",
			3861 => "1111111011110001101001",
			3862 => "0000001011110001101001",
			3863 => "0001110010001000000100",
			3864 => "1111111011110001101001",
			3865 => "0000000011110001101001",
			3866 => "0011000100011000000100",
			3867 => "1111111011110100001101",
			3868 => "0000011010011000111100",
			3869 => "0001000000010100101100",
			3870 => "0010110000110100011000",
			3871 => "0011100110111000010000",
			3872 => "0011000001101000001000",
			3873 => "0001000011001100000100",
			3874 => "1111111011110100001101",
			3875 => "0000000011110100001101",
			3876 => "0011011100010100000100",
			3877 => "0000000011110100001101",
			3878 => "0000000011110100001101",
			3879 => "0011001111011100000100",
			3880 => "1111111011110100001101",
			3881 => "0000000011110100001101",
			3882 => "0011000100000100001000",
			3883 => "0010011010100100000100",
			3884 => "0000000011110100001101",
			3885 => "0000001011110100001101",
			3886 => "0011101000110100001000",
			3887 => "0001000110001100000100",
			3888 => "0000000011110100001101",
			3889 => "1111111011110100001101",
			3890 => "0000000011110100001101",
			3891 => "0001101001111100001100",
			3892 => "0011011100010000001000",
			3893 => "0010011011001100000100",
			3894 => "0000000011110100001101",
			3895 => "0000001011110100001101",
			3896 => "0000000011110100001101",
			3897 => "1111111011110100001101",
			3898 => "0000110101000000000100",
			3899 => "0000001011110100001101",
			3900 => "0000000111000000000100",
			3901 => "1111111011110100001101",
			3902 => "0010000111000100001000",
			3903 => "0011000001101000000100",
			3904 => "0000000011110100001101",
			3905 => "0000001011110100001101",
			3906 => "0000000011110100001101",
			3907 => "0010010100111100000100",
			3908 => "1111111011110111001001",
			3909 => "0000111110100100101100",
			3910 => "0000100011000000001000",
			3911 => "0010110001001000000100",
			3912 => "1111111011110111001001",
			3913 => "0000000011110111001001",
			3914 => "0000011100011000011100",
			3915 => "0011101000101000010000",
			3916 => "0000010111101000001000",
			3917 => "0011111111101000000100",
			3918 => "0000000011110111001001",
			3919 => "0000000011110111001001",
			3920 => "0001110110110100000100",
			3921 => "0000001011110111001001",
			3922 => "0000000011110111001001",
			3923 => "0001001110111000001000",
			3924 => "0001100100111100000100",
			3925 => "0000000011110111001001",
			3926 => "1111111011110111001001",
			3927 => "0000000011110111001001",
			3928 => "0011001001110100000100",
			3929 => "0000000011110111001001",
			3930 => "0000001011110111001001",
			3931 => "0001110110110100010100",
			3932 => "0000011101011000001000",
			3933 => "0010010010101100000100",
			3934 => "0000000011110111001001",
			3935 => "1111111011110111001001",
			3936 => "0011100110001100000100",
			3937 => "0000000011110111001001",
			3938 => "0010001001101000000100",
			3939 => "0000000011110111001001",
			3940 => "0000000011110111001001",
			3941 => "0001111011110100010100",
			3942 => "0010010010101100001100",
			3943 => "0001101001111100001000",
			3944 => "0010011010100100000100",
			3945 => "0000000011110111001001",
			3946 => "0000000011110111001001",
			3947 => "0000000011110111001001",
			3948 => "0001001100001100000100",
			3949 => "0000000011110111001001",
			3950 => "0000001011110111001001",
			3951 => "0011000100000100000100",
			3952 => "0000000011110111001001",
			3953 => "0000000011110111001001",
			3954 => "0011001000000000000100",
			3955 => "1111111011111010010101",
			3956 => "0010110110100001000100",
			3957 => "0011001000011000101000",
			3958 => "0001111111011100010000",
			3959 => "0001111000011000000100",
			3960 => "0000000011111010010101",
			3961 => "0000001000110000000100",
			3962 => "0000000011111010010101",
			3963 => "0011111000110100000100",
			3964 => "0000001011111010010101",
			3965 => "0000000011111010010101",
			3966 => "0001100101010000010000",
			3967 => "0010110001001000001000",
			3968 => "0000101000000100000100",
			3969 => "0000000011111010010101",
			3970 => "0000000011111010010101",
			3971 => "0000011101111100000100",
			3972 => "0000000011111010010101",
			3973 => "0000000011111010010101",
			3974 => "0000101110100100000100",
			3975 => "0000000011111010010101",
			3976 => "1111111011111010010101",
			3977 => "0000011101111100001000",
			3978 => "0011001000011000000100",
			3979 => "0000000011111010010101",
			3980 => "0000000011111010010101",
			3981 => "0011101000011100001000",
			3982 => "0011110011110000000100",
			3983 => "0000001011111010010101",
			3984 => "0000000011111010010101",
			3985 => "0000110110001100000100",
			3986 => "0000000011111010010101",
			3987 => "0011111010110100000100",
			3988 => "0000000011111010010101",
			3989 => "0000000011111010010101",
			3990 => "0000011101011000010000",
			3991 => "0001101000010000000100",
			3992 => "0000000011111010010101",
			3993 => "0011101110100100001000",
			3994 => "0001010010000100000100",
			3995 => "1111111011111010010101",
			3996 => "0000000011111010010101",
			3997 => "0000000011111010010101",
			3998 => "0001100100101100001100",
			3999 => "0001110100010000001000",
			4000 => "0011001010001100000100",
			4001 => "0000000011111010010101",
			4002 => "0000000011111010010101",
			4003 => "0000001011111010010101",
			4004 => "0000000011111010010101",
			4005 => "0010010100111100000100",
			4006 => "1111111011111101100011",
			4007 => "0001100101010001001100",
			4008 => "0000000111000000101000",
			4009 => "0001101000010000010100",
			4010 => "0001111011011100001100",
			4011 => "0000011010011000001000",
			4012 => "0010111110101100000100",
			4013 => "0000000011111101100011",
			4014 => "0000000011111101100011",
			4015 => "0000000011111101100011",
			4016 => "0000010100110100000100",
			4017 => "0000000011111101100011",
			4018 => "0000001011111101100011",
			4019 => "0010110110100000001100",
			4020 => "0000011100011000000100",
			4021 => "1111111011111101100011",
			4022 => "0000111110000000000100",
			4023 => "0000000011111101100011",
			4024 => "0000000011111101100011",
			4025 => "0011111000011100000100",
			4026 => "0000000011111101100011",
			4027 => "1111111011111101100011",
			4028 => "0000100010110000011100",
			4029 => "0011001011000000001100",
			4030 => "0011100010000000001000",
			4031 => "0000110110010000000100",
			4032 => "0000000011111101100011",
			4033 => "0000000011111101100011",
			4034 => "0000000011111101100011",
			4035 => "0000101110000000001000",
			4036 => "0000011100011000000100",
			4037 => "0000000011111101100011",
			4038 => "0000000011111101100011",
			4039 => "0001110001101000000100",
			4040 => "0000000011111101100011",
			4041 => "0000001011111101100011",
			4042 => "0000011011001100000100",
			4043 => "0000000011111101100011",
			4044 => "0000000011111101100011",
			4045 => "0000011101011000001100",
			4046 => "0000000000110000001000",
			4047 => "0001110111110000000100",
			4048 => "1111111011111101100011",
			4049 => "0000000011111101100011",
			4050 => "0000000011111101100011",
			4051 => "0010001111001000001000",
			4052 => "0000100101000000000100",
			4053 => "0000000011111101100011",
			4054 => "0000000011111101100011",
			4055 => "0000000011111101100011",
			4056 => "0000000011111101100101",
			4057 => "0001011111010100000100",
			4058 => "0000000011111101110001",
			4059 => "1111111011111101110001",
			4060 => "0011001011011100000100",
			4061 => "0000000011111101111101",
			4062 => "0000000011111101111101",
			4063 => "0001000011010100000100",
			4064 => "0000000011111110010001",
			4065 => "0001000001100100000100",
			4066 => "0000000011111110010001",
			4067 => "0000000011111110010001",
			4068 => "0010000110001000001000",
			4069 => "0010000001010100000100",
			4070 => "0000000011111110100101",
			4071 => "0000000011111110100101",
			4072 => "0000000011111110100101",
			4073 => "0001011111100100000100",
			4074 => "0000000011111110111001",
			4075 => "0011011000101000000100",
			4076 => "1111110011111110111001",
			4077 => "0000000011111110111001",
			4078 => "0001110001001000001100",
			4079 => "0001000100001100000100",
			4080 => "0000000011111111010101",
			4081 => "0001000001100100000100",
			4082 => "0000000011111111010101",
			4083 => "0000000011111111010101",
			4084 => "0000000011111111010101",
			4085 => "0001110001001000001100",
			4086 => "0001000000010100000100",
			4087 => "0000000011111111110001",
			4088 => "0001000001100100000100",
			4089 => "0000000011111111110001",
			4090 => "0000000011111111110001",
			4091 => "0000000011111111110001",
			4092 => "0001000100001100001100",
			4093 => "0001001110100100000100",
			4094 => "0000000100000000010101",
			4095 => "0001000000010100000100",
			4096 => "0000000100000000010101",
			4097 => "0000000100000000010101",
			4098 => "0001000001100100000100",
			4099 => "0000000100000000010101",
			4100 => "0000000100000000010101",
			4101 => "0000011100011000001100",
			4102 => "0010100110011100001000",
			4103 => "0010101000010100000100",
			4104 => "0000000100000000111001",
			4105 => "0000000100000000111001",
			4106 => "0000000100000000111001",
			4107 => "0010101010110000000100",
			4108 => "0000000100000000111001",
			4109 => "0000000100000000111001",
			4110 => "0011000111010000001100",
			4111 => "0011001010111000000100",
			4112 => "0000000100000001011101",
			4113 => "0010110110100000000100",
			4114 => "0000000100000001011101",
			4115 => "0000000100000001011101",
			4116 => "0001111011011100000100",
			4117 => "0000000100000001011101",
			4118 => "0000000100000001011101",
			4119 => "0001000100001100001100",
			4120 => "0001001100001100000100",
			4121 => "0000000100000010001001",
			4122 => "0010011000100100000100",
			4123 => "0000000100000010001001",
			4124 => "0000000100000010001001",
			4125 => "0010011001111100000100",
			4126 => "0000000100000010001001",
			4127 => "0001100100101100000100",
			4128 => "0000000100000010001001",
			4129 => "0000000100000010001001",
			4130 => "0010011010100100001100",
			4131 => "0001111000011000001000",
			4132 => "0011001010111000000100",
			4133 => "0000000100000010110101",
			4134 => "0000000100000010110101",
			4135 => "0000000100000010110101",
			4136 => "0011000001101000000100",
			4137 => "0000000100000010110101",
			4138 => "0001111011110100000100",
			4139 => "0000000100000010110101",
			4140 => "0000000100000010110101",
			4141 => "0011000111010000010000",
			4142 => "0011001010111000000100",
			4143 => "0000000100000011011001",
			4144 => "0011011010000100001000",
			4145 => "0011011110101100000100",
			4146 => "0000000100000011011001",
			4147 => "0000000100000011011001",
			4148 => "0000000100000011011001",
			4149 => "0000000100000011011001",
			4150 => "0011011100111000010000",
			4151 => "0011000100011000000100",
			4152 => "0000000100000011111101",
			4153 => "0001100100101100001000",
			4154 => "0001101001100100000100",
			4155 => "0000000100000011111101",
			4156 => "0000000100000011111101",
			4157 => "0000000100000011111101",
			4158 => "0000000100000011111101",
			4159 => "0011111110100100000100",
			4160 => "0000000100000100100001",
			4161 => "0000011111000000001100",
			4162 => "0010101000010100000100",
			4163 => "0000000100000100100001",
			4164 => "0000110011101100000100",
			4165 => "0000000100000100100001",
			4166 => "0000000100000100100001",
			4167 => "0000000100000100100001",
			4168 => "0010011010100100001000",
			4169 => "0010110101110100000100",
			4170 => "0000000100000101001101",
			4171 => "0000000100000101001101",
			4172 => "0011000001101000000100",
			4173 => "0000000100000101001101",
			4174 => "0010000111000100001000",
			4175 => "0000000111000000000100",
			4176 => "0000000100000101001101",
			4177 => "0000000100000101001101",
			4178 => "0000000100000101001101",
			4179 => "0001110001001000010100",
			4180 => "0001000000010100001000",
			4181 => "0000011101011000000100",
			4182 => "0000000100000101111001",
			4183 => "0000000100000101111001",
			4184 => "0010011001111100000100",
			4185 => "0000000100000101111001",
			4186 => "0001100100101100000100",
			4187 => "0000000100000101111001",
			4188 => "0000000100000101111001",
			4189 => "1111111100000101111001",
			4190 => "0001000000010100001100",
			4191 => "0001001110100100000100",
			4192 => "0000000100000110101101",
			4193 => "0011111010110100000100",
			4194 => "0000000100000110101101",
			4195 => "0000000100000110101101",
			4196 => "0001000001100100001100",
			4197 => "0000101101101100000100",
			4198 => "0000000100000110101101",
			4199 => "0000101110100100000100",
			4200 => "0000000100000110101101",
			4201 => "0000000100000110101101",
			4202 => "0000000100000110101101",
			4203 => "0010001111001000010000",
			4204 => "0001000000010100000100",
			4205 => "0000000100000111100001",
			4206 => "0001110001101000000100",
			4207 => "0000000100000111100001",
			4208 => "0000000010011000000100",
			4209 => "0000000100000111100001",
			4210 => "0000000100000111100001",
			4211 => "0001000000101100001000",
			4212 => "0010101100011100000100",
			4213 => "0000000100000111100001",
			4214 => "0000000100000111100001",
			4215 => "0000000100000111100001",
			4216 => "0010000110001000010100",
			4217 => "0001001110100100000100",
			4218 => "0000000100001000010101",
			4219 => "0011001001110100000100",
			4220 => "0000000100001000010101",
			4221 => "0001111011110100001000",
			4222 => "0000011110010100000100",
			4223 => "0000000100001000010101",
			4224 => "0000000100001000010101",
			4225 => "0000000100001000010101",
			4226 => "0001001001000000000100",
			4227 => "0000000100001000010101",
			4228 => "0000000100001000010101",
			4229 => "0010110110100000010100",
			4230 => "0010111010011100000100",
			4231 => "0000000100001001000001",
			4232 => "0000100010110000001100",
			4233 => "0000101100111000000100",
			4234 => "0000000100001001000001",
			4235 => "0000110101000000000100",
			4236 => "0000000100001001000001",
			4237 => "0000000100001001000001",
			4238 => "0000000100001001000001",
			4239 => "0000000100001001000001",
			4240 => "0010110101110100010000",
			4241 => "0011000100011000000100",
			4242 => "0000000100001010000101",
			4243 => "0001000100001100000100",
			4244 => "0000000100001010000101",
			4245 => "0010000111000000000100",
			4246 => "0000001100001010000101",
			4247 => "0000000100001010000101",
			4248 => "0010000110001000001100",
			4249 => "0011000001101000000100",
			4250 => "0000000100001010000101",
			4251 => "0011000100000100000100",
			4252 => "0000000100001010000101",
			4253 => "0000000100001010000101",
			4254 => "0011100011010100000100",
			4255 => "0000000100001010000101",
			4256 => "0000000100001010000101",
			4257 => "0001111011110100010100",
			4258 => "0010011001111100000100",
			4259 => "0000000100001011000001",
			4260 => "0000100110111000000100",
			4261 => "0000000100001011000001",
			4262 => "0010000111000100001000",
			4263 => "0011001001110100000100",
			4264 => "0000000100001011000001",
			4265 => "0000000100001011000001",
			4266 => "0000000100001011000001",
			4267 => "0001101000010000000100",
			4268 => "0000000100001011000001",
			4269 => "0010111101000100000100",
			4270 => "0000000100001011000001",
			4271 => "0000000100001011000001",
			4272 => "0001000100001100010100",
			4273 => "0000011101011000010000",
			4274 => "0010000101000100000100",
			4275 => "0000000100001100000101",
			4276 => "0001011110110100001000",
			4277 => "0001100100111100000100",
			4278 => "0000000100001100000101",
			4279 => "0000000100001100000101",
			4280 => "0000000100001100000101",
			4281 => "0000000100001100000101",
			4282 => "0010000111000100001100",
			4283 => "0000011011111100000100",
			4284 => "0000000100001100000101",
			4285 => "0010100001010000000100",
			4286 => "0000000100001100000101",
			4287 => "0000000100001100000101",
			4288 => "0000000100001100000101",
			4289 => "0001000000010100010100",
			4290 => "0010110000110100010000",
			4291 => "0001111011011100001100",
			4292 => "0000011011001100001000",
			4293 => "0010000101000100000100",
			4294 => "0000000100001101001001",
			4295 => "0000000100001101001001",
			4296 => "0000000100001101001001",
			4297 => "0000000100001101001001",
			4298 => "0000000100001101001001",
			4299 => "0010001111001000001100",
			4300 => "0000011011111100000100",
			4301 => "0000000100001101001001",
			4302 => "0010001001101000000100",
			4303 => "0000000100001101001001",
			4304 => "0000000100001101001001",
			4305 => "0000000100001101001001",
			4306 => "0011001011011100011100",
			4307 => "0010010010101100001100",
			4308 => "0011111111101000000100",
			4309 => "0000000100001110001101",
			4310 => "0001100100111100000100",
			4311 => "0000000100001110001101",
			4312 => "0000000100001110001101",
			4313 => "0001101000010000000100",
			4314 => "0000000100001110001101",
			4315 => "0010011001000100001000",
			4316 => "0011001001110100000100",
			4317 => "0000000100001110001101",
			4318 => "0000000100001110001101",
			4319 => "0000000100001110001101",
			4320 => "0010111111010000000100",
			4321 => "0000000100001110001101",
			4322 => "1111111100001110001101",
			4323 => "0001111000011000010100",
			4324 => "0011000100011000000100",
			4325 => "0000000100001111100001",
			4326 => "0001001000001000000100",
			4327 => "0000000100001111100001",
			4328 => "0010000111000000001000",
			4329 => "0011111000011100000100",
			4330 => "0000001100001111100001",
			4331 => "0000000100001111100001",
			4332 => "0000000100001111100001",
			4333 => "0010000110001000001100",
			4334 => "0011001001110100000100",
			4335 => "0000000100001111100001",
			4336 => "0011000100000100000100",
			4337 => "0000000100001111100001",
			4338 => "0000000100001111100001",
			4339 => "0001101000010000000100",
			4340 => "0000000100001111100001",
			4341 => "0000011001100100000100",
			4342 => "0000000100001111100001",
			4343 => "0000000100001111100001",
			4344 => "0001101000010000011000",
			4345 => "0000101101101100000100",
			4346 => "0000000100010000011101",
			4347 => "0010101000010100000100",
			4348 => "0000000100010000011101",
			4349 => "0010011011001100000100",
			4350 => "0000000100010000011101",
			4351 => "0011000001011000001000",
			4352 => "0011001010111000000100",
			4353 => "0000000100010000011101",
			4354 => "0000001100010000011101",
			4355 => "0000000100010000011101",
			4356 => "0010001111001000000100",
			4357 => "0000000100010000011101",
			4358 => "0000000100010000011101",
			4359 => "0011001011011100011000",
			4360 => "0001001100001100000100",
			4361 => "0000000100010001011001",
			4362 => "0010011011001100000100",
			4363 => "0000000100010001011001",
			4364 => "0000100011110000001100",
			4365 => "0001000011110000000100",
			4366 => "0000000100010001011001",
			4367 => "0011001010111000000100",
			4368 => "0000000100010001011001",
			4369 => "0000000100010001011001",
			4370 => "0000000100010001011001",
			4371 => "0010000110001000000100",
			4372 => "0000000100010001011001",
			4373 => "1111111100010001011001",
			4374 => "0000101000000100010100",
			4375 => "0000101101101100000100",
			4376 => "0000000100010010100101",
			4377 => "0001100101010000001100",
			4378 => "0000011001011000000100",
			4379 => "0000000100010010100101",
			4380 => "0001101111000000000100",
			4381 => "0000000100010010100101",
			4382 => "0000000100010010100101",
			4383 => "0000000100010010100101",
			4384 => "0000011101011000010000",
			4385 => "0000001010101100000100",
			4386 => "0000000100010010100101",
			4387 => "0001100100111100000100",
			4388 => "0000000100010010100101",
			4389 => "0010101000010100000100",
			4390 => "0000000100010010100101",
			4391 => "0000000100010010100101",
			4392 => "0000000100010010100101",
			4393 => "0011011100111000011000",
			4394 => "0011000100011000000100",
			4395 => "0000000100010011011001",
			4396 => "0001100100101100010000",
			4397 => "0000101101101100000100",
			4398 => "0000000100010011011001",
			4399 => "0001101111000000000100",
			4400 => "0000000100010011011001",
			4401 => "0010110110100000000100",
			4402 => "0000000100010011011001",
			4403 => "0000000100010011011001",
			4404 => "0000000100010011011001",
			4405 => "0000000100010011011001",
			4406 => "0000101000000100011000",
			4407 => "0001101001100100000100",
			4408 => "0000000100010100100101",
			4409 => "0011111000110100010000",
			4410 => "0001100101010000001100",
			4411 => "0011011110101100000100",
			4412 => "0000000100010100100101",
			4413 => "0000101100111000000100",
			4414 => "0000000100010100100101",
			4415 => "0000000100010100100101",
			4416 => "0000000100010100100101",
			4417 => "0000000100010100100101",
			4418 => "0011000111010000000100",
			4419 => "0000000100010100100101",
			4420 => "0001000110001100000100",
			4421 => "0000000100010100100101",
			4422 => "0001101000010000000100",
			4423 => "0000000100010100100101",
			4424 => "0000000100010100100101",
			4425 => "0001000100001100011100",
			4426 => "0010110000110100010100",
			4427 => "0010000101000100000100",
			4428 => "0000000100010101111001",
			4429 => "0010010011101000001100",
			4430 => "0011001111011100001000",
			4431 => "0001110110110100000100",
			4432 => "0000000100010101111001",
			4433 => "0000000100010101111001",
			4434 => "0000000100010101111001",
			4435 => "0000000100010101111001",
			4436 => "0011011010000100000100",
			4437 => "0000000100010101111001",
			4438 => "0000000100010101111001",
			4439 => "0010001111001000001100",
			4440 => "0010010101010000000100",
			4441 => "0000000100010101111001",
			4442 => "0011000101100100000100",
			4443 => "0000000100010101111001",
			4444 => "0000000100010101111001",
			4445 => "0000000100010101111001",
			4446 => "0000001011000100100100",
			4447 => "0001100101010000011000",
			4448 => "0010110110100000001100",
			4449 => "0010110000110100000100",
			4450 => "0000000100010111010101",
			4451 => "0001100101010000000100",
			4452 => "0000000100010111010101",
			4453 => "0000000100010111010101",
			4454 => "0001101000010000000100",
			4455 => "0000000100010111010101",
			4456 => "0001101000010000000100",
			4457 => "0000000100010111010101",
			4458 => "0000000100010111010101",
			4459 => "0010111111010000001000",
			4460 => "0010110010001000000100",
			4461 => "0000000100010111010101",
			4462 => "0000000100010111010101",
			4463 => "0000000100010111010101",
			4464 => "0000000000101000001000",
			4465 => "0000100110111100000100",
			4466 => "0000000100010111010101",
			4467 => "0000001100010111010101",
			4468 => "0000000100010111010101",
			4469 => "0001000000010100100000",
			4470 => "0010110000110100010100",
			4471 => "0010000101000100000100",
			4472 => "0000000100011000110001",
			4473 => "0000011010011000001100",
			4474 => "0001110110110100001000",
			4475 => "0010101000100100000100",
			4476 => "0000000100011000110001",
			4477 => "0000000100011000110001",
			4478 => "0000000100011000110001",
			4479 => "0000000100011000110001",
			4480 => "0010100001010000001000",
			4481 => "0010101000100100000100",
			4482 => "0000000100011000110001",
			4483 => "0000000100011000110001",
			4484 => "0000000100011000110001",
			4485 => "0010001111001000001100",
			4486 => "0000011011111100000100",
			4487 => "0000000100011000110001",
			4488 => "0010001001101000000100",
			4489 => "0000000100011000110001",
			4490 => "0000000100011000110001",
			4491 => "0000000100011000110001",
			4492 => "0001000000010100010100",
			4493 => "0000001010101100000100",
			4494 => "0000000100011010000101",
			4495 => "0010011000100100001100",
			4496 => "0001110111110000001000",
			4497 => "0010101000010100000100",
			4498 => "0000000100011010000101",
			4499 => "0000000100011010000101",
			4500 => "0000000100011010000101",
			4501 => "0000000100011010000101",
			4502 => "0010100101000100010100",
			4503 => "0010011011001100000100",
			4504 => "0000000100011010000101",
			4505 => "0000000010011000000100",
			4506 => "0000000100011010000101",
			4507 => "0001100100101100001000",
			4508 => "0001111011000000000100",
			4509 => "0000000100011010000101",
			4510 => "0000000100011010000101",
			4511 => "0000000100011010000101",
			4512 => "0000000100011010000101",
			4513 => "0011011010000100100000",
			4514 => "0011001001110100001000",
			4515 => "0001000000101100000100",
			4516 => "0000000100011011010001",
			4517 => "0000000100011011010001",
			4518 => "0001001110100100000100",
			4519 => "0000000100011011010001",
			4520 => "0010000111000100010000",
			4521 => "0011101000011100001100",
			4522 => "0011000001011000001000",
			4523 => "0000011110010100000100",
			4524 => "0000000100011011010001",
			4525 => "0000000100011011010001",
			4526 => "0000000100011011010001",
			4527 => "0000000100011011010001",
			4528 => "0000000100011011010001",
			4529 => "0000011101011000000100",
			4530 => "0000000100011011010001",
			4531 => "0000000100011011010001",
			4532 => "0011011010000100011100",
			4533 => "0010011001111100000100",
			4534 => "0000000100011100011101",
			4535 => "0001101001111100010100",
			4536 => "0000100110111000000100",
			4537 => "0000000100011100011101",
			4538 => "0011000100000100001100",
			4539 => "0000101010110100001000",
			4540 => "0011001001110100000100",
			4541 => "0000000100011100011101",
			4542 => "0000000100011100011101",
			4543 => "0000000100011100011101",
			4544 => "0000000100011100011101",
			4545 => "0000000100011100011101",
			4546 => "0011100011010100001000",
			4547 => "0001101000010000000100",
			4548 => "0000000100011100011101",
			4549 => "0000000100011100011101",
			4550 => "0000000100011100011101",
			4551 => "0001000011011000100100",
			4552 => "0010000110001000011000",
			4553 => "0010010111101100000100",
			4554 => "0000000100011101111001",
			4555 => "0010110110100000010000",
			4556 => "0011101000011100001100",
			4557 => "0000110001011100000100",
			4558 => "0000000100011101111001",
			4559 => "0010110100010000000100",
			4560 => "0000000100011101111001",
			4561 => "0000000100011101111001",
			4562 => "0000000100011101111001",
			4563 => "0000000100011101111001",
			4564 => "0001001001000000001000",
			4565 => "0000111110111000000100",
			4566 => "0000000100011101111001",
			4567 => "0000000100011101111001",
			4568 => "0000000100011101111001",
			4569 => "0010100101000100001000",
			4570 => "0001101000010000000100",
			4571 => "0000000100011101111001",
			4572 => "0000001100011101111001",
			4573 => "0000000100011101111001",
			4574 => "0001000100001100011100",
			4575 => "0010000101000100000100",
			4576 => "0000000100011111001101",
			4577 => "0001011110110100010100",
			4578 => "0010010111110100010000",
			4579 => "0001100100111100000100",
			4580 => "0000000100011111001101",
			4581 => "0010111101000100001000",
			4582 => "0000000001110100000100",
			4583 => "0000000100011111001101",
			4584 => "0000000100011111001101",
			4585 => "0000000100011111001101",
			4586 => "0000000100011111001101",
			4587 => "0000000100011111001101",
			4588 => "0010000111000100001100",
			4589 => "0010010101010000000100",
			4590 => "0000000100011111001101",
			4591 => "0010100001010000000100",
			4592 => "0000000100011111001101",
			4593 => "0000000100011111001101",
			4594 => "0000000100011111001101",
			4595 => "0011001011011100100100",
			4596 => "0001000100001100001100",
			4597 => "0001111011011100001000",
			4598 => "0010111110101100000100",
			4599 => "0000000100100000100001",
			4600 => "0000000100100000100001",
			4601 => "0000000100100000100001",
			4602 => "0010100101000100010100",
			4603 => "0010011011001100000100",
			4604 => "0000000100100000100001",
			4605 => "0000101010110100001100",
			4606 => "0011011100000000001000",
			4607 => "0001111011000000000100",
			4608 => "0000000100100000100001",
			4609 => "0000000100100000100001",
			4610 => "0000000100100000100001",
			4611 => "0000000100100000100001",
			4612 => "0000000100100000100001",
			4613 => "0010000110001000000100",
			4614 => "0000000100100000100001",
			4615 => "1111111100100000100001",
			4616 => "0011111111101000011000",
			4617 => "0000011001011000000100",
			4618 => "0000000100100001111101",
			4619 => "0000101101101100000100",
			4620 => "0000000100100001111101",
			4621 => "0001100101010000001100",
			4622 => "0011001010111000000100",
			4623 => "0000000100100001111101",
			4624 => "0000011010011000000100",
			4625 => "0000000100100001111101",
			4626 => "0000000100100001111101",
			4627 => "0000000100100001111101",
			4628 => "0010000001010100000100",
			4629 => "0000000100100001111101",
			4630 => "0011100011010100010000",
			4631 => "0010101000010100000100",
			4632 => "0000000100100001111101",
			4633 => "0000001010101100000100",
			4634 => "0000000100100001111101",
			4635 => "0000110011101100000100",
			4636 => "0000000100100001111101",
			4637 => "0000000100100001111101",
			4638 => "0000000100100001111101",
			4639 => "0000101011110000011000",
			4640 => "0000101101101100000100",
			4641 => "0000000100100011110001",
			4642 => "0001101000010000010000",
			4643 => "0001101111000000000100",
			4644 => "0000000100100011110001",
			4645 => "0011001010111000000100",
			4646 => "0000000100100011110001",
			4647 => "0000000001110100000100",
			4648 => "0000000100100011110001",
			4649 => "0000001100100011110001",
			4650 => "0000000100100011110001",
			4651 => "0010001111001000011000",
			4652 => "0000000111000000001100",
			4653 => "0000001010101100000100",
			4654 => "0000000100100011110001",
			4655 => "0000000111000000000100",
			4656 => "0000000100100011110001",
			4657 => "0000000100100011110001",
			4658 => "0010110100010000000100",
			4659 => "0000000100100011110001",
			4660 => "0010110111100000000100",
			4661 => "0000000100100011110001",
			4662 => "0000000100100011110001",
			4663 => "0011100011010100001000",
			4664 => "0000110011101100000100",
			4665 => "0000000100100011110001",
			4666 => "0000000100100011110001",
			4667 => "0000000100100011110001",
			4668 => "0001000011011000101000",
			4669 => "0000011010011000011000",
			4670 => "0010000101000100000100",
			4671 => "0000000100100101010101",
			4672 => "0001000111011100010000",
			4673 => "0010110110100000001100",
			4674 => "0001010110010000001000",
			4675 => "0010010011101000000100",
			4676 => "0000000100100101010101",
			4677 => "0000000100100101010101",
			4678 => "0000000100100101010101",
			4679 => "0000000100100101010101",
			4680 => "0000000100100101010101",
			4681 => "0010111110101000001100",
			4682 => "0010000110001000001000",
			4683 => "0010111010010100000100",
			4684 => "0000000100100101010101",
			4685 => "0000000100100101010101",
			4686 => "0000000100100101010101",
			4687 => "0000000100100101010101",
			4688 => "0010100101000100001000",
			4689 => "0000011001011000000100",
			4690 => "0000000100100101010101",
			4691 => "0000001100100101010101",
			4692 => "0000000100100101010101",
			4693 => "0010011010100000001000",
			4694 => "0011111110100100000100",
			4695 => "0000000100100110110001",
			4696 => "0000000100100110110001",
			4697 => "0011101000011100011000",
			4698 => "0001101001111100010100",
			4699 => "0010110100010000000100",
			4700 => "0000000100100110110001",
			4701 => "0000111100001100001100",
			4702 => "0010110110100000001000",
			4703 => "0001011001010000000100",
			4704 => "0000000100100110110001",
			4705 => "0000000100100110110001",
			4706 => "0000000100100110110001",
			4707 => "0000000100100110110001",
			4708 => "0000000100100110110001",
			4709 => "0010011000100100001100",
			4710 => "0001110111110000001000",
			4711 => "0001000100001100000100",
			4712 => "0000000100100110110001",
			4713 => "0000000100100110110001",
			4714 => "0000000100100110110001",
			4715 => "0000000100100110110001",
			4716 => "0001011110000100010000",
			4717 => "0011001010111000000100",
			4718 => "0000000100101000011101",
			4719 => "0001001111100000000100",
			4720 => "0000000100101000011101",
			4721 => "0010001101010000000100",
			4722 => "0000001100101000011101",
			4723 => "0000000100101000011101",
			4724 => "0000011010011000011000",
			4725 => "0001100100111100000100",
			4726 => "0000000100101000011101",
			4727 => "0001111111011100000100",
			4728 => "0000000100101000011101",
			4729 => "0010010011101000001100",
			4730 => "0001011110110100001000",
			4731 => "0010000101000100000100",
			4732 => "0000000100101000011101",
			4733 => "0000000100101000011101",
			4734 => "0000000100101000011101",
			4735 => "0000000100101000011101",
			4736 => "0001100100101100001100",
			4737 => "0001110111010000000100",
			4738 => "0000000100101000011101",
			4739 => "0000001010101100000100",
			4740 => "0000000100101000011101",
			4741 => "0000000100101000011101",
			4742 => "0000000100101000011101",
			4743 => "0000001011000100110000",
			4744 => "0011000111010000100000",
			4745 => "0001010111111100001100",
			4746 => "0000100110111000001000",
			4747 => "0000000001110100000100",
			4748 => "0000000100101010001001",
			4749 => "0000000100101010001001",
			4750 => "0000000100101010001001",
			4751 => "0001100100101100010000",
			4752 => "0011011111010100001100",
			4753 => "0000011101111100000100",
			4754 => "0000000100101010001001",
			4755 => "0000110010111000000100",
			4756 => "0000000100101010001001",
			4757 => "0000000100101010001001",
			4758 => "0000000100101010001001",
			4759 => "0000000100101010001001",
			4760 => "0000101000000100000100",
			4761 => "0000000100101010001001",
			4762 => "0010011000100100001000",
			4763 => "0001101000010000000100",
			4764 => "0000000100101010001001",
			4765 => "0000000100101010001001",
			4766 => "0000000100101010001001",
			4767 => "0000000000101000000100",
			4768 => "0000001100101010001001",
			4769 => "0000000100101010001001",
			4770 => "0000101011110000011100",
			4771 => "0000101101101100000100",
			4772 => "0000000100101011111101",
			4773 => "0001101000010000010100",
			4774 => "0001101111000000000100",
			4775 => "0000000100101011111101",
			4776 => "0011001010111000000100",
			4777 => "0000000100101011111101",
			4778 => "0001000110111000000100",
			4779 => "0000000100101011111101",
			4780 => "0010101000100100000100",
			4781 => "0000000100101011111101",
			4782 => "0000001100101011111101",
			4783 => "0000000100101011111101",
			4784 => "0011011100000000001100",
			4785 => "0010010100101100000100",
			4786 => "0000000100101011111101",
			4787 => "0000010111101000000100",
			4788 => "0000000100101011111101",
			4789 => "0000000100101011111101",
			4790 => "0010011000100100010000",
			4791 => "0001101000010000000100",
			4792 => "0000000100101011111101",
			4793 => "0010000001010100000100",
			4794 => "0000000100101011111101",
			4795 => "0001001110100100000100",
			4796 => "0000000100101011111101",
			4797 => "0000000100101011111101",
			4798 => "0000000100101011111101",
			4799 => "0000011100011000100100",
			4800 => "0010011010100000010000",
			4801 => "0000011011111100000100",
			4802 => "1111111100101110010001",
			4803 => "0000101110000000000100",
			4804 => "1111111100101110010001",
			4805 => "0011101011101100000100",
			4806 => "0000001100101110010001",
			4807 => "1111111100101110010001",
			4808 => "0001111111011100000100",
			4809 => "1111111100101110010001",
			4810 => "0011100010010100001000",
			4811 => "0000010100110100000100",
			4812 => "0000010100101110010001",
			4813 => "0000001100101110010001",
			4814 => "0011001000011000000100",
			4815 => "1111111100101110010001",
			4816 => "0000000100101110010001",
			4817 => "0011011100010100001100",
			4818 => "0011101101101100001000",
			4819 => "0001111000011000000100",
			4820 => "0000000100101110010001",
			4821 => "0000000100101110010001",
			4822 => "1111111100101110010001",
			4823 => "0010101100011100010100",
			4824 => "0001110111010000000100",
			4825 => "0000000100101110010001",
			4826 => "0011000101100100001100",
			4827 => "0010111110101000001000",
			4828 => "0010011010100100000100",
			4829 => "0000001100101110010001",
			4830 => "0000001100101110010001",
			4831 => "0000000100101110010001",
			4832 => "0000000100101110010001",
			4833 => "0001011100010000000100",
			4834 => "1111111100101110010001",
			4835 => "0000000100101110010001",
			4836 => "0010011010100100100000",
			4837 => "0010011010100100010100",
			4838 => "0010011001111100000100",
			4839 => "1111111100110000010101",
			4840 => "0001110001101000000100",
			4841 => "1111111100110000010101",
			4842 => "0011101111101000001000",
			4843 => "0000101110000000000100",
			4844 => "1111111100110000010101",
			4845 => "0000001100110000010101",
			4846 => "1111111100110000010101",
			4847 => "0001010101110000000100",
			4848 => "1111111100110000010101",
			4849 => "0000111011110000000100",
			4850 => "0000001100110000010101",
			4851 => "0000000100110000010101",
			4852 => "0010110101110100000100",
			4853 => "1111111100110000010101",
			4854 => "0010000110001000011000",
			4855 => "0001110111010000001000",
			4856 => "0001010101110000000100",
			4857 => "1111111100110000010101",
			4858 => "0000000100110000010101",
			4859 => "0011000101100100001100",
			4860 => "0010111110101000001000",
			4861 => "0010011010100100000100",
			4862 => "0000001100110000010101",
			4863 => "0000001100110000010101",
			4864 => "0000001100110000010101",
			4865 => "0000000100110000010101",
			4866 => "0001000111011100000100",
			4867 => "1111111100110000010101",
			4868 => "0000000100110000010101",
			4869 => "0000010100110100101100",
			4870 => "0010011010100100011100",
			4871 => "0000010101011100000100",
			4872 => "1111111100110010100001",
			4873 => "0001000011110100010000",
			4874 => "0001001110111000000100",
			4875 => "1111111100110010100001",
			4876 => "0001001110111000000100",
			4877 => "0000001100110010100001",
			4878 => "0010111011110100000100",
			4879 => "0000000100110010100001",
			4880 => "1111111100110010100001",
			4881 => "0011001000011000000100",
			4882 => "0000010100110010100001",
			4883 => "1111111100110010100001",
			4884 => "0001110111010000001000",
			4885 => "0011001001110100000100",
			4886 => "1111111100110010100001",
			4887 => "0000000100110010100001",
			4888 => "0011101011110000000100",
			4889 => "0000001100110010100001",
			4890 => "0000000100110010100001",
			4891 => "0011011100010100000100",
			4892 => "1111111100110010100001",
			4893 => "0001100100101100010100",
			4894 => "0011001001110100000100",
			4895 => "0000000100110010100001",
			4896 => "0001100100101100001100",
			4897 => "0001001111100000001000",
			4898 => "0001100101010000000100",
			4899 => "0000001100110010100001",
			4900 => "0000001100110010100001",
			4901 => "0000010100110010100001",
			4902 => "0000000100110010100001",
			4903 => "1111111100110010100001",
			4904 => "0000011100011000110000",
			4905 => "0010011010100100101000",
			4906 => "0010011010100100011100",
			4907 => "0001100100111100000100",
			4908 => "1101110100110100111101",
			4909 => "0011111110000000010000",
			4910 => "0000101110000000001000",
			4911 => "0001111000011000000100",
			4912 => "1101110100110100111101",
			4913 => "1101110100110100111101",
			4914 => "0000011011111100000100",
			4915 => "1101110100110100111101",
			4916 => "1110011100110100111101",
			4917 => "0001101000010000000100",
			4918 => "1101110100110100111101",
			4919 => "1101110100110100111101",
			4920 => "0011000001101000001000",
			4921 => "0001011001010000000100",
			4922 => "1101110100110100111101",
			4923 => "1101111100110100111101",
			4924 => "1110010100110100111101",
			4925 => "0001101000010000000100",
			4926 => "1110101100110100111101",
			4927 => "1101110100110100111101",
			4928 => "0001010111111100001000",
			4929 => "0001110111010000000100",
			4930 => "1101110100110100111101",
			4931 => "1110010100110100111101",
			4932 => "0010001111001000010000",
			4933 => "0001110000011100001000",
			4934 => "0010101001000100000100",
			4935 => "1110101100110100111101",
			4936 => "1110010100110100111101",
			4937 => "0011001011011100000100",
			4938 => "1110110100110100111101",
			4939 => "1110100100110100111101",
			4940 => "0001100100101100000100",
			4941 => "1110000100110100111101",
			4942 => "1101110100110100111101",
			4943 => "0011001001110100001000",
			4944 => "0010100110011100000100",
			4945 => "0000000100110111000001",
			4946 => "0000000100110111000001",
			4947 => "0011010110111100100000",
			4948 => "0000011100011000011000",
			4949 => "0011011110110100010000",
			4950 => "0011011010001000000100",
			4951 => "0000000100110111000001",
			4952 => "0000001110111100001000",
			4953 => "0000001111001000000100",
			4954 => "0000000100110111000001",
			4955 => "0000000100110111000001",
			4956 => "0000000100110111000001",
			4957 => "0000001010101100000100",
			4958 => "0000000100110111000001",
			4959 => "0000000100110111000001",
			4960 => "0010110001001000000100",
			4961 => "0000000100110111000001",
			4962 => "0000000100110111000001",
			4963 => "0010010011101000001000",
			4964 => "0011000100000100000100",
			4965 => "0000000100110111000001",
			4966 => "0000000100110111000001",
			4967 => "0011000111010000010000",
			4968 => "0001011110110100001100",
			4969 => "0000110101000000000100",
			4970 => "0000000100110111000001",
			4971 => "0000011111000000000100",
			4972 => "0000000100110111000001",
			4973 => "0000000100110111000001",
			4974 => "0000000100110111000001",
			4975 => "0000000100110111000001",
			4976 => "0011001011000000000100",
			4977 => "1111111100111000110101",
			4978 => "0001101000010000001100",
			4979 => "0011110010010100000100",
			4980 => "0000000100111000110101",
			4981 => "0000010100110100000100",
			4982 => "0000000100111000110101",
			4983 => "0000000100111000110101",
			4984 => "0000001010101100010000",
			4985 => "0011111000110100000100",
			4986 => "0000000100111000110101",
			4987 => "0011000111010000001000",
			4988 => "0000001010101100000100",
			4989 => "0000000100111000110101",
			4990 => "0000000100111000110101",
			4991 => "0000000100111000110101",
			4992 => "0001100101010000010000",
			4993 => "0001001100001100000100",
			4994 => "0000000100111000110101",
			4995 => "0000011011111100000100",
			4996 => "0000000100111000110101",
			4997 => "0011100110001100000100",
			4998 => "0000000100111000110101",
			4999 => "0000000100111000110101",
			5000 => "0000011010011000000100",
			5001 => "0000000100111000110101",
			5002 => "0001100100101100000100",
			5003 => "0000000100111000110101",
			5004 => "0000000100111000110101",
			5005 => "0000010100110100110100",
			5006 => "0010011010100100100100",
			5007 => "0000010101011100000100",
			5008 => "1111111100111011001001",
			5009 => "0001000011110100010000",
			5010 => "0001001110111000000100",
			5011 => "1111111100111011001001",
			5012 => "0001001110111000000100",
			5013 => "0000001100111011001001",
			5014 => "0010111011110100000100",
			5015 => "0000000100111011001001",
			5016 => "1111111100111011001001",
			5017 => "0000100110001100000100",
			5018 => "0000010100111011001001",
			5019 => "0001001011100000001000",
			5020 => "0001010010000100000100",
			5021 => "0000001100111011001001",
			5022 => "0000000100111011001001",
			5023 => "1111111100111011001001",
			5024 => "0001110111010000001000",
			5025 => "0011001001110100000100",
			5026 => "1111111100111011001001",
			5027 => "0000000100111011001001",
			5028 => "0011101011110000000100",
			5029 => "0000010100111011001001",
			5030 => "0000000100111011001001",
			5031 => "0011011100010100000100",
			5032 => "1111111100111011001001",
			5033 => "0010000001110100010000",
			5034 => "0011001001110100000100",
			5035 => "0000000100111011001001",
			5036 => "0010001111001000001000",
			5037 => "0011001011011100000100",
			5038 => "0000001100111011001001",
			5039 => "0000001100111011001001",
			5040 => "0000001100111011001001",
			5041 => "1111111100111011001001",
			5042 => "0000011100011000100100",
			5043 => "0000010101011100000100",
			5044 => "1111111100111101110101",
			5045 => "0001000100001100010100",
			5046 => "0001110000011100001000",
			5047 => "0001011110010000000100",
			5048 => "1111111100111101110101",
			5049 => "0000000100111101110101",
			5050 => "0001101000010000001000",
			5051 => "0000011101111100000100",
			5052 => "1111111100111101110101",
			5053 => "0000001100111101110101",
			5054 => "1111111100111101110101",
			5055 => "0000100110001100000100",
			5056 => "0000010100111101110101",
			5057 => "0001100101010000000100",
			5058 => "0000001100111101110101",
			5059 => "1111111100111101110101",
			5060 => "0011001001110100001100",
			5061 => "0010101001000100001000",
			5062 => "0001001100001100000100",
			5063 => "1111111100111101110101",
			5064 => "0000001100111101110101",
			5065 => "1111111100111101110101",
			5066 => "0001100100101100100000",
			5067 => "0010110001001000001100",
			5068 => "0011100110111000000100",
			5069 => "0000001100111101110101",
			5070 => "0010010011101000000100",
			5071 => "1111111100111101110101",
			5072 => "0000001100111101110101",
			5073 => "0001101001111100001100",
			5074 => "0010110110100000000100",
			5075 => "0000001100111101110101",
			5076 => "0010111101000100000100",
			5077 => "0000001100111101110101",
			5078 => "0000001100111101110101",
			5079 => "0000011011001100000100",
			5080 => "0000000100111101110101",
			5081 => "0000001100111101110101",
			5082 => "0001000011011000000100",
			5083 => "1111111100111101110101",
			5084 => "0000000100111101110101",
			5085 => "0000010111101000000100",
			5086 => "1111111100111111110001",
			5087 => "0001000011110000100100",
			5088 => "0010110000110100010000",
			5089 => "0010000101000100000100",
			5090 => "0000000100111111110001",
			5091 => "0000011010011000001000",
			5092 => "0011001111011100000100",
			5093 => "1111111100111111110001",
			5094 => "0000000100111111110001",
			5095 => "0000000100111111110001",
			5096 => "0000111100001100001100",
			5097 => "0010111101000100001000",
			5098 => "0010101001000100000100",
			5099 => "0000000100111111110001",
			5100 => "0000000100111111110001",
			5101 => "0000000100111111110001",
			5102 => "0010101000010100000100",
			5103 => "0000000100111111110001",
			5104 => "0000000100111111110001",
			5105 => "0001100100101100010100",
			5106 => "0011001011011100010000",
			5107 => "0011001001110100000100",
			5108 => "0000000100111111110001",
			5109 => "0011100110001100001000",
			5110 => "0000010100110100000100",
			5111 => "0000000100111111110001",
			5112 => "0000000100111111110001",
			5113 => "0000000100111111110001",
			5114 => "0000000100111111110001",
			5115 => "0000000100111111110001",
			5116 => "0000100011000000001000",
			5117 => "0010110001001000000100",
			5118 => "1111111101000010001101",
			5119 => "0000000101000010001101",
			5120 => "0001100101010000101100",
			5121 => "0011011111010100011100",
			5122 => "0000011010011000011000",
			5123 => "0011100110111000001100",
			5124 => "0010010100111100000100",
			5125 => "0000000101000010001101",
			5126 => "0001001000001000000100",
			5127 => "0000000101000010001101",
			5128 => "0000000101000010001101",
			5129 => "0001111011011100001000",
			5130 => "0000000010011000000100",
			5131 => "0000000101000010001101",
			5132 => "0000000101000010001101",
			5133 => "0000000101000010001101",
			5134 => "0000001101000010001101",
			5135 => "0010010011101000001000",
			5136 => "0000011100011000000100",
			5137 => "0000000101000010001101",
			5138 => "0000000101000010001101",
			5139 => "0000000111000000000100",
			5140 => "1111111101000010001101",
			5141 => "0000000101000010001101",
			5142 => "0010011000100100001100",
			5143 => "0001000011101100001000",
			5144 => "0010100110011000000100",
			5145 => "0000000101000010001101",
			5146 => "1111111101000010001101",
			5147 => "0000000101000010001101",
			5148 => "0010011000010100001000",
			5149 => "0000011001100100000100",
			5150 => "0000000101000010001101",
			5151 => "0000000101000010001101",
			5152 => "0010100110011100000100",
			5153 => "0000000101000010001101",
			5154 => "0000000101000010001101",
			5155 => "0000010101011100000100",
			5156 => "1111111101000100001001",
			5157 => "0001100101010000101100",
			5158 => "0010010011101000011000",
			5159 => "0010011010100100010000",
			5160 => "0000000010011000001100",
			5161 => "0001100100111100000100",
			5162 => "0000000101000100001001",
			5163 => "0000011100011000000100",
			5164 => "0000000101000100001001",
			5165 => "0000000101000100001001",
			5166 => "0000000101000100001001",
			5167 => "0011011100010100000100",
			5168 => "0000000101000100001001",
			5169 => "0000001101000100001001",
			5170 => "0010101000010100010000",
			5171 => "0011101110000000000100",
			5172 => "0000000101000100001001",
			5173 => "0011001010001100001000",
			5174 => "0011010111011000000100",
			5175 => "0000000101000100001001",
			5176 => "1111111101000100001001",
			5177 => "0000000101000100001001",
			5178 => "0000000101000100001001",
			5179 => "0001111111011100000100",
			5180 => "0000000101000100001001",
			5181 => "0000011101011000000100",
			5182 => "0000000101000100001001",
			5183 => "0010000111000100000100",
			5184 => "0000000101000100001001",
			5185 => "0000000101000100001001",
			5186 => "0000100011000000001100",
			5187 => "0010000101000100000100",
			5188 => "0000000101000110011101",
			5189 => "0011111111101000000100",
			5190 => "0000000101000110011101",
			5191 => "0000000101000110011101",
			5192 => "0001010110010000011000",
			5193 => "0001101001111100010100",
			5194 => "0010010100111100000100",
			5195 => "0000000101000110011101",
			5196 => "0011110010111000001100",
			5197 => "0001001110100100000100",
			5198 => "0000000101000110011101",
			5199 => "0001100100111100000100",
			5200 => "0000000101000110011101",
			5201 => "0000000101000110011101",
			5202 => "0000000101000110011101",
			5203 => "0000000101000110011101",
			5204 => "0001110100010000010100",
			5205 => "0010010011101000000100",
			5206 => "0000000101000110011101",
			5207 => "0000110101000000000100",
			5208 => "0000000101000110011101",
			5209 => "0010111101000100001000",
			5210 => "0011010110111100000100",
			5211 => "0000000101000110011101",
			5212 => "0000000101000110011101",
			5213 => "0000000101000110011101",
			5214 => "0001100100101100010000",
			5215 => "0011111000011100000100",
			5216 => "0000000101000110011101",
			5217 => "0011101011110000000100",
			5218 => "0000000101000110011101",
			5219 => "0010011010100100000100",
			5220 => "0000000101000110011101",
			5221 => "0000000101000110011101",
			5222 => "0000000101000110011101",
			5223 => "0010010100101100001000",
			5224 => "0001001100111100000100",
			5225 => "1111111101001000100001",
			5226 => "0000000101001000100001",
			5227 => "0001110111010000001000",
			5228 => "0000000010111100000100",
			5229 => "0000000101001000100001",
			5230 => "0000000101001000100001",
			5231 => "0010110110100000011000",
			5232 => "0011000100000100010000",
			5233 => "0011101000001000001100",
			5234 => "0000000001110100000100",
			5235 => "0000000101001000100001",
			5236 => "0010010111101100000100",
			5237 => "0000000101001000100001",
			5238 => "0000001101001000100001",
			5239 => "0000000101001000100001",
			5240 => "0010010010101100000100",
			5241 => "0000000101001000100001",
			5242 => "0000000101001000100001",
			5243 => "0011101110000000001000",
			5244 => "0001001100001100000100",
			5245 => "0000000101001000100001",
			5246 => "0000000101001000100001",
			5247 => "0001100100101100010000",
			5248 => "0001110100010000001000",
			5249 => "0001110010001000000100",
			5250 => "0000000101001000100001",
			5251 => "0000000101001000100001",
			5252 => "0000011100011000000100",
			5253 => "0000000101001000100001",
			5254 => "0000001101001000100001",
			5255 => "0000000101001000100001",
			5256 => "0011001011000000000100",
			5257 => "0000000101001010011101",
			5258 => "0001101001111100110000",
			5259 => "0001000011110000011100",
			5260 => "0010110000110100010000",
			5261 => "0001100100111100000100",
			5262 => "0000000101001010011101",
			5263 => "0000011010011000001000",
			5264 => "0011001111011100000100",
			5265 => "0000000101001010011101",
			5266 => "0000000101001010011101",
			5267 => "0000000101001010011101",
			5268 => "0010110110100000001000",
			5269 => "0000010100110100000100",
			5270 => "0000000101001010011101",
			5271 => "0000000101001010011101",
			5272 => "0000000101001010011101",
			5273 => "0011101000001000010000",
			5274 => "0010010101010000000100",
			5275 => "0000000101001010011101",
			5276 => "0001110001101000000100",
			5277 => "0000000101001010011101",
			5278 => "0000011011111100000100",
			5279 => "0000000101001010011101",
			5280 => "0000000101001010011101",
			5281 => "0000000101001010011101",
			5282 => "0000011001100100000100",
			5283 => "0000000101001010011101",
			5284 => "0010000111000100000100",
			5285 => "0000000101001010011101",
			5286 => "0000000101001010011101",
			5287 => "0011001011000000000100",
			5288 => "1111111101001100100001",
			5289 => "0001101000010000010000",
			5290 => "0000110001011100000100",
			5291 => "0000000101001100100001",
			5292 => "0000010100110100000100",
			5293 => "0000000101001100100001",
			5294 => "0011110010010100000100",
			5295 => "0000000101001100100001",
			5296 => "0000000101001100100001",
			5297 => "0000001010101100010000",
			5298 => "0011111000110100000100",
			5299 => "0000000101001100100001",
			5300 => "0011000111010000001000",
			5301 => "0010000001010100000100",
			5302 => "0000000101001100100001",
			5303 => "0000000101001100100001",
			5304 => "0000000101001100100001",
			5305 => "0001100101010000010000",
			5306 => "0010101000010100000100",
			5307 => "0000000101001100100001",
			5308 => "0000011011111100000100",
			5309 => "0000000101001100100001",
			5310 => "0011110011001100000100",
			5311 => "0000000101001100100001",
			5312 => "0000000101001100100001",
			5313 => "0000011010011000000100",
			5314 => "0000000101001100100001",
			5315 => "0001100100101100001000",
			5316 => "0000000011010000000100",
			5317 => "0000000101001100100001",
			5318 => "0000000101001100100001",
			5319 => "0000000101001100100001",
			5320 => "0010010100111100000100",
			5321 => "1111111101001110110101",
			5322 => "0001100101010000110000",
			5323 => "0000000111000000100000",
			5324 => "0000111100001100011000",
			5325 => "0001110001011000001100",
			5326 => "0001001110100100001000",
			5327 => "0010110000110100000100",
			5328 => "1111111101001110110101",
			5329 => "0000000101001110110101",
			5330 => "0000000101001110110101",
			5331 => "0001110101110100001000",
			5332 => "0000010100110100000100",
			5333 => "0000000101001110110101",
			5334 => "0000001101001110110101",
			5335 => "0000000101001110110101",
			5336 => "0010010011101000000100",
			5337 => "0000000101001110110101",
			5338 => "1111111101001110110101",
			5339 => "0001000110001100000100",
			5340 => "0000000101001110110101",
			5341 => "0011111101001000001000",
			5342 => "0011111111100100000100",
			5343 => "0000000101001110110101",
			5344 => "0000001101001110110101",
			5345 => "0000000101001110110101",
			5346 => "0010011000100100001100",
			5347 => "0001000011101100001000",
			5348 => "0010001100000100000100",
			5349 => "0000000101001110110101",
			5350 => "1111111101001110110101",
			5351 => "0000000101001110110101",
			5352 => "0010000111000100001000",
			5353 => "0011001000011000000100",
			5354 => "0000000101001110110101",
			5355 => "0000000101001110110101",
			5356 => "0000000101001110110101",
			5357 => "0000010100110100101000",
			5358 => "0001100100111100000100",
			5359 => "1111111101010010010001",
			5360 => "0011110110111000010000",
			5361 => "0001000111011100001000",
			5362 => "0000111100111000000100",
			5363 => "1111111101010010010001",
			5364 => "0000000101010010010001",
			5365 => "0010011011001100000100",
			5366 => "0000000101010010010001",
			5367 => "0000001101010010010001",
			5368 => "0001101000010000001000",
			5369 => "0001101000010000000100",
			5370 => "0000000101010010010001",
			5371 => "0000000101010010010001",
			5372 => "0000111000101000001000",
			5373 => "0000110001011100000100",
			5374 => "0000000101010010010001",
			5375 => "0000000101010010010001",
			5376 => "1111111101010010010001",
			5377 => "0000011100011000100100",
			5378 => "0001100100111100010000",
			5379 => "0000110001011100000100",
			5380 => "1111111101010010010001",
			5381 => "0011110010010100001000",
			5382 => "0000101111101000000100",
			5383 => "0000001101010010010001",
			5384 => "0000000101010010010001",
			5385 => "0000001101010010010001",
			5386 => "0001001110111000010000",
			5387 => "0011101000101000001000",
			5388 => "0011011110010000000100",
			5389 => "0000000101010010010001",
			5390 => "0000000101010010010001",
			5391 => "0001001000011100000100",
			5392 => "0000000101010010010001",
			5393 => "1111111101010010010001",
			5394 => "0000000101010010010001",
			5395 => "0010000110001000011100",
			5396 => "0011011010000100010100",
			5397 => "0001010101110000000100",
			5398 => "0000000101010010010001",
			5399 => "0011000100000100001000",
			5400 => "0011101000001000000100",
			5401 => "0000001101010010010001",
			5402 => "0000000101010010010001",
			5403 => "0011010110111100000100",
			5404 => "0000001101010010010001",
			5405 => "0000000101010010010001",
			5406 => "0010000001010100000100",
			5407 => "1111111101010010010001",
			5408 => "0000001101010010010001",
			5409 => "0000100101010100000100",
			5410 => "0000000101010010010001",
			5411 => "1111111101010010010001",
			5412 => "0011001000000000001100",
			5413 => "0000100110111000000100",
			5414 => "1111111101010101001101",
			5415 => "0000100110111000000100",
			5416 => "0000000101010101001101",
			5417 => "1111111101010101001101",
			5418 => "0000011101011001000000",
			5419 => "0000111110100100100100",
			5420 => "0010011001111100001100",
			5421 => "0011001000000000001000",
			5422 => "0000010101011100000100",
			5423 => "0000000101010101001101",
			5424 => "0000000101010101001101",
			5425 => "1111111101010101001101",
			5426 => "0001100100111100001000",
			5427 => "0011111000101000000100",
			5428 => "0000000101010101001101",
			5429 => "0000001101010101001101",
			5430 => "0001001101001000001000",
			5431 => "0000011100011000000100",
			5432 => "1111111101010101001101",
			5433 => "0000000101010101001101",
			5434 => "0001101001111100000100",
			5435 => "0000001101010101001101",
			5436 => "0000000101010101001101",
			5437 => "0001110110110100010000",
			5438 => "0010010010101100001000",
			5439 => "0001100101010000000100",
			5440 => "0000000101010101001101",
			5441 => "0000000101010101001101",
			5442 => "0010010011101000000100",
			5443 => "1111111101010101001101",
			5444 => "1111110101010101001101",
			5445 => "0010100110011000000100",
			5446 => "0000001101010101001101",
			5447 => "0011011100010000000100",
			5448 => "0000000101010101001101",
			5449 => "1111111101010101001101",
			5450 => "0010101000010100001000",
			5451 => "0010010011101000000100",
			5452 => "0000001101010101001101",
			5453 => "1111111101010101001101",
			5454 => "0001100100101100001000",
			5455 => "0011011110110100000100",
			5456 => "0000000101010101001101",
			5457 => "0000001101010101001101",
			5458 => "0000000101010101001101",
			5459 => "0011001011000000000100",
			5460 => "1111111101010111110001",
			5461 => "0000110110001100110100",
			5462 => "0001001100001100011100",
			5463 => "0001101000010000001100",
			5464 => "0010011010100100000100",
			5465 => "0000000101010111110001",
			5466 => "0001110111010000000100",
			5467 => "0000000101010111110001",
			5468 => "0000000101010111110001",
			5469 => "0011001010001100001100",
			5470 => "0011111000110100000100",
			5471 => "0000000101010111110001",
			5472 => "0010000001010100000100",
			5473 => "0000000101010111110001",
			5474 => "0000000101010111110001",
			5475 => "0000000101010111110001",
			5476 => "0010010100101100001000",
			5477 => "0011111111101000000100",
			5478 => "0000000101010111110001",
			5479 => "0000000101010111110001",
			5480 => "0001101001111100001100",
			5481 => "0011000001011000001000",
			5482 => "0011001001110100000100",
			5483 => "0000000101010111110001",
			5484 => "0000001101010111110001",
			5485 => "0000000101010111110001",
			5486 => "0000000101010111110001",
			5487 => "0011000111010000010000",
			5488 => "0010101001000100000100",
			5489 => "0000000101010111110001",
			5490 => "0011110110001100000100",
			5491 => "0000000101010111110001",
			5492 => "0011101000011100000100",
			5493 => "0000000101010111110001",
			5494 => "0000000101010111110001",
			5495 => "0001100100101100001000",
			5496 => "0000011100011000000100",
			5497 => "0000000101010111110001",
			5498 => "0000000101010111110001",
			5499 => "0000000101010111110001",
			5500 => "0010011010100100100000",
			5501 => "0000101101101100000100",
			5502 => "1111111101011010110101",
			5503 => "0011101111101000011000",
			5504 => "0011000100011000000100",
			5505 => "1111111101011010110101",
			5506 => "0001001110111000001000",
			5507 => "0000010100110100000100",
			5508 => "1111111101011010110101",
			5509 => "0000000101011010110101",
			5510 => "0011001000000000000100",
			5511 => "0000001101011010110101",
			5512 => "0010010111101100000100",
			5513 => "1111111101011010110101",
			5514 => "0000001101011010110101",
			5515 => "1111111101011010110101",
			5516 => "0010110001001000011100",
			5517 => "0001000011110000010000",
			5518 => "0001100100111100001000",
			5519 => "0001010101110000000100",
			5520 => "1111111101011010110101",
			5521 => "0000001101011010110101",
			5522 => "0000011010011000000100",
			5523 => "1111111101011010110101",
			5524 => "0000000101011010110101",
			5525 => "0011100110111000000100",
			5526 => "0000001101011010110101",
			5527 => "0001011110010000000100",
			5528 => "1111111101011010110101",
			5529 => "0000000101011010110101",
			5530 => "0011001011011100100100",
			5531 => "0001101001111100011000",
			5532 => "0011011010000100010000",
			5533 => "0011000100000100001000",
			5534 => "0001011110110100000100",
			5535 => "0000001101011010110101",
			5536 => "0000001101011010110101",
			5537 => "0001010010000000000100",
			5538 => "0000000101011010110101",
			5539 => "0000001101011010110101",
			5540 => "0000100101000000000100",
			5541 => "1111111101011010110101",
			5542 => "0000001101011010110101",
			5543 => "0000011001100100000100",
			5544 => "1111111101011010110101",
			5545 => "0011001111011100000100",
			5546 => "0000000101011010110101",
			5547 => "0000001101011010110101",
			5548 => "0000000101011010110101",
			5549 => "0010011010100100101000",
			5550 => "0000101101101100000100",
			5551 => "1111111101011101110001",
			5552 => "0001100101010000100000",
			5553 => "0001001110111000001100",
			5554 => "0011001000011000000100",
			5555 => "1111111101011101110001",
			5556 => "0001110001011000000100",
			5557 => "0000000101011101110001",
			5558 => "0000000101011101110001",
			5559 => "0010011011001100000100",
			5560 => "1111111101011101110001",
			5561 => "0000101100001100001000",
			5562 => "0001111011000000000100",
			5563 => "0000000101011101110001",
			5564 => "0000010101011101110001",
			5565 => "0010010100101100000100",
			5566 => "1111111101011101110001",
			5567 => "0000001101011101110001",
			5568 => "1111111101011101110001",
			5569 => "0011001001110100001000",
			5570 => "0001010111111100000100",
			5571 => "1111111101011101110001",
			5572 => "0000000101011101110001",
			5573 => "0010100001010000011100",
			5574 => "0011011010000100010100",
			5575 => "0010110001001000001000",
			5576 => "0011100110111000000100",
			5577 => "0000001101011101110001",
			5578 => "0000000101011101110001",
			5579 => "0011010110111100000100",
			5580 => "0000001101011101110001",
			5581 => "0010111110101100000100",
			5582 => "0000000101011101110001",
			5583 => "0000001101011101110001",
			5584 => "0000000111000000000100",
			5585 => "1111111101011101110001",
			5586 => "0000001101011101110001",
			5587 => "0001000100001100001000",
			5588 => "0010010111110100000100",
			5589 => "1111111101011101110001",
			5590 => "0000001101011101110001",
			5591 => "0001100100101100001000",
			5592 => "0011100010111000000100",
			5593 => "0000001101011101110001",
			5594 => "0000000101011101110001",
			5595 => "1111111101011101110001",
			5596 => "0000101101101100001000",
			5597 => "0000110001011100000100",
			5598 => "1111111101100000011101",
			5599 => "0000000101100000011101",
			5600 => "0011111000000100100000",
			5601 => "0001100101010000010100",
			5602 => "0011001010111000000100",
			5603 => "0000000101100000011101",
			5604 => "0010011011001100000100",
			5605 => "0000000101100000011101",
			5606 => "0001000110111000000100",
			5607 => "0000000101100000011101",
			5608 => "0001101111000000000100",
			5609 => "0000000101100000011101",
			5610 => "0000001101100000011101",
			5611 => "0011111011110000001000",
			5612 => "0000010001111000000100",
			5613 => "0000000101100000011101",
			5614 => "0000000101100000011101",
			5615 => "0000000101100000011101",
			5616 => "0000011101011000101000",
			5617 => "0010110110100000011100",
			5618 => "0011101000011100010000",
			5619 => "0010010010101100001000",
			5620 => "0000101000110100000100",
			5621 => "1111111101100000011101",
			5622 => "0000000101100000011101",
			5623 => "0001010101110000000100",
			5624 => "0000000101100000011101",
			5625 => "0000001101100000011101",
			5626 => "0011010110111100001000",
			5627 => "0011000100000100000100",
			5628 => "1111111101100000011101",
			5629 => "0000000101100000011101",
			5630 => "0000000101100000011101",
			5631 => "0010010011101000001000",
			5632 => "0001001101001000000100",
			5633 => "0000000101100000011101",
			5634 => "1111111101100000011101",
			5635 => "1111111101100000011101",
			5636 => "0010000111000100000100",
			5637 => "0000001101100000011101",
			5638 => "0000000101100000011101",
			5639 => "0010011010100100100100",
			5640 => "0001100100111100000100",
			5641 => "1111111101100100010001",
			5642 => "0001101000010000001100",
			5643 => "0001001110111000000100",
			5644 => "1111111101100100010001",
			5645 => "0010011011001100000100",
			5646 => "0000000101100100010001",
			5647 => "0000001101100100010001",
			5648 => "0010010100101100000100",
			5649 => "1111111101100100010001",
			5650 => "0001000011101100001100",
			5651 => "0010010111101100001000",
			5652 => "0010010111101100000100",
			5653 => "0000000101100100010001",
			5654 => "0000000101100100010001",
			5655 => "1111111101100100010001",
			5656 => "0000001101100100010001",
			5657 => "0010110000110100101000",
			5658 => "0011100110111000010100",
			5659 => "0001001000001000010000",
			5660 => "0001010111111100001000",
			5661 => "0010000101000100000100",
			5662 => "0000000101100100010001",
			5663 => "1111111101100100010001",
			5664 => "0001101000010000000100",
			5665 => "0000001101100100010001",
			5666 => "0000000101100100010001",
			5667 => "0000001101100100010001",
			5668 => "0011001000011000010000",
			5669 => "0001000110001100000100",
			5670 => "1111110101100100010001",
			5671 => "0010100110011000000100",
			5672 => "0000000101100100010001",
			5673 => "0000000011111100000100",
			5674 => "1111111101100100010001",
			5675 => "0000000101100100010001",
			5676 => "0000001101100100010001",
			5677 => "0011010110111100010000",
			5678 => "0011000001011000001000",
			5679 => "0011100011110000000100",
			5680 => "0000001101100100010001",
			5681 => "0000000101100100010001",
			5682 => "0010110110100000000100",
			5683 => "0000000101100100010001",
			5684 => "0000000101100100010001",
			5685 => "0000101000110100010000",
			5686 => "0000110101000000001000",
			5687 => "0001001100001100000100",
			5688 => "0000001101100100010001",
			5689 => "0000000101100100010001",
			5690 => "0010101000010100000100",
			5691 => "1111110101100100010001",
			5692 => "0000001101100100010001",
			5693 => "0010001111001000001000",
			5694 => "0011101000000100000100",
			5695 => "0000000101100100010001",
			5696 => "0000001101100100010001",
			5697 => "0001000011011000000100",
			5698 => "1111111101100100010001",
			5699 => "0000000101100100010001",
			5700 => "0011001011000000000100",
			5701 => "1111111101100110111101",
			5702 => "0010110110100000111000",
			5703 => "0010010010101100100100",
			5704 => "0011100110111000010100",
			5705 => "0010010101010000000100",
			5706 => "0000000101100110111101",
			5707 => "0001000010110000001000",
			5708 => "0001110111010000000100",
			5709 => "0000000101100110111101",
			5710 => "0000000101100110111101",
			5711 => "0001100101010000000100",
			5712 => "0000001101100110111101",
			5713 => "0000000101100110111101",
			5714 => "0001101000010000000100",
			5715 => "0000000101100110111101",
			5716 => "0000011010011000001000",
			5717 => "0001011110110100000100",
			5718 => "1111111101100110111101",
			5719 => "0000000101100110111101",
			5720 => "0000000101100110111101",
			5721 => "0011000001101000001100",
			5722 => "0011001001110100000100",
			5723 => "0000000101100110111101",
			5724 => "0001110001011000000100",
			5725 => "0000000101100110111101",
			5726 => "0000000101100110111101",
			5727 => "0010011000010100000100",
			5728 => "0000001101100110111101",
			5729 => "0000000101100110111101",
			5730 => "0000011101011000010000",
			5731 => "0010010011101000001100",
			5732 => "0001100101010000001000",
			5733 => "0000011100011000000100",
			5734 => "0000000101100110111101",
			5735 => "0000000101100110111101",
			5736 => "0000000101100110111101",
			5737 => "1111111101100110111101",
			5738 => "0010000111000100001000",
			5739 => "0010110110100000000100",
			5740 => "0000000101100110111101",
			5741 => "0000000101100110111101",
			5742 => "0000000101100110111101",
			5743 => "0010010111101100001000",
			5744 => "0001000000100000000100",
			5745 => "1111111101101001101001",
			5746 => "0000000101101001101001",
			5747 => "0001100100111100001100",
			5748 => "0001110111010000001000",
			5749 => "0001000110001100000100",
			5750 => "0000000101101001101001",
			5751 => "0000000101101001101001",
			5752 => "0000000101101001101001",
			5753 => "0000000111000000011000",
			5754 => "0011111000011100001100",
			5755 => "0010110000110100001000",
			5756 => "0001110000011100000100",
			5757 => "0000000101101001101001",
			5758 => "0000000101101001101001",
			5759 => "0000000101101001101001",
			5760 => "0010010011101000000100",
			5761 => "0000000101101001101001",
			5762 => "0011010110111100000100",
			5763 => "0000000101101001101001",
			5764 => "1111111101101001101001",
			5765 => "0001100101010000010000",
			5766 => "0000101000000100000100",
			5767 => "0000000101101001101001",
			5768 => "0001111111011100000100",
			5769 => "0000000101101001101001",
			5770 => "0001110111110000000100",
			5771 => "0000001101101001101001",
			5772 => "0000000101101001101001",
			5773 => "0001000100001100001100",
			5774 => "0010011000100100001000",
			5775 => "0010100110011000000100",
			5776 => "0000000101101001101001",
			5777 => "0000000101101001101001",
			5778 => "0000000101101001101001",
			5779 => "0000000011010000001000",
			5780 => "0010011010100100000100",
			5781 => "0000000101101001101001",
			5782 => "0000000101101001101001",
			5783 => "0001001011001000000100",
			5784 => "0000000101101001101001",
			5785 => "0000000101101001101001",
			5786 => "0011001011000000000100",
			5787 => "1111111101101100011101",
			5788 => "0010110110100000111000",
			5789 => "0000100010110000101000",
			5790 => "0001001110100100010100",
			5791 => "0001110001011000001100",
			5792 => "0001101111000000000100",
			5793 => "0000000101101100011101",
			5794 => "0010110000110100000100",
			5795 => "1111111101101100011101",
			5796 => "0000000101101100011101",
			5797 => "0000010100110100000100",
			5798 => "0000000101101100011101",
			5799 => "0000001101101100011101",
			5800 => "0011000100000100001100",
			5801 => "0010010101010000000100",
			5802 => "0000000101101100011101",
			5803 => "0001111000011000000100",
			5804 => "0000000101101100011101",
			5805 => "0000001101101100011101",
			5806 => "0001010010000000000100",
			5807 => "0000000101101100011101",
			5808 => "0000000101101100011101",
			5809 => "0010010111110100001000",
			5810 => "0011000100000100000100",
			5811 => "1111111101101100011101",
			5812 => "0000000101101100011101",
			5813 => "0010101010110000000100",
			5814 => "0000000101101100011101",
			5815 => "0000000101101100011101",
			5816 => "0000011101011000010100",
			5817 => "0001101000010000000100",
			5818 => "0000000101101100011101",
			5819 => "0011001111011100000100",
			5820 => "0000000101101100011101",
			5821 => "0011101110100100001000",
			5822 => "0001010110010000000100",
			5823 => "0000000101101100011101",
			5824 => "1111111101101100011101",
			5825 => "0000000101101100011101",
			5826 => "0010100110011100001000",
			5827 => "0010110110100000000100",
			5828 => "0000000101101100011101",
			5829 => "0000000101101100011101",
			5830 => "0000000101101100011101",
			5831 => "0000101101101100001000",
			5832 => "0010111010010100000100",
			5833 => "1111111101101111101001",
			5834 => "0000000101101111101001",
			5835 => "0010010010101100111100",
			5836 => "0011100110111000011100",
			5837 => "0010011010100100010100",
			5838 => "0001000100001100001000",
			5839 => "0001100100111100000100",
			5840 => "0000000101101111101001",
			5841 => "1111111101101111101001",
			5842 => "0010100101000100001000",
			5843 => "0011000001101000000100",
			5844 => "0000001101101111101001",
			5845 => "0000000101101111101001",
			5846 => "0000000101101111101001",
			5847 => "0011011100010100000100",
			5848 => "0000000101101111101001",
			5849 => "0000001101101111101001",
			5850 => "0011001000011000010000",
			5851 => "0001000000010100001100",
			5852 => "0010111110101100001000",
			5853 => "0011111000110100000100",
			5854 => "0000000101101111101001",
			5855 => "1111111101101111101001",
			5856 => "0000000101101111101001",
			5857 => "0000000101101111101001",
			5858 => "0011000100000100001100",
			5859 => "0010101010110000001000",
			5860 => "0010011010100100000100",
			5861 => "0000000101101111101001",
			5862 => "0000001101101111101001",
			5863 => "0000000101101111101001",
			5864 => "1111111101101111101001",
			5865 => "0011000110100100001100",
			5866 => "0011001001110100001000",
			5867 => "0010001001101000000100",
			5868 => "0000000101101111101001",
			5869 => "0000000101101111101001",
			5870 => "1111111101101111101001",
			5871 => "0011010110111100000100",
			5872 => "0000001101101111101001",
			5873 => "0011000111010000001100",
			5874 => "0000110101000000000100",
			5875 => "0000000101101111101001",
			5876 => "0010000001010100000100",
			5877 => "1111111101101111101001",
			5878 => "0000000101101111101001",
			5879 => "0011001011011100000100",
			5880 => "0000001101101111101001",
			5881 => "0000000101101111101001",
			5882 => "0000010100110100011100",
			5883 => "0000101110000000000100",
			5884 => "1111111101110011000101",
			5885 => "0011111110100100010100",
			5886 => "0011001011000000000100",
			5887 => "1111111101110011000101",
			5888 => "0011001000011000001000",
			5889 => "0001001110111000000100",
			5890 => "0000000101110011000101",
			5891 => "0000001101110011000101",
			5892 => "0010110001001000000100",
			5893 => "0000000101110011000101",
			5894 => "1111111101110011000101",
			5895 => "1111111101110011000101",
			5896 => "0011001000011000101000",
			5897 => "0011100110001100100100",
			5898 => "0001000011110000010000",
			5899 => "0010110001001000001100",
			5900 => "0001100100111100001000",
			5901 => "0011101111100100000100",
			5902 => "0000000101110011000101",
			5903 => "0000000101110011000101",
			5904 => "1111111101110011000101",
			5905 => "0000001101110011000101",
			5906 => "0001100101010000001000",
			5907 => "0010110100010000000100",
			5908 => "0000000101110011000101",
			5909 => "0000001101110011000101",
			5910 => "0001001001001100001000",
			5911 => "0011111000110100000100",
			5912 => "0000000101110011000101",
			5913 => "0000000101110011000101",
			5914 => "0000000101110011000101",
			5915 => "1111111101110011000101",
			5916 => "0010110110100000010100",
			5917 => "0001101001111100010000",
			5918 => "0010110000110100001100",
			5919 => "0011101000011100001000",
			5920 => "0011001000011000000100",
			5921 => "0000000101110011000101",
			5922 => "0000001101110011000101",
			5923 => "1111111101110011000101",
			5924 => "0000001101110011000101",
			5925 => "0000000101110011000101",
			5926 => "0001110110110100000100",
			5927 => "1111101101110011000101",
			5928 => "0000001010101100001000",
			5929 => "0011111000011100000100",
			5930 => "0000000101110011000101",
			5931 => "1111111101110011000101",
			5932 => "0010101010110000000100",
			5933 => "0000001101110011000101",
			5934 => "0001000111011100000100",
			5935 => "1111111101110011000101",
			5936 => "0000000101110011000101",
			5937 => "0000101101101100001000",
			5938 => "0010111010010100000100",
			5939 => "1111111101110110011001",
			5940 => "0000000101110110011001",
			5941 => "0000011100011000111000",
			5942 => "0001100101010000101100",
			5943 => "0001001000001000010100",
			5944 => "0011001000011000001100",
			5945 => "0001100100111100000100",
			5946 => "0000000101110110011001",
			5947 => "0010000101000100000100",
			5948 => "0000000101110110011001",
			5949 => "1111111101110110011001",
			5950 => "0000010100110100000100",
			5951 => "0000000101110110011001",
			5952 => "0000000101110110011001",
			5953 => "0000010111101000001100",
			5954 => "0011110010010100001000",
			5955 => "0010011011001100000100",
			5956 => "0000000101110110011001",
			5957 => "0000001101110110011001",
			5958 => "1111111101110110011001",
			5959 => "0010110100010000000100",
			5960 => "0000000101110110011001",
			5961 => "0011010010000100000100",
			5962 => "0000001101110110011001",
			5963 => "0000000101110110011001",
			5964 => "0010110000110100001000",
			5965 => "0010111011110100000100",
			5966 => "1111111101110110011001",
			5967 => "0000000101110110011001",
			5968 => "1111111101110110011001",
			5969 => "0011000110100100010000",
			5970 => "0010010010101100001000",
			5971 => "0010010010101100000100",
			5972 => "0000000101110110011001",
			5973 => "0000000101110110011001",
			5974 => "0001010011001000000100",
			5975 => "1111111101110110011001",
			5976 => "0000000101110110011001",
			5977 => "0011010110111100001000",
			5978 => "0010110001001000000100",
			5979 => "0000000101110110011001",
			5980 => "0000001101110110011001",
			5981 => "0010111110101100000100",
			5982 => "1111111101110110011001",
			5983 => "0000011101011000001000",
			5984 => "0000011101011000000100",
			5985 => "0000000101110110011001",
			5986 => "1111111101110110011001",
			5987 => "0010000111000100000100",
			5988 => "0000001101110110011001",
			5989 => "0000000101110110011001",
			5990 => "0010010100111100000100",
			5991 => "1111111101111001001101",
			5992 => "0011100110111000100100",
			5993 => "0001001001000000100000",
			5994 => "0010011010100000001000",
			5995 => "0011111000011100000100",
			5996 => "0000000101111001001101",
			5997 => "0000000101111001001101",
			5998 => "0011110010010100001100",
			5999 => "0001101111000000000100",
			6000 => "0000000101111001001101",
			6001 => "0011000001101000000100",
			6002 => "0000000101111001001101",
			6003 => "0000000101111001001101",
			6004 => "0001100101010000001000",
			6005 => "0011011010001000000100",
			6006 => "0000000101111001001101",
			6007 => "0000000101111001001101",
			6008 => "0000000101111001001101",
			6009 => "0000000101111001001101",
			6010 => "0000011101011000101000",
			6011 => "0010111110101100010000",
			6012 => "0011111000110100000100",
			6013 => "0000000101111001001101",
			6014 => "0010011010100100000100",
			6015 => "0000000101111001001101",
			6016 => "0001100100111100000100",
			6017 => "0000000101111001001101",
			6018 => "1111111101111001001101",
			6019 => "0010010011101000001100",
			6020 => "0001001101001000001000",
			6021 => "0000010100110100000100",
			6022 => "0000000101111001001101",
			6023 => "0000000101111001001101",
			6024 => "0000000101111001001101",
			6025 => "0010111101000100001000",
			6026 => "0011111000011100000100",
			6027 => "0000000101111001001101",
			6028 => "0000000101111001001101",
			6029 => "0000000101111001001101",
			6030 => "0001100100101100001000",
			6031 => "0000111000000100000100",
			6032 => "0000000101111001001101",
			6033 => "0000000101111001001101",
			6034 => "0000000101111001001101",
			6035 => "0011001011000000000100",
			6036 => "1111111101111011100011",
			6037 => "0000011011111100000100",
			6038 => "1111111101111011100011",
			6039 => "0010110110100000101000",
			6040 => "0010110000110100011000",
			6041 => "0011101000011100010000",
			6042 => "0000101110000000001000",
			6043 => "0010110000110100000100",
			6044 => "0000000101111011100011",
			6045 => "0000001101111011100011",
			6046 => "0001101001111100000100",
			6047 => "0000001101111011100011",
			6048 => "1111111101111011100011",
			6049 => "0000011101011000000100",
			6050 => "1111111101111011100011",
			6051 => "0000001101111011100011",
			6052 => "0001101001111100001100",
			6053 => "0000010100110100001000",
			6054 => "0011110101000000000100",
			6055 => "0000000101111011100011",
			6056 => "0000000101111011100011",
			6057 => "0000001101111011100011",
			6058 => "1111111101111011100011",
			6059 => "0001110110110100000100",
			6060 => "1111110101111011100011",
			6061 => "0000001010101100001000",
			6062 => "0011111000011100000100",
			6063 => "0000000101111011100011",
			6064 => "1111111101111011100011",
			6065 => "0010101010110000001000",
			6066 => "0000011100011000000100",
			6067 => "0000000101111011100011",
			6068 => "0000001101111011100011",
			6069 => "0000011001100100000100",
			6070 => "1111111101111011100011",
			6071 => "0000000101111011100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1980, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(4056, initial_addr_3'length));
	end generate gen_rom_8;

	gen_rom_9: if SELECT_ROM = 9 generate
		bank <= (
			0 => "0011011110110000010100",
			1 => "0001000000101100000100",
			2 => "1111111000000010110101",
			3 => "0010001101010000001000",
			4 => "0010100001110000000100",
			5 => "0000000000000010110101",
			6 => "0000000000000010110101",
			7 => "0000101111010100000100",
			8 => "0000000000000010110101",
			9 => "0000000000000010110101",
			10 => "0011000100000000010000",
			11 => "0011110011001000001000",
			12 => "0001101011001100000100",
			13 => "0000000000000010110101",
			14 => "0000001000000010110101",
			15 => "0000010111100100000100",
			16 => "1111111000000010110101",
			17 => "0000000000000010110101",
			18 => "0011011011000000011000",
			19 => "0001000011011000010000",
			20 => "0001111000111100000100",
			21 => "0000000000000010110101",
			22 => "0010000110001000000100",
			23 => "0000000000000010110101",
			24 => "0011111101000100000100",
			25 => "0000000000000010110101",
			26 => "1111111000000010110101",
			27 => "0001101001100100000100",
			28 => "0000000000000010110101",
			29 => "0000000000000010110101",
			30 => "0001111000111000000100",
			31 => "0000001000000010110101",
			32 => "0010110110000100001100",
			33 => "0001101001100100001000",
			34 => "0000101100010000000100",
			35 => "0000001000000010110101",
			36 => "1111111000000010110101",
			37 => "0000001000000010110101",
			38 => "0000011011101000001000",
			39 => "0011000011011100000100",
			40 => "0000000000000010110101",
			41 => "1111111000000010110101",
			42 => "0010111001110100000100",
			43 => "0000001000000010110101",
			44 => "0000000000000010110101",
			45 => "0001011010111100010100",
			46 => "0000101100000000001000",
			47 => "0011011010111000000100",
			48 => "1111111000000101101001",
			49 => "0000000000000101101001",
			50 => "0011010001111100000100",
			51 => "0000000000000101101001",
			52 => "0000001100001000000100",
			53 => "0000000000000101101001",
			54 => "0000000000000101101001",
			55 => "0011011101101101000100",
			56 => "0011000000101000010100",
			57 => "0001111000111000001100",
			58 => "0010111101100000001000",
			59 => "0000000010011000000100",
			60 => "0000000000000101101001",
			61 => "0000000000000101101001",
			62 => "0000000000000101101001",
			63 => "0001101011001100000100",
			64 => "0000000000000101101001",
			65 => "0000001000000101101001",
			66 => "0000110010000000100000",
			67 => "0000000010011000010000",
			68 => "0000101001100000001000",
			69 => "0000110111110000000100",
			70 => "0000000000000101101001",
			71 => "0000000000000101101001",
			72 => "0011000100000000000100",
			73 => "0000000000000101101001",
			74 => "1111111000000101101001",
			75 => "0000101100000000001000",
			76 => "0000111111011100000100",
			77 => "0000000000000101101001",
			78 => "0000000000000101101001",
			79 => "0001101111000000000100",
			80 => "1111111000000101101001",
			81 => "0000000000000101101001",
			82 => "0001110001111100000100",
			83 => "0000001000000101101001",
			84 => "0000110010000100000100",
			85 => "1111111000000101101001",
			86 => "0001010111100000000100",
			87 => "0000000000000101101001",
			88 => "0000000000000101101001",
			89 => "1111111000000101101001",
			90 => "0000010110101001000000",
			91 => "0001000011011000101000",
			92 => "0011001000111000011100",
			93 => "0000110000011100001100",
			94 => "0011000100010100000100",
			95 => "0000000000001010001101",
			96 => "0001000111011100000100",
			97 => "0000000000001010001101",
			98 => "0000000000001010001101",
			99 => "0011110111111100000100",
			100 => "0000000000001010001101",
			101 => "0001000010111000000100",
			102 => "1111111000001010001101",
			103 => "0011111110010000000100",
			104 => "0000000000001010001101",
			105 => "0000000000001010001101",
			106 => "0011000011011100001000",
			107 => "0001111000111000000100",
			108 => "0000000000001010001101",
			109 => "1111111000001010001101",
			110 => "0000000000001010001101",
			111 => "0010001111000100001000",
			112 => "0001101011001100000100",
			113 => "0000000000001010001101",
			114 => "0000001000001010001101",
			115 => "0001000110110000000100",
			116 => "0000000000001010001101",
			117 => "0011110100010000000100",
			118 => "0000000000001010001101",
			119 => "0000101111100100000100",
			120 => "0000000000001010001101",
			121 => "0000000000001010001101",
			122 => "0011100101110100010100",
			123 => "0001000101010100001100",
			124 => "0000111011011100000100",
			125 => "0000000000001010001101",
			126 => "0001101010011000000100",
			127 => "0000000000001010001101",
			128 => "0000001000001010001101",
			129 => "0001100100111100000100",
			130 => "0000000000001010001101",
			131 => "0000000000001010001101",
			132 => "0010011110010100001100",
			133 => "0001101000010000001000",
			134 => "0001000010010100000100",
			135 => "0000000000001010001101",
			136 => "0000000000001010001101",
			137 => "0000000000001010001101",
			138 => "0010011101111100010100",
			139 => "0011110010000000001000",
			140 => "0010110000001100000100",
			141 => "0000000000001010001101",
			142 => "0000000000001010001101",
			143 => "0011100111111100001000",
			144 => "0001000110111000000100",
			145 => "0000000000001010001101",
			146 => "0000001000001010001101",
			147 => "0000000000001010001101",
			148 => "0011111011110000010000",
			149 => "0010000001010100001000",
			150 => "0001010010011100000100",
			151 => "0000000000001010001101",
			152 => "0000000000001010001101",
			153 => "0001100101010000000100",
			154 => "0000000000001010001101",
			155 => "0000000000001010001101",
			156 => "0000111110000000001000",
			157 => "0000000111000000000100",
			158 => "0000000000001010001101",
			159 => "0000000000001010001101",
			160 => "0001100100101100000100",
			161 => "0000000000001010001101",
			162 => "0000000000001010001101",
			163 => "0000010110101001000100",
			164 => "0010100101000100100100",
			165 => "0011000000101000001000",
			166 => "0011011110110000000100",
			167 => "0000000000001110110001",
			168 => "0000000000001110110001",
			169 => "0011011000000000001000",
			170 => "0001110100000000000100",
			171 => "0000000000001110110001",
			172 => "1111111000001110110001",
			173 => "0011100101100100010000",
			174 => "0011001000111000001000",
			175 => "0001111001110000000100",
			176 => "0000000000001110110001",
			177 => "0000000000001110110001",
			178 => "0000101100000000000100",
			179 => "0000000000001110110001",
			180 => "0000000000001110110001",
			181 => "1111111000001110110001",
			182 => "0010001111000100010000",
			183 => "0001001001000000000100",
			184 => "0000000000001110110001",
			185 => "0000111101010100000100",
			186 => "0000000000001110110001",
			187 => "0011010111001000000100",
			188 => "0000000000001110110001",
			189 => "0000000000001110110001",
			190 => "0001000110110000000100",
			191 => "0000000000001110110001",
			192 => "0011110100010000000100",
			193 => "0000000000001110110001",
			194 => "0000101111100100000100",
			195 => "0000000000001110110001",
			196 => "0000000000001110110001",
			197 => "0011100101110100010100",
			198 => "0001000101010100001100",
			199 => "0000111011011100000100",
			200 => "0000000000001110110001",
			201 => "0000000001110000000100",
			202 => "0000000000001110110001",
			203 => "0000001000001110110001",
			204 => "0010100110011100000100",
			205 => "0000000000001110110001",
			206 => "0000000000001110110001",
			207 => "0010011011111100001000",
			208 => "0011110110010000000100",
			209 => "0000000000001110110001",
			210 => "0000000000001110110001",
			211 => "0010111101000100100000",
			212 => "0000101000110100010000",
			213 => "0000100011000000001000",
			214 => "0010000110001000000100",
			215 => "0000000000001110110001",
			216 => "0000000000001110110001",
			217 => "0010010111101100000100",
			218 => "0000000000001110110001",
			219 => "0000000000001110110001",
			220 => "0010000010101000001000",
			221 => "0011001001001000000100",
			222 => "0000001000001110110001",
			223 => "0000000000001110110001",
			224 => "0000010000111100000100",
			225 => "0000000000001110110001",
			226 => "0000000000001110110001",
			227 => "0010010111101100001000",
			228 => "0000000011010000000100",
			229 => "0000000000001110110001",
			230 => "0000000000001110110001",
			231 => "0000001010101100000100",
			232 => "0000000000001110110001",
			233 => "0010011001000100000100",
			234 => "1111111000001110110001",
			235 => "0000000000001110110001",
			236 => "0011011110110000010100",
			237 => "0001000000101100000100",
			238 => "1111111000010010011101",
			239 => "0000000011011100001000",
			240 => "0010100001010100000100",
			241 => "0000000000010010011101",
			242 => "0000000000010010011101",
			243 => "0010101111001000000100",
			244 => "0000000000010010011101",
			245 => "0000000000010010011101",
			246 => "0001100100101101010100",
			247 => "0011111000110100101000",
			248 => "0011000100000000010000",
			249 => "0011110011001000001000",
			250 => "0001101011001100000100",
			251 => "0000000000010010011101",
			252 => "0000001000010010011101",
			253 => "0010111100101100000100",
			254 => "1111111000010010011101",
			255 => "0000000000010010011101",
			256 => "0011000100000000001000",
			257 => "0000010111100100000100",
			258 => "1111111000010010011101",
			259 => "0000000000010010011101",
			260 => "0001010111100000001000",
			261 => "0001000110111000000100",
			262 => "0000000000010010011101",
			263 => "0000000000010010011101",
			264 => "0011011100010100000100",
			265 => "0000000000010010011101",
			266 => "0000000000010010011101",
			267 => "0001000100001100011000",
			268 => "0000011101011000001100",
			269 => "0010000001010100000100",
			270 => "0000000000010010011101",
			271 => "0000001010101100000100",
			272 => "0000000000010010011101",
			273 => "0000001000010010011101",
			274 => "0000001010101100000100",
			275 => "0000000000010010011101",
			276 => "0001010011001000000100",
			277 => "0000000000010010011101",
			278 => "0000000000010010011101",
			279 => "0001011110010000000100",
			280 => "1111111000010010011101",
			281 => "0011001111011100001000",
			282 => "0000111110100100000100",
			283 => "0000000000010010011101",
			284 => "0000001000010010011101",
			285 => "0010101010110000000100",
			286 => "0000000000010010011101",
			287 => "0000000000010010011101",
			288 => "0011100011110000000100",
			289 => "0000000000010010011101",
			290 => "0011101011100000000100",
			291 => "1111111000010010011101",
			292 => "0001101010100000000100",
			293 => "0000000000010010011101",
			294 => "0000000000010010011101",
			295 => "0011111001010001000000",
			296 => "0000111001110100011100",
			297 => "0001000010010000001000",
			298 => "0011011000011000000100",
			299 => "0000000000010110110001",
			300 => "0000000000010110110001",
			301 => "0010111000111100000100",
			302 => "0000000000010110110001",
			303 => "0000100010000100000100",
			304 => "0000000000010110110001",
			305 => "0000101000100000001000",
			306 => "0010111100101100000100",
			307 => "0000000000010110110001",
			308 => "0000000000010110110001",
			309 => "0000000000010110110001",
			310 => "0001101011001100011000",
			311 => "0011000100000000001000",
			312 => "0010011011101000000100",
			313 => "0000000000010110110001",
			314 => "0000000000010110110001",
			315 => "0011000100000000001000",
			316 => "0011010011100000000100",
			317 => "0000000000010110110001",
			318 => "0000000000010110110001",
			319 => "0010010001111000000100",
			320 => "0000000000010110110001",
			321 => "0000000000010110110001",
			322 => "0000100010000000000100",
			323 => "0000000000010110110001",
			324 => "0011011001001000000100",
			325 => "0000001000010110110001",
			326 => "0000000000010110110001",
			327 => "0000110001011000000100",
			328 => "1111111000010110110001",
			329 => "0010000001110100110000",
			330 => "0000000000111000100000",
			331 => "0000011001011000010000",
			332 => "0011001001110000001000",
			333 => "0001101001100100000100",
			334 => "0000000000010110110001",
			335 => "0000000000010110110001",
			336 => "0001001110111000000100",
			337 => "1111111000010110110001",
			338 => "0000000000010110110001",
			339 => "0000010101011100001000",
			340 => "0001101010011000000100",
			341 => "0000000000010110110001",
			342 => "0000001000010110110001",
			343 => "0011111110000000000100",
			344 => "0000000000010110110001",
			345 => "0000000000010110110001",
			346 => "0000000000110000001000",
			347 => "0011001100110000000100",
			348 => "0000001000010110110001",
			349 => "0000000000010110110001",
			350 => "0010101100011100000100",
			351 => "0000000000010110110001",
			352 => "0000000000010110110001",
			353 => "0010100101000100001000",
			354 => "0011100101100100000100",
			355 => "0000000000010110110001",
			356 => "1111111000010110110001",
			357 => "0010001111000100001100",
			358 => "0011000011011100000100",
			359 => "0000000000010110110001",
			360 => "0010011010100100000100",
			361 => "0000000000010110110001",
			362 => "0000000000010110110001",
			363 => "0000000000010110110001",
			364 => "0001101010011000100100",
			365 => "0000010101011100010000",
			366 => "0010101010100000001100",
			367 => "0000001100000100000100",
			368 => "1111111000011011001101",
			369 => "0011101100110000000100",
			370 => "0000000000011011001101",
			371 => "0000001000011011001101",
			372 => "1111111000011011001101",
			373 => "0001101010011000001100",
			374 => "0011010010011100001000",
			375 => "0001110110100100000100",
			376 => "1111111000011011001101",
			377 => "0000001000011011001101",
			378 => "0000010000011011001101",
			379 => "0010010100101100000100",
			380 => "1111111000011011001101",
			381 => "0000000000011011001101",
			382 => "0010101001101001011100",
			383 => "0001101000010000111000",
			384 => "0001000011000000011000",
			385 => "0000001111001000001100",
			386 => "0010100011101000001000",
			387 => "0000011101111100000100",
			388 => "0000000000011011001101",
			389 => "0000011000011011001101",
			390 => "1111111000011011001101",
			391 => "0000100000010000001000",
			392 => "0011000100011000000100",
			393 => "0000001000011011001101",
			394 => "0000010000011011001101",
			395 => "1111111000011011001101",
			396 => "0011001000111100010000",
			397 => "0011011110110000001000",
			398 => "0001001100111100000100",
			399 => "1111111000011011001101",
			400 => "0000001000011011001101",
			401 => "0000000011010000000100",
			402 => "0000000000011011001101",
			403 => "0000001000011011001101",
			404 => "0000111011011100001000",
			405 => "0001000011010100000100",
			406 => "1111111000011011001101",
			407 => "0000000000011011001101",
			408 => "0001110101101100000100",
			409 => "0000001000011011001101",
			410 => "0000000000011011001101",
			411 => "0001111111011100010100",
			412 => "0001000111011100001100",
			413 => "0001000011110100001000",
			414 => "0000010101011100000100",
			415 => "0000000000011011001101",
			416 => "0000001000011011001101",
			417 => "0000001000011011001101",
			418 => "0000011101011100000100",
			419 => "0000001000011011001101",
			420 => "1111111000011011001101",
			421 => "0010100110011000000100",
			422 => "1111111000011011001101",
			423 => "0000111011110000000100",
			424 => "1111111000011011001101",
			425 => "0001100101010000000100",
			426 => "0000001000011011001101",
			427 => "0000000000011011001101",
			428 => "0011000100000000000100",
			429 => "0000000000011011001101",
			430 => "0000000110000100000100",
			431 => "1111110000011011001101",
			432 => "0000001100101100000100",
			433 => "0000000000011011001101",
			434 => "1111111000011011001101",
			435 => "0000110111110001001000",
			436 => "0010111100101100111000",
			437 => "0011100010001000110000",
			438 => "0011011000000000100000",
			439 => "0001111000111000010000",
			440 => "0001011101010100001000",
			441 => "0000101100000000000100",
			442 => "0000000000011111110001",
			443 => "0000000000011111110001",
			444 => "0000100010000100000100",
			445 => "0000000000011111110001",
			446 => "0000000000011111110001",
			447 => "0001001110111000001000",
			448 => "0010111100101100000100",
			449 => "1111111000011111110001",
			450 => "0000000000011111110001",
			451 => "0000001010000000000100",
			452 => "0000000000011111110001",
			453 => "0000000000011111110001",
			454 => "0001101001100100001100",
			455 => "0010011001011000001000",
			456 => "0000100010000100000100",
			457 => "0000000000011111110001",
			458 => "0000000000011111110001",
			459 => "0000000000011111110001",
			460 => "0000001000011111110001",
			461 => "0000110101110100000100",
			462 => "1111111000011111110001",
			463 => "0000000000011111110001",
			464 => "0001101111000000001000",
			465 => "0000100001000000000100",
			466 => "0000000000011111110001",
			467 => "1111111000011111110001",
			468 => "0011010001101000000100",
			469 => "0000000000011111110001",
			470 => "0000000000011111110001",
			471 => "0001010100000100010100",
			472 => "0000001000101100000100",
			473 => "0000000000011111110001",
			474 => "0010011011111100001100",
			475 => "0010111110001100000100",
			476 => "0000000000011111110001",
			477 => "0001001010110100000100",
			478 => "0000000000011111110001",
			479 => "0000000000011111110001",
			480 => "0000001000011111110001",
			481 => "0010011100011000001100",
			482 => "0000110010000000000100",
			483 => "1111111000011111110001",
			484 => "0010010001111000000100",
			485 => "0000000000011111110001",
			486 => "0000000000011111110001",
			487 => "0001010000110100010100",
			488 => "0001001100111100010000",
			489 => "0010011000010000001000",
			490 => "0011101110101100000100",
			491 => "0000000000011111110001",
			492 => "0000001000011111110001",
			493 => "0001100100111100000100",
			494 => "0000000000011111110001",
			495 => "0000000000011111110001",
			496 => "0000000000011111110001",
			497 => "0011011110101000001000",
			498 => "0010010000001000000100",
			499 => "1111111000011111110001",
			500 => "0000000000011111110001",
			501 => "0011011111010000001000",
			502 => "0011101100000000000100",
			503 => "0000000000011111110001",
			504 => "0000000000011111110001",
			505 => "0000110110111000000100",
			506 => "0000000000011111110001",
			507 => "0000000000011111110001",
			508 => "0001101101011000101100",
			509 => "0000010001000100010100",
			510 => "0010001001000100010000",
			511 => "0001010110110100001100",
			512 => "0010000011101000000100",
			513 => "1111111000100100110101",
			514 => "0001011100101100000100",
			515 => "0000000000100100110101",
			516 => "0000001000100100110101",
			517 => "1111111000100100110101",
			518 => "1111111000100100110101",
			519 => "0000111111010100010000",
			520 => "0000100111011000001100",
			521 => "0001000111011000000100",
			522 => "0000001000100100110101",
			523 => "0011111100000000000100",
			524 => "1111111000100100110101",
			525 => "0000000000100100110101",
			526 => "0000001000100100110101",
			527 => "0000100110111100000100",
			528 => "0000000000100100110101",
			529 => "1111111000100100110101",
			530 => "0011001000011001010100",
			531 => "0001101000010000110000",
			532 => "0001001000000100011100",
			533 => "0011001001110000001100",
			534 => "0001101011001100000100",
			535 => "1111111000100100110101",
			536 => "0011001000111000000100",
			537 => "0000001000100100110101",
			538 => "0000001000100100110101",
			539 => "0011010001000000001000",
			540 => "0001001100111000000100",
			541 => "0000000000100100110101",
			542 => "1111111000100100110101",
			543 => "0011010101110000000100",
			544 => "0000001000100100110101",
			545 => "0000000000100100110101",
			546 => "0001101011001100000100",
			547 => "1111111000100100110101",
			548 => "0011000100000000001000",
			549 => "0010111000111100000100",
			550 => "1111111000100100110101",
			551 => "0000001000100100110101",
			552 => "0000111000011000000100",
			553 => "1111111000100100110101",
			554 => "0000000000100100110101",
			555 => "0010100001010100011100",
			556 => "0001010101110000010000",
			557 => "0010011001111100001000",
			558 => "0010000111000100000100",
			559 => "0000000000100100110101",
			560 => "0000001000100100110101",
			561 => "0010001100000100000100",
			562 => "0000000000100100110101",
			563 => "0000001000100100110101",
			564 => "0011111101001000001000",
			565 => "0011001000011000000100",
			566 => "1111111000100100110101",
			567 => "0000001000100100110101",
			568 => "0000001000100100110101",
			569 => "0001100101010000000100",
			570 => "0000001000100100110101",
			571 => "1111111000100100110101",
			572 => "0011010110111100001100",
			573 => "0000010101011100001000",
			574 => "0001010010000000000100",
			575 => "0000000000100100110101",
			576 => "0000001000100100110101",
			577 => "1111111000100100110101",
			578 => "0010001000101100010100",
			579 => "0000101000110100001000",
			580 => "0011111000011100000100",
			581 => "0000000000100100110101",
			582 => "0000011000100100110101",
			583 => "0011011111010100000100",
			584 => "1111111000100100110101",
			585 => "0010010111101100000100",
			586 => "0000001000100100110101",
			587 => "0000000000100100110101",
			588 => "1111111000100100110101",
			589 => "0001011010111000011000",
			590 => "0001001111100000000100",
			591 => "1111111000101001001001",
			592 => "0011010001111100000100",
			593 => "1111111000101001001001",
			594 => "0011111110000100001100",
			595 => "0001101011001100001000",
			596 => "0011000000101000000100",
			597 => "0000000000101001001001",
			598 => "0000000000101001001001",
			599 => "0000001000101001001001",
			600 => "1111111000101001001001",
			601 => "0001010100011000011100",
			602 => "0011011011000000010100",
			603 => "0010110101101100001000",
			604 => "0000011001111000000100",
			605 => "0000000000101001001001",
			606 => "1111111000101001001001",
			607 => "0001101101011000000100",
			608 => "0000000000101001001001",
			609 => "0000100010000100000100",
			610 => "0000001000101001001001",
			611 => "0000000000101001001001",
			612 => "0001101101011000000100",
			613 => "0000000000101001001001",
			614 => "0000001000101001001001",
			615 => "0011011000000000011100",
			616 => "0001000010100100010000",
			617 => "0011110101110000001100",
			618 => "0000010110101000001000",
			619 => "0000001010000000000100",
			620 => "1111111000101001001001",
			621 => "0000000000101001001001",
			622 => "0000000000101001001001",
			623 => "1111111000101001001001",
			624 => "0000100111010100001000",
			625 => "0011001100110000000100",
			626 => "0000001000101001001001",
			627 => "0000000000101001001001",
			628 => "0000000000101001001001",
			629 => "0010111100101100011100",
			630 => "0011111001011100010000",
			631 => "0000001111000100001000",
			632 => "0001010011100000000100",
			633 => "0000000000101001001001",
			634 => "0000000000101001001001",
			635 => "0001010011100000000100",
			636 => "0000001000101001001001",
			637 => "0000000000101001001001",
			638 => "0001101001100100000100",
			639 => "1111111000101001001001",
			640 => "0000101111010100000100",
			641 => "0000001000101001001001",
			642 => "0000000000101001001001",
			643 => "0011100101100100010000",
			644 => "0000000001110100001000",
			645 => "0011000110000100000100",
			646 => "0000000000101001001001",
			647 => "0000000000101001001001",
			648 => "0001101111000000000100",
			649 => "1111111000101001001001",
			650 => "0000000000101001001001",
			651 => "0001011001001000001000",
			652 => "0010100001010000000100",
			653 => "0000000000101001001001",
			654 => "0000001000101001001001",
			655 => "0010010100110100000100",
			656 => "0000000000101001001001",
			657 => "0000000000101001001001",
			658 => "0001101010011000100100",
			659 => "0000010101011100010000",
			660 => "0010101010100000001100",
			661 => "0000001100000100000100",
			662 => "1111111000101110000101",
			663 => "0011101100110000000100",
			664 => "0000000000101110000101",
			665 => "0000001000101110000101",
			666 => "1111111000101110000101",
			667 => "0001101010011000001100",
			668 => "0011010010011100001000",
			669 => "0001110110100100000100",
			670 => "1111111000101110000101",
			671 => "0000001000101110000101",
			672 => "0000010000101110000101",
			673 => "0010010100101100000100",
			674 => "1111111000101110000101",
			675 => "0000000000101110000101",
			676 => "0011001000011001010100",
			677 => "0001101000010000110000",
			678 => "0000111001110100010000",
			679 => "0001101001100100000100",
			680 => "1111111000101110000101",
			681 => "0001111101100000001000",
			682 => "0011010111001000000100",
			683 => "0000000000101110000101",
			684 => "0000001000101110000101",
			685 => "1111111000101110000101",
			686 => "0011001000111100010000",
			687 => "0001101001100100001000",
			688 => "0010011101011100000100",
			689 => "0000001000101110000101",
			690 => "0000000000101110000101",
			691 => "0000110000011100000100",
			692 => "0000000000101110000101",
			693 => "0000001000101110000101",
			694 => "0000111011011100001000",
			695 => "0001000011010100000100",
			696 => "1111111000101110000101",
			697 => "0000000000101110000101",
			698 => "0010110000001100000100",
			699 => "0000001000101110000101",
			700 => "0000000000101110000101",
			701 => "0001000111011100011000",
			702 => "0010111011110100001100",
			703 => "0010101001000100000100",
			704 => "0000000000101110000101",
			705 => "0010011010011000000100",
			706 => "0000000000101110000101",
			707 => "0000001000101110000101",
			708 => "0010010010101100000100",
			709 => "1111111000101110000101",
			710 => "0000011101011000000100",
			711 => "0000001000101110000101",
			712 => "0000000000101110000101",
			713 => "0010011110010100000100",
			714 => "0000001000101110000101",
			715 => "0001001101110100000100",
			716 => "0000000000101110000101",
			717 => "1111111000101110000101",
			718 => "0011010110111100001000",
			719 => "0001101111000000000100",
			720 => "0000000000101110000101",
			721 => "1111111000101110000101",
			722 => "0001111011011100000100",
			723 => "0001001000101110000101",
			724 => "0011101110100100010000",
			725 => "0010110110100000001000",
			726 => "0011100110111000000100",
			727 => "0000000000101110000101",
			728 => "1111111000101110000101",
			729 => "0010010011101000000100",
			730 => "0000001000101110000101",
			731 => "0000010000101110000101",
			732 => "0000001011000100001000",
			733 => "0010111111010000000100",
			734 => "1111111000101110000101",
			735 => "0000000000101110000101",
			736 => "1111111000101110000101",
			737 => "0001010111001000011000",
			738 => "0001000001101100000100",
			739 => "1111111000110010111001",
			740 => "0010110011011100010000",
			741 => "0000100111011000000100",
			742 => "0000000000110010111001",
			743 => "0000100000010000001000",
			744 => "0001010011011100000100",
			745 => "0000000000110010111001",
			746 => "0000000000110010111001",
			747 => "0000000000110010111001",
			748 => "0000000000110010111001",
			749 => "0011111111010000111100",
			750 => "0001111001110000011100",
			751 => "0010101010110000001100",
			752 => "0011000100000000000100",
			753 => "1111111000110010111001",
			754 => "0011000100000000000100",
			755 => "0000001000110010111001",
			756 => "0000000000110010111001",
			757 => "0011100100001000000100",
			758 => "0000000000110010111001",
			759 => "0001101101011000000100",
			760 => "0000000000110010111001",
			761 => "0011000100000000000100",
			762 => "0000001000110010111001",
			763 => "0000000000110010111001",
			764 => "0011101011011100011000",
			765 => "0011111110000100001100",
			766 => "0010110110000100000100",
			767 => "0000000000110010111001",
			768 => "0000100001000000000100",
			769 => "0000000000110010111001",
			770 => "1111111000110010111001",
			771 => "0000000100010100000100",
			772 => "0000000000110010111001",
			773 => "0010110000001100000100",
			774 => "0000000000110010111001",
			775 => "0000000000110010111001",
			776 => "0001100111101000000100",
			777 => "0000000000110010111001",
			778 => "0000001000110010111001",
			779 => "0000010110101000100100",
			780 => "0011110111111100010100",
			781 => "0001111001110000001000",
			782 => "0001101011001100000100",
			783 => "0000000000110010111001",
			784 => "0000001000110010111001",
			785 => "0000000011010000000100",
			786 => "1111111000110010111001",
			787 => "0010100110011100000100",
			788 => "0000000000110010111001",
			789 => "0000000000110010111001",
			790 => "0011001000111000001100",
			791 => "0001000010111000000100",
			792 => "1111111000110010111001",
			793 => "0000001010000000000100",
			794 => "0000000000110010111001",
			795 => "1111111000110010111001",
			796 => "0000000000110010111001",
			797 => "0001011000000000001100",
			798 => "0011011001110100001000",
			799 => "0011000100000000000100",
			800 => "0000000000110010111001",
			801 => "0000000000110010111001",
			802 => "0000001000110010111001",
			803 => "0010010111101000001100",
			804 => "0011010110100100000100",
			805 => "0000000000110010111001",
			806 => "0000101010000100000100",
			807 => "1111111000110010111001",
			808 => "0000000000110010111001",
			809 => "0001011000011000000100",
			810 => "0000001000110010111001",
			811 => "0011011011101100000100",
			812 => "0000000000110010111001",
			813 => "1111111000110010111001",
			814 => "0010110011011100001100",
			815 => "0000101111010100000100",
			816 => "1111111000110110001101",
			817 => "0000001100110000000100",
			818 => "0000000000110110001101",
			819 => "0000001000110110001101",
			820 => "0010101001101001011000",
			821 => "0000010111100100110100",
			822 => "0000000010011000011000",
			823 => "0001111001110000001000",
			824 => "0000001111000100000100",
			825 => "1111111000110110001101",
			826 => "1111101000110110001101",
			827 => "0011001000111100001000",
			828 => "0010101001000100000100",
			829 => "0000000000110110001101",
			830 => "0000001000110110001101",
			831 => "0011000110000100000100",
			832 => "1111111000110110001101",
			833 => "0000001000110110001101",
			834 => "0001000010100100010000",
			835 => "0010111110001100001000",
			836 => "0000110000011100000100",
			837 => "0000000000110110001101",
			838 => "0000000000110110001101",
			839 => "0010111101111000000100",
			840 => "1111110000110110001101",
			841 => "1111111000110110001101",
			842 => "0011000011011100001000",
			843 => "0000111010001100000100",
			844 => "0000000000110110001101",
			845 => "0000001000110110001101",
			846 => "1111111000110110001101",
			847 => "0001010001101000000100",
			848 => "0000001000110110001101",
			849 => "0010011100011000010000",
			850 => "0001110001111100001000",
			851 => "0010100110011100000100",
			852 => "1111111000110110001101",
			853 => "0000000000110110001101",
			854 => "0001001110000000000100",
			855 => "0000001000110110001101",
			856 => "1111111000110110001101",
			857 => "0010100010101100001000",
			858 => "0010010101010000000100",
			859 => "0000000000110110001101",
			860 => "0000001000110110001101",
			861 => "0011111000110100000100",
			862 => "0000000000110110001101",
			863 => "0000000000110110001101",
			864 => "0011001000111100000100",
			865 => "0000001000110110001101",
			866 => "1111111000110110001101",
			867 => "0001000011000000111000",
			868 => "0010110000011100011000",
			869 => "0010101001000100010100",
			870 => "0010001010110000001100",
			871 => "0001001011101100001000",
			872 => "0000000110001000000100",
			873 => "0000000000111011011001",
			874 => "0000000000111011011001",
			875 => "0000000000111011011001",
			876 => "0001000000010000000100",
			877 => "0000000000111011011001",
			878 => "1111111000111011011001",
			879 => "0000000000111011011001",
			880 => "0001110001101000010100",
			881 => "0010011010100000010000",
			882 => "0000010101011100000100",
			883 => "0000000000111011011001",
			884 => "0001111001001000000100",
			885 => "0000000000111011011001",
			886 => "0001010111100000000100",
			887 => "0000001000111011011001",
			888 => "0000000000111011011001",
			889 => "0000000000111011011001",
			890 => "0001101101011000001000",
			891 => "0001101101011000000100",
			892 => "0000000000111011011001",
			893 => "0000000000111011011001",
			894 => "0000000000111011011001",
			895 => "0001000110001100111100",
			896 => "0000010111100100011000",
			897 => "0000000010011000000100",
			898 => "1111111000111011011001",
			899 => "0001010100011000001100",
			900 => "0010001011010100000100",
			901 => "0000000000111011011001",
			902 => "0000000011111100000100",
			903 => "1111111000111011011001",
			904 => "0000000000111011011001",
			905 => "0001111101100000000100",
			906 => "0000000000111011011001",
			907 => "0000000000111011011001",
			908 => "0010110000001100000100",
			909 => "0000001000111011011001",
			910 => "0000000111000000010000",
			911 => "0000001010101100001000",
			912 => "0001001000000100000100",
			913 => "0000000000111011011001",
			914 => "0000000000111011011001",
			915 => "0001100100111100000100",
			916 => "0000000000111011011001",
			917 => "0000000000111011011001",
			918 => "0010010111101100001000",
			919 => "0001001000110100000100",
			920 => "0000000000111011011001",
			921 => "1111111000111011011001",
			922 => "0010110100010000000100",
			923 => "0000000000111011011001",
			924 => "0000000000111011011001",
			925 => "0001101101011000000100",
			926 => "1111111000111011011001",
			927 => "0001111000111000010100",
			928 => "0001011101010100001100",
			929 => "0010111000111100000100",
			930 => "0000000000111011011001",
			931 => "0001000011011000000100",
			932 => "0000000000111011011001",
			933 => "0000000000111011011001",
			934 => "0011010011100000000100",
			935 => "0000000000111011011001",
			936 => "0000001000111011011001",
			937 => "0010000111000000010000",
			938 => "0001001101001000001000",
			939 => "0010000111000100000100",
			940 => "0000000000111011011001",
			941 => "1111111000111011011001",
			942 => "0000111010011100000100",
			943 => "0000000000111011011001",
			944 => "0000000000111011011001",
			945 => "0011100100001000001000",
			946 => "0011011110110000000100",
			947 => "0000000000111011011001",
			948 => "0000000000111011011001",
			949 => "1111111000111011011001",
			950 => "0001101010011000101000",
			951 => "0000010101011100010100",
			952 => "0010101010100000010000",
			953 => "0010001000010100001100",
			954 => "0001001010000100000100",
			955 => "1111111001000000011101",
			956 => "0000110111010100000100",
			957 => "0000000001000000011101",
			958 => "0000000001000000011101",
			959 => "0000001001000000011101",
			960 => "1111111001000000011101",
			961 => "0001101010011000001100",
			962 => "0011010010011100001000",
			963 => "0001110110100100000100",
			964 => "0000000001000000011101",
			965 => "0000001001000000011101",
			966 => "0000010001000000011101",
			967 => "0010010100101100000100",
			968 => "1111111001000000011101",
			969 => "0000000001000000011101",
			970 => "0010101001101001101100",
			971 => "0001101000010000111100",
			972 => "0001000011000000011100",
			973 => "0010010100101100001100",
			974 => "0000101000001100001000",
			975 => "0011111111010100000100",
			976 => "0000001001000000011101",
			977 => "1111111001000000011101",
			978 => "0000010001000000011101",
			979 => "0001011100100100001000",
			980 => "0011100010000100000100",
			981 => "1111111001000000011101",
			982 => "0000001001000000011101",
			983 => "0011011001011100000100",
			984 => "1111111001000000011101",
			985 => "0000001001000000011101",
			986 => "0011001000111100010000",
			987 => "0011011110110000001000",
			988 => "0001001100111100000100",
			989 => "1111111001000000011101",
			990 => "0000001001000000011101",
			991 => "0001101001100100000100",
			992 => "0000000001000000011101",
			993 => "0000001001000000011101",
			994 => "0000111011011100001000",
			995 => "0001000011010100000100",
			996 => "1111111001000000011101",
			997 => "0000000001000000011101",
			998 => "0001011001110100000100",
			999 => "0000001001000000011101",
			1000 => "0000000001000000011101",
			1001 => "0001111111011100010100",
			1002 => "0001000111011100001100",
			1003 => "0010011010011000000100",
			1004 => "0000000001000000011101",
			1005 => "0010000001110000000100",
			1006 => "0000000001000000011101",
			1007 => "0000001001000000011101",
			1008 => "0000011101011100000100",
			1009 => "0000001001000000011101",
			1010 => "1111111001000000011101",
			1011 => "0011100010110000010000",
			1012 => "0011010111010100001000",
			1013 => "0001010111111100000100",
			1014 => "0000000001000000011101",
			1015 => "1111111001000000011101",
			1016 => "0011000001011000000100",
			1017 => "0000001001000000011101",
			1018 => "0000000001000000011101",
			1019 => "0001110110110100000100",
			1020 => "0000001001000000011101",
			1021 => "0001000001101100000100",
			1022 => "0000000001000000011101",
			1023 => "0000001001000000011101",
			1024 => "0011000100000000000100",
			1025 => "0000000001000000011101",
			1026 => "0010011011101000001000",
			1027 => "0000011100100000000100",
			1028 => "1111111001000000011101",
			1029 => "0000000001000000011101",
			1030 => "1111111001000000011101",
			1031 => "0010110011011100010000",
			1032 => "0000100111011000000100",
			1033 => "1111111001000100101001",
			1034 => "0000100000010000001000",
			1035 => "0011010001111100000100",
			1036 => "0000000001000100101001",
			1037 => "0000000001000100101001",
			1038 => "0000000001000100101001",
			1039 => "0010111100101100111000",
			1040 => "0011010110100100110000",
			1041 => "0001000010111000010100",
			1042 => "0010000111000100010000",
			1043 => "0000110000011100001000",
			1044 => "0001110100000000000100",
			1045 => "0000000001000100101001",
			1046 => "1111111001000100101001",
			1047 => "0000101110110100000100",
			1048 => "0000001001000100101001",
			1049 => "0000000001000100101001",
			1050 => "1111111001000100101001",
			1051 => "0011000100000000001100",
			1052 => "0000101010000100001000",
			1053 => "0001010111001000000100",
			1054 => "0000000001000100101001",
			1055 => "0000001001000100101001",
			1056 => "0000000001000100101001",
			1057 => "0000111010011100001000",
			1058 => "0001000010010000000100",
			1059 => "1111111001000100101001",
			1060 => "0000000001000100101001",
			1061 => "0000101111010100000100",
			1062 => "0000001001000100101001",
			1063 => "0000000001000100101001",
			1064 => "0010100001010000000100",
			1065 => "0000000001000100101001",
			1066 => "0000001001000100101001",
			1067 => "0011000100000000001100",
			1068 => "0001000110001100001000",
			1069 => "0001101001100100000100",
			1070 => "0000000001000100101001",
			1071 => "0000000001000100101001",
			1072 => "1111111001000100101001",
			1073 => "0001001110100100010100",
			1074 => "0010001011010100010000",
			1075 => "0011001110001100001000",
			1076 => "0001000010010100000100",
			1077 => "0000000001000100101001",
			1078 => "1111111001000100101001",
			1079 => "0010101000100100000100",
			1080 => "0000000001000100101001",
			1081 => "0000000001000100101001",
			1082 => "0000001001000100101001",
			1083 => "0000110110111000010000",
			1084 => "0010101010110000001000",
			1085 => "0000001111000100000100",
			1086 => "0000000001000100101001",
			1087 => "1111111001000100101001",
			1088 => "0001000000010100000100",
			1089 => "0000001001000100101001",
			1090 => "0000000001000100101001",
			1091 => "0010000001110100001000",
			1092 => "0010000001010100000100",
			1093 => "0000000001000100101001",
			1094 => "0000000001000100101001",
			1095 => "0001000001101100000100",
			1096 => "1111111001000100101001",
			1097 => "0000000001000100101001",
			1098 => "0010010001111001000000",
			1099 => "0001111101100000101000",
			1100 => "0011001001110000100000",
			1101 => "0011111001100000011100",
			1102 => "0000010110101000010000",
			1103 => "0001000010111000001000",
			1104 => "0011110101110000000100",
			1105 => "0000000001001001010101",
			1106 => "1111111001001001010101",
			1107 => "0011011011000000000100",
			1108 => "0000000001001001010101",
			1109 => "0000001001001001010101",
			1110 => "0001101011001100000100",
			1111 => "0000000001001001010101",
			1112 => "0001111001110000000100",
			1113 => "0000000001001001010101",
			1114 => "0000001001001001010101",
			1115 => "1111111001001001010101",
			1116 => "0010100101000100000100",
			1117 => "1111111001001001010101",
			1118 => "0000000001001001010101",
			1119 => "0001111110001100001000",
			1120 => "0000101100111000000100",
			1121 => "1111111001001001010101",
			1122 => "0000000001001001010101",
			1123 => "0010100001110000001100",
			1124 => "0001010111010000000100",
			1125 => "0000000001001001010101",
			1126 => "0000101110010000000100",
			1127 => "0000000001001001010101",
			1128 => "0000000001001001010101",
			1129 => "0000000001001001010101",
			1130 => "0001011010011100000100",
			1131 => "0000001001001001010101",
			1132 => "0000110010000000011000",
			1133 => "0001001010110100001000",
			1134 => "0000101100010000000100",
			1135 => "0000000001001001010101",
			1136 => "1111111001001001010101",
			1137 => "0001001100111100001100",
			1138 => "0001111101111000001000",
			1139 => "0000101111100100000100",
			1140 => "0000000001001001010101",
			1141 => "0000001001001001010101",
			1142 => "0000000001001001010101",
			1143 => "0000000001001001010101",
			1144 => "0000111010000100011100",
			1145 => "0011111111010100010000",
			1146 => "0010001000100100001000",
			1147 => "0000010101011100000100",
			1148 => "0000000001001001010101",
			1149 => "0000001001001001010101",
			1150 => "0000011011111100000100",
			1151 => "0000000001001001010101",
			1152 => "0000000001001001010101",
			1153 => "0000100010010100001000",
			1154 => "0010010000001000000100",
			1155 => "0000001001001001010101",
			1156 => "0000000001001001010101",
			1157 => "0000000001001001010101",
			1158 => "0001011101000100010000",
			1159 => "0011000100011000001000",
			1160 => "0000011011111100000100",
			1161 => "0000000001001001010101",
			1162 => "0000001001001001010101",
			1163 => "0001100100111100000100",
			1164 => "0000000001001001010101",
			1165 => "0000000001001001010101",
			1166 => "0011000100011000001000",
			1167 => "0000010100110100000100",
			1168 => "1111111001001001010101",
			1169 => "0000000001001001010101",
			1170 => "0011001011000000000100",
			1171 => "0000000001001001010101",
			1172 => "0000000001001001010101",
			1173 => "0011111011110001111000",
			1174 => "0011110010010101100100",
			1175 => "0011110101110000111000",
			1176 => "0000111010011100011100",
			1177 => "0001000000101100010000",
			1178 => "0001111000111000001000",
			1179 => "0001011101010100000100",
			1180 => "0000000001001111000001",
			1181 => "0000000001001111000001",
			1182 => "0010110001111100000100",
			1183 => "1111111001001111000001",
			1184 => "0000000001001111000001",
			1185 => "0001010100011000001000",
			1186 => "0011010111001000000100",
			1187 => "0000000001001111000001",
			1188 => "0000001001001111000001",
			1189 => "0000000001001111000001",
			1190 => "0001111001110000001100",
			1191 => "0011010011100000000100",
			1192 => "0000000001001111000001",
			1193 => "0001101101011000000100",
			1194 => "0000000001001111000001",
			1195 => "0000001001001111000001",
			1196 => "0010000001110100001000",
			1197 => "0000010111100100000100",
			1198 => "1111111001001111000001",
			1199 => "0000000001001111000001",
			1200 => "0011001001110000000100",
			1201 => "0000000001001111000001",
			1202 => "0000000001001111000001",
			1203 => "0000110101110100010100",
			1204 => "0001101111000000001100",
			1205 => "0010111100101100001000",
			1206 => "0001000011110000000100",
			1207 => "0000000001001111000001",
			1208 => "0000000001001111000001",
			1209 => "1111111001001111000001",
			1210 => "0001001110111000000100",
			1211 => "0000000001001111000001",
			1212 => "0000000001001111000001",
			1213 => "0010111100101100001000",
			1214 => "0010001001101000000100",
			1215 => "0000000001001111000001",
			1216 => "0000001001001111000001",
			1217 => "0000010111100100001000",
			1218 => "0000111001010100000100",
			1219 => "0000000001001111000001",
			1220 => "0000001001001111000001",
			1221 => "0000110010000000000100",
			1222 => "0000000001001111000001",
			1223 => "0000000001001111000001",
			1224 => "0000010001111000000100",
			1225 => "1111111001001111000001",
			1226 => "0010110010001000000100",
			1227 => "0000000001001111000001",
			1228 => "0010110001001000000100",
			1229 => "0000000001001111000001",
			1230 => "0001001000011100000100",
			1231 => "0000000001001111000001",
			1232 => "0000000001001111000001",
			1233 => "0010100110011100101100",
			1234 => "0010110100010000001000",
			1235 => "0011111110000000000100",
			1236 => "0000000001001111000001",
			1237 => "0000001001001111000001",
			1238 => "0001000010100100011100",
			1239 => "0010110110100000010000",
			1240 => "0001001110100100001000",
			1241 => "0000011100011000000100",
			1242 => "0000000001001111000001",
			1243 => "0000000001001111000001",
			1244 => "0000011110010100000100",
			1245 => "0000000001001111000001",
			1246 => "0000000001001111000001",
			1247 => "0010001001101000001000",
			1248 => "0011011111010100000100",
			1249 => "0000000001001111000001",
			1250 => "0000000001001111000001",
			1251 => "0000000001001111000001",
			1252 => "0000000000111000000100",
			1253 => "0000001001001111000001",
			1254 => "0000000001001111000001",
			1255 => "0011111011001000001100",
			1256 => "0000101101001000000100",
			1257 => "0000000001001111000001",
			1258 => "0001100100101100000100",
			1259 => "0000000001001111000001",
			1260 => "1111111001001111000001",
			1261 => "0010101001101000000100",
			1262 => "0000001001001111000001",
			1263 => "0000000001001111000001",
			1264 => "0001101011001101100000",
			1265 => "0011110110111100111100",
			1266 => "0001101101011000100100",
			1267 => "0000010101011100010000",
			1268 => "0000010110101000000100",
			1269 => "1111111001010101100101",
			1270 => "0010011001011000000100",
			1271 => "0000001001010101100101",
			1272 => "0010001000010100000100",
			1273 => "1111111001010101100101",
			1274 => "0000000001010101100101",
			1275 => "0010001000100100000100",
			1276 => "0000011001010101100101",
			1277 => "0011100110010000001000",
			1278 => "0010010101010000000100",
			1279 => "0000001001010101100101",
			1280 => "1111111001010101100101",
			1281 => "0011011111010000000100",
			1282 => "0000011001010101100101",
			1283 => "1111111001010101100101",
			1284 => "0000101110110100010100",
			1285 => "0000111001110100000100",
			1286 => "1111111001010101100101",
			1287 => "0001000010110000001000",
			1288 => "0000110001011000000100",
			1289 => "1111111001010101100101",
			1290 => "0000010001010101100101",
			1291 => "0011001000111000000100",
			1292 => "0000110001010101100101",
			1293 => "0000000001010101100101",
			1294 => "1111111001010101100101",
			1295 => "0011000100011000010000",
			1296 => "0000101111010100000100",
			1297 => "0000101001010101100101",
			1298 => "0011110000010000001000",
			1299 => "0001110001101000000100",
			1300 => "1111111001010101100101",
			1301 => "0000000001010101100101",
			1302 => "0000011001010101100101",
			1303 => "0001001101101100001100",
			1304 => "0010111011011100001000",
			1305 => "0010000001010000000100",
			1306 => "0000010001010101100101",
			1307 => "1111111001010101100101",
			1308 => "1111111001010101100101",
			1309 => "0001000011000000000100",
			1310 => "0000101001010101100101",
			1311 => "0000000001010101100101",
			1312 => "0011000110100101001000",
			1313 => "0010101000010100100000",
			1314 => "0001101111000000010000",
			1315 => "0010011001111100000100",
			1316 => "0000011001010101100101",
			1317 => "0010100011101000000100",
			1318 => "0000010001010101100101",
			1319 => "0001110110100100000100",
			1320 => "1111111001010101100101",
			1321 => "0000000001010101100101",
			1322 => "0001111001001000000100",
			1323 => "0000100001010101100101",
			1324 => "0001100100111100000100",
			1325 => "0000011001010101100101",
			1326 => "0000010100110100000100",
			1327 => "0000000001010101100101",
			1328 => "0000010001010101100101",
			1329 => "0001000011111000100000",
			1330 => "0001101001100100010000",
			1331 => "0001110101101100001000",
			1332 => "0010110011011100000100",
			1333 => "1111111001010101100101",
			1334 => "0000011001010101100101",
			1335 => "0010001100000100000100",
			1336 => "0000001001010101100101",
			1337 => "1111111001010101100101",
			1338 => "0001110111010000001000",
			1339 => "0001111101100000000100",
			1340 => "0000011001010101100101",
			1341 => "0000011001010101100101",
			1342 => "0000101100001100000100",
			1343 => "1111111001010101100101",
			1344 => "0000010001010101100101",
			1345 => "0011001000111100000100",
			1346 => "0000010001010101100101",
			1347 => "1111111001010101100101",
			1348 => "0011001000011000011000",
			1349 => "0001100101010000010000",
			1350 => "0000011100011000001100",
			1351 => "0001110101100100001000",
			1352 => "0010011010100000000100",
			1353 => "1111111001010101100101",
			1354 => "0000000001010101100101",
			1355 => "0000011001010101100101",
			1356 => "1111111001010101100101",
			1357 => "0000011100011000000100",
			1358 => "0000000001010101100101",
			1359 => "0000110001010101100101",
			1360 => "0000011000010000010000",
			1361 => "0010011000010100001100",
			1362 => "0001101111000000000100",
			1363 => "0000000001010101100101",
			1364 => "0001110000011100000100",
			1365 => "0000000001010101100101",
			1366 => "1111111001010101100101",
			1367 => "0000000001010101100101",
			1368 => "0000010001010101100101",
			1369 => "0001101001100101010100",
			1370 => "0001010111001000000100",
			1371 => "1111111001011010100001",
			1372 => "0011111110000100100100",
			1373 => "0010101010110000010100",
			1374 => "0000100001000000001100",
			1375 => "0011000110000100000100",
			1376 => "0000000001011010100001",
			1377 => "0001011011011100000100",
			1378 => "0000000001011010100001",
			1379 => "0000000001011010100001",
			1380 => "0011110001000000000100",
			1381 => "1111111001011010100001",
			1382 => "0000000001011010100001",
			1383 => "0001101101011000000100",
			1384 => "0000000001011010100001",
			1385 => "0011001000111000001000",
			1386 => "0011100100001000000100",
			1387 => "0000000001011010100001",
			1388 => "0000001001011010100001",
			1389 => "0000000001011010100001",
			1390 => "0001001000000100011000",
			1391 => "0010011110010100001000",
			1392 => "0001001011110000000100",
			1393 => "0000000001011010100001",
			1394 => "0000001001011010100001",
			1395 => "0010010111101100001000",
			1396 => "0001110111010000000100",
			1397 => "0000000001011010100001",
			1398 => "0000000001011010100001",
			1399 => "0010001010110000000100",
			1400 => "0000000001011010100001",
			1401 => "0000000001011010100001",
			1402 => "0000101100010000001100",
			1403 => "0000100110010000000100",
			1404 => "0000000001011010100001",
			1405 => "0011001000111000000100",
			1406 => "0000000001011010100001",
			1407 => "0000000001011010100001",
			1408 => "0011000111001000000100",
			1409 => "1111111001011010100001",
			1410 => "0000000001011010100001",
			1411 => "0001111101100000011000",
			1412 => "0010111100101100010100",
			1413 => "0011111110010000010000",
			1414 => "0010011001011000001100",
			1415 => "0001000100001100000100",
			1416 => "1111111001011010100001",
			1417 => "0000101010000100000100",
			1418 => "0000001001011010100001",
			1419 => "0000000001011010100001",
			1420 => "0000001001011010100001",
			1421 => "0000000001011010100001",
			1422 => "0000001001011010100001",
			1423 => "0011000100000000001000",
			1424 => "0010001011010100000100",
			1425 => "0000000001011010100001",
			1426 => "1111111001011010100001",
			1427 => "0000000111111000011100",
			1428 => "0010101100011100010000",
			1429 => "0010000111000100001000",
			1430 => "0011001001110000000100",
			1431 => "0000001001011010100001",
			1432 => "0000000001011010100001",
			1433 => "0011110110010000000100",
			1434 => "0000000001011010100001",
			1435 => "1111111001011010100001",
			1436 => "0011001000000000000100",
			1437 => "0000001001011010100001",
			1438 => "0011110000010100000100",
			1439 => "1111111001011010100001",
			1440 => "0000000001011010100001",
			1441 => "0001111101100000000100",
			1442 => "0000000001011010100001",
			1443 => "0011101011001000000100",
			1444 => "1111111001011010100001",
			1445 => "0011000101110100000100",
			1446 => "0000000001011010100001",
			1447 => "0000000001011010100001",
			1448 => "0011101110101101010100",
			1449 => "0010111100101100101100",
			1450 => "0001001000000100001100",
			1451 => "0011000100000000000100",
			1452 => "0000000001100000010101",
			1453 => "0011011001110100000100",
			1454 => "1111111001100000010101",
			1455 => "0000000001100000010101",
			1456 => "0000110000011100010000",
			1457 => "0010101010110000000100",
			1458 => "1111111001100000010101",
			1459 => "0011111001010000001000",
			1460 => "0000111001110100000100",
			1461 => "0000000001100000010101",
			1462 => "0000000001100000010101",
			1463 => "0000000001100000010101",
			1464 => "0011111110010000001000",
			1465 => "0011011011000000000100",
			1466 => "0000000001100000010101",
			1467 => "0000001001100000010101",
			1468 => "0011010110100100000100",
			1469 => "1111111001100000010101",
			1470 => "0000000001100000010101",
			1471 => "0000010111100100010100",
			1472 => "0011011001001000000100",
			1473 => "0000000001100000010101",
			1474 => "0001101000010000001100",
			1475 => "0001101001011000000100",
			1476 => "0000000001100000010101",
			1477 => "0010100110011100000100",
			1478 => "1111111001100000010101",
			1479 => "0000000001100000010101",
			1480 => "0000000001100000010101",
			1481 => "0010110000001100000100",
			1482 => "0000000001100000010101",
			1483 => "0001101101011000001100",
			1484 => "0011001110001100000100",
			1485 => "0000000001100000010101",
			1486 => "0011010001011000000100",
			1487 => "0000000001100000010101",
			1488 => "0000000001100000010101",
			1489 => "0000000001100000010101",
			1490 => "0011111111100100110100",
			1491 => "0001100100111100110000",
			1492 => "0011110110111100011000",
			1493 => "0000101100010000010000",
			1494 => "0011100101001000001000",
			1495 => "0001110011100000000100",
			1496 => "0000000001100000010101",
			1497 => "0000000001100000010101",
			1498 => "0010110101100100000100",
			1499 => "0000000001100000010101",
			1500 => "0000000001100000010101",
			1501 => "0010110000001100000100",
			1502 => "0000000001100000010101",
			1503 => "1111111001100000010101",
			1504 => "0000111010000100001100",
			1505 => "0000011101111100001000",
			1506 => "0000111100010000000100",
			1507 => "0000000001100000010101",
			1508 => "0000000001100000010101",
			1509 => "0000000001100000010101",
			1510 => "0001110110100100000100",
			1511 => "0000000001100000010101",
			1512 => "0001001111100100000100",
			1513 => "0000000001100000010101",
			1514 => "0000000001100000010101",
			1515 => "0000001001100000010101",
			1516 => "0000111110110100000100",
			1517 => "1111111001100000010101",
			1518 => "0000010111101000010100",
			1519 => "0010000010101000001100",
			1520 => "0010001011010100001000",
			1521 => "0010100110011000000100",
			1522 => "0000000001100000010101",
			1523 => "0000000001100000010101",
			1524 => "0000001001100000010101",
			1525 => "0000010000111100000100",
			1526 => "0000000001100000010101",
			1527 => "0000000001100000010101",
			1528 => "0000010001111000001100",
			1529 => "0010101100011100001000",
			1530 => "0010111011011100000100",
			1531 => "0000000001100000010101",
			1532 => "1111111001100000010101",
			1533 => "0000000001100000010101",
			1534 => "0001000100001100001000",
			1535 => "0000000001110100000100",
			1536 => "0000000001100000010101",
			1537 => "0000000001100000010101",
			1538 => "0010100001010100000100",
			1539 => "0000000001100000010101",
			1540 => "0000000001100000010101",
			1541 => "0001101011001101011000",
			1542 => "0010011000010000110100",
			1543 => "0001101011001100100000",
			1544 => "0001101001011000001000",
			1545 => "0000001100000100000100",
			1546 => "1111111001100110110001",
			1547 => "0000010001100110110001",
			1548 => "0001101101011000001100",
			1549 => "0011101011011100000100",
			1550 => "1111111001100110110001",
			1551 => "0011010100010000000100",
			1552 => "0000001001100110110001",
			1553 => "1111111001100110110001",
			1554 => "0011101011000000000100",
			1555 => "1111111001100110110001",
			1556 => "0011100110100100000100",
			1557 => "0000001001100110110001",
			1558 => "1111111001100110110001",
			1559 => "0000100010000100010000",
			1560 => "0011101010111000000100",
			1561 => "1111111001100110110001",
			1562 => "0010101010110000001000",
			1563 => "0000000010011000000100",
			1564 => "0000000001100110110001",
			1565 => "1111111001100110110001",
			1566 => "0000001001100110110001",
			1567 => "1111111001100110110001",
			1568 => "0011101110110100001100",
			1569 => "0001111110110000001000",
			1570 => "0001001100111000000100",
			1571 => "0000010001100110110001",
			1572 => "1111111001100110110001",
			1573 => "1111111001100110110001",
			1574 => "0011000100011000001000",
			1575 => "0001010110100000000100",
			1576 => "0000000001100110110001",
			1577 => "1111111001100110110001",
			1578 => "0001001101101100001100",
			1579 => "0001010111100000001000",
			1580 => "0010100010101100000100",
			1581 => "0000010001100110110001",
			1582 => "0000000001100110110001",
			1583 => "1111111001100110110001",
			1584 => "0000011001100110110001",
			1585 => "0010110001001001001100",
			1586 => "0010000001010100100000",
			1587 => "0001001000110100011100",
			1588 => "0010010111101100001100",
			1589 => "0011000100011000001000",
			1590 => "0001101011001100000100",
			1591 => "1111111001100110110001",
			1592 => "0000001001100110110001",
			1593 => "0000010001100110110001",
			1594 => "0010100111110100001000",
			1595 => "0010100011101000000100",
			1596 => "0000000001100110110001",
			1597 => "1111111001100110110001",
			1598 => "0010110110110100000100",
			1599 => "0000001001100110110001",
			1600 => "1111111001100110110001",
			1601 => "1111111001100110110001",
			1602 => "0001000100001100010100",
			1603 => "0011011110110000000100",
			1604 => "1111111001100110110001",
			1605 => "0000011011101000001000",
			1606 => "0001110101101100000100",
			1607 => "0000001001100110110001",
			1608 => "1111111001100110110001",
			1609 => "0000001010101100000100",
			1610 => "0000000001100110110001",
			1611 => "0000001001100110110001",
			1612 => "0011001000111000001100",
			1613 => "0001010100001000000100",
			1614 => "1111111001100110110001",
			1615 => "0010011101101000000100",
			1616 => "0000010001100110110001",
			1617 => "0000001001100110110001",
			1618 => "0001101111000000000100",
			1619 => "1111111001100110110001",
			1620 => "0011000110000100000100",
			1621 => "0000001001100110110001",
			1622 => "0000000001100110110001",
			1623 => "0010011000100100100100",
			1624 => "0001110001011000001100",
			1625 => "0011011100010000000100",
			1626 => "1111111001100110110001",
			1627 => "0011101000000100000100",
			1628 => "0000011001100110110001",
			1629 => "0000000001100110110001",
			1630 => "0000010001111000001100",
			1631 => "0010101010110000001000",
			1632 => "0011010110111100000100",
			1633 => "0000000001100110110001",
			1634 => "0000011001100110110001",
			1635 => "1111111001100110110001",
			1636 => "0011011010000100000100",
			1637 => "1111111001100110110001",
			1638 => "0011101110100100000100",
			1639 => "0000011001100110110001",
			1640 => "1111111001100110110001",
			1641 => "0011100000010100000100",
			1642 => "1111111001100110110001",
			1643 => "0000001001100110110001",
			1644 => "0001101011001100111100",
			1645 => "0000010101011100011100",
			1646 => "0001101001011000001000",
			1647 => "0000010111100100000100",
			1648 => "1111111001101100100101",
			1649 => "0000001001101100100101",
			1650 => "0011101011000000000100",
			1651 => "1111111001101100100101",
			1652 => "0011010100010000001100",
			1653 => "0001111101010100001000",
			1654 => "0000001110111100000100",
			1655 => "1111111001101100100101",
			1656 => "0000001001101100100101",
			1657 => "0000011001101100100101",
			1658 => "1111111001101100100101",
			1659 => "0011111111010100010000",
			1660 => "0011100111111100000100",
			1661 => "0000001001101100100101",
			1662 => "0011101110110100000100",
			1663 => "1111111001101100100101",
			1664 => "0001011101000100000100",
			1665 => "0000001001101100100101",
			1666 => "1111111001101100100101",
			1667 => "0001010101110000001100",
			1668 => "0001010111100000001000",
			1669 => "0001011100100100000100",
			1670 => "0000000001101100100101",
			1671 => "0000011001101100100101",
			1672 => "1111111001101100100101",
			1673 => "0000011001101100100101",
			1674 => "0011001000011001011100",
			1675 => "0001101000010000111000",
			1676 => "0001111101100000011100",
			1677 => "0011011110110000001100",
			1678 => "0001000000101100001000",
			1679 => "0011110000110100000100",
			1680 => "0000000001101100100101",
			1681 => "1111111001101100100101",
			1682 => "0000001001101100100101",
			1683 => "0011111001011100001000",
			1684 => "0011011011000000000100",
			1685 => "0000001001101100100101",
			1686 => "0000001001101100100101",
			1687 => "0010011001011000000100",
			1688 => "1111111001101100100101",
			1689 => "0000001001101100100101",
			1690 => "0001010010110100010000",
			1691 => "0001001111101000001000",
			1692 => "0000011110010100000100",
			1693 => "0000010001101100100101",
			1694 => "1111111001101100100101",
			1695 => "0001110101101100000100",
			1696 => "0000000001101100100101",
			1697 => "1111111001101100100101",
			1698 => "0000011100011000001000",
			1699 => "0000000110001000000100",
			1700 => "0000000001101100100101",
			1701 => "0000001001101100100101",
			1702 => "1111111001101100100101",
			1703 => "0000001010101100001000",
			1704 => "0011111111101000000100",
			1705 => "0000000001101100100101",
			1706 => "1111111001101100100101",
			1707 => "0010111011110100010000",
			1708 => "0001000100001100001000",
			1709 => "0000011011101000000100",
			1710 => "0000001001101100100101",
			1711 => "0000001001101100100101",
			1712 => "0011001110001100000100",
			1713 => "0000001001101100100101",
			1714 => "1111111001101100100101",
			1715 => "0001101000010000000100",
			1716 => "0000011001101100100101",
			1717 => "0011111000001000000100",
			1718 => "1111111001101100100101",
			1719 => "0000001001101100100101",
			1720 => "0000011000010000100000",
			1721 => "0010100110011100011100",
			1722 => "0000010111101000010000",
			1723 => "0011010110111100001000",
			1724 => "0001000100001100000100",
			1725 => "1111111001101100100101",
			1726 => "0000001001101100100101",
			1727 => "0010100001010000000100",
			1728 => "0000110001101100100101",
			1729 => "0000001001101100100101",
			1730 => "0001000011101100001000",
			1731 => "0011011010000100000100",
			1732 => "1111111001101100100101",
			1733 => "0000000001101100100101",
			1734 => "0000001001101100100101",
			1735 => "1111111001101100100101",
			1736 => "0000001001101100100101",
			1737 => "0010110011011100001100",
			1738 => "0000101111010100000100",
			1739 => "1111111001110000011001",
			1740 => "0000001100110000000100",
			1741 => "0000000001110000011001",
			1742 => "0000001001110000011001",
			1743 => "0010001111000101101000",
			1744 => "0001100100111100110100",
			1745 => "0010001010110000011000",
			1746 => "0001001111100100001100",
			1747 => "0010110101100100001000",
			1748 => "0011100111011000000100",
			1749 => "0000000001110000011001",
			1750 => "1111111001110000011001",
			1751 => "1111111001110000011001",
			1752 => "0011001001110100001000",
			1753 => "0011000100011000000100",
			1754 => "0000000001110000011001",
			1755 => "0000001001110000011001",
			1756 => "0000000001110000011001",
			1757 => "0011001000111100001100",
			1758 => "0001101101011000000100",
			1759 => "1111111001110000011001",
			1760 => "0011110010000000000100",
			1761 => "0000000001110000011001",
			1762 => "1111111001110000011001",
			1763 => "0001001000000100001000",
			1764 => "0010001001101000000100",
			1765 => "0000000001110000011001",
			1766 => "1111111001110000011001",
			1767 => "0010011001111100000100",
			1768 => "0000000001110000011001",
			1769 => "1111111001110000011001",
			1770 => "0011001100110000011000",
			1771 => "0011000100000000001000",
			1772 => "0001011001110100000100",
			1773 => "1111111001110000011001",
			1774 => "0000000001110000011001",
			1775 => "0010011010011000001000",
			1776 => "0000101111010100000100",
			1777 => "0000000001110000011001",
			1778 => "0000001001110000011001",
			1779 => "0011000011011100000100",
			1780 => "0000000001110000011001",
			1781 => "0000001001110000011001",
			1782 => "0010011100011000001100",
			1783 => "0000011011101000000100",
			1784 => "1111111001110000011001",
			1785 => "0000011111001100000100",
			1786 => "0000001001110000011001",
			1787 => "0000000001110000011001",
			1788 => "0011010111111100001000",
			1789 => "0000011110010100000100",
			1790 => "0000000001110000011001",
			1791 => "0000001001110000011001",
			1792 => "0011111000110100000100",
			1793 => "0000000001110000011001",
			1794 => "0000000001110000011001",
			1795 => "0011001000111100000100",
			1796 => "0000001001110000011001",
			1797 => "1111111001110000011001",
			1798 => "0001101101011001001100",
			1799 => "0010011000010000100100",
			1800 => "0000010110101000001100",
			1801 => "0000111010001100000100",
			1802 => "1111111001110110101101",
			1803 => "0000110100000100000100",
			1804 => "0000001001110110101101",
			1805 => "1111111001110110101101",
			1806 => "0010011001011000000100",
			1807 => "0000001001110110101101",
			1808 => "0011010010110100010000",
			1809 => "0000011101011100001000",
			1810 => "0011100010001000000100",
			1811 => "1111111001110110101101",
			1812 => "0000000001110110101101",
			1813 => "0010110011100000000100",
			1814 => "0000000001110110101101",
			1815 => "0000011001110110101101",
			1816 => "1111111001110110101101",
			1817 => "0001111001001000001000",
			1818 => "0011011110101100000100",
			1819 => "0000001001110110101101",
			1820 => "1111111001110110101101",
			1821 => "0001110110100100010000",
			1822 => "0011100010000000000100",
			1823 => "1111111001110110101101",
			1824 => "0000010001000100000100",
			1825 => "0000000001110110101101",
			1826 => "0010001001000100000100",
			1827 => "0000011001110110101101",
			1828 => "0000001001110110101101",
			1829 => "0000001001101000001000",
			1830 => "0010110101100100000100",
			1831 => "0000001001110110101101",
			1832 => "1111111001110110101101",
			1833 => "0011001001110100000100",
			1834 => "0000010001110110101101",
			1835 => "1111111001110110101101",
			1836 => "0011001000011001011000",
			1837 => "0001101000010000110100",
			1838 => "0011001000111100010100",
			1839 => "0010110011011100001000",
			1840 => "0001000110110000000100",
			1841 => "1111111001110110101101",
			1842 => "0000000001110110101101",
			1843 => "0000010111100100001000",
			1844 => "0011111110010000000100",
			1845 => "0000001001110110101101",
			1846 => "0000000001110110101101",
			1847 => "0000001001110110101101",
			1848 => "0010001001101000010000",
			1849 => "0010000001110000001000",
			1850 => "0010110110110100000100",
			1851 => "0000000001110110101101",
			1852 => "0000000001110110101101",
			1853 => "0001101001100100000100",
			1854 => "0000000001110110101101",
			1855 => "0000001001110110101101",
			1856 => "0001110101101100001000",
			1857 => "0000111011011100000100",
			1858 => "1111111001110110101101",
			1859 => "0000001001110110101101",
			1860 => "0010100110011100000100",
			1861 => "1111111001110110101101",
			1862 => "0000000001110110101101",
			1863 => "0010111011110100010100",
			1864 => "0001000011010100001100",
			1865 => "0000111100010100000100",
			1866 => "0000001001110110101101",
			1867 => "0010101001000100000100",
			1868 => "0000001001110110101101",
			1869 => "0000001001110110101101",
			1870 => "0011000110000100000100",
			1871 => "0000001001110110101101",
			1872 => "1111111001110110101101",
			1873 => "0011101011110000000100",
			1874 => "1111111001110110101101",
			1875 => "0011001001110100000100",
			1876 => "1111111001110110101101",
			1877 => "0001100101010000000100",
			1878 => "1111111001110110101101",
			1879 => "0000001001110110101101",
			1880 => "0010011000010100100000",
			1881 => "0010101010110000011100",
			1882 => "0011011010000100010000",
			1883 => "0010011001111100001000",
			1884 => "0011011100000000000100",
			1885 => "1111111001110110101101",
			1886 => "0000010001110110101101",
			1887 => "0010110110100000000100",
			1888 => "1111111001110110101101",
			1889 => "0000000001110110101101",
			1890 => "0010000001010100000100",
			1891 => "0000100001110110101101",
			1892 => "0010011010100000000100",
			1893 => "0000010001110110101101",
			1894 => "1111111001110110101101",
			1895 => "1111111001110110101101",
			1896 => "0011110000010100000100",
			1897 => "0000000001110110101101",
			1898 => "0000001001110110101101",
			1899 => "0001001011110001001100",
			1900 => "0001101001100100111100",
			1901 => "0011000100001000001100",
			1902 => "0000100010110100000100",
			1903 => "0000000001111101011001",
			1904 => "0011000100000000000100",
			1905 => "0000000001111101011001",
			1906 => "0000000001111101011001",
			1907 => "0011000100011000011000",
			1908 => "0011101100000000001100",
			1909 => "0001011001010100001000",
			1910 => "0000011011111100000100",
			1911 => "0000000001111101011001",
			1912 => "0000000001111101011001",
			1913 => "0000000001111101011001",
			1914 => "0001010111100000001000",
			1915 => "0010110000011100000100",
			1916 => "0000000001111101011001",
			1917 => "0000000001111101011001",
			1918 => "0000000001111101011001",
			1919 => "0011101100000000001100",
			1920 => "0011111111010100000100",
			1921 => "0000000001111101011001",
			1922 => "0011110111010100000100",
			1923 => "0000000001111101011001",
			1924 => "0000000001111101011001",
			1925 => "0010100010101100000100",
			1926 => "0000000001111101011001",
			1927 => "0000011011111100000100",
			1928 => "0000000001111101011001",
			1929 => "0000000001111101011001",
			1930 => "0010100111110100000100",
			1931 => "0000000001111101011001",
			1932 => "0011101100111000001000",
			1933 => "0001111111011100000100",
			1934 => "0000000001111101011001",
			1935 => "0000000001111101011001",
			1936 => "0000000001111101011001",
			1937 => "0001001110111001000100",
			1938 => "0001100100111100011000",
			1939 => "0001111000111000001100",
			1940 => "0011011011000000001000",
			1941 => "0010110101101100000100",
			1942 => "0000000001111101011001",
			1943 => "0000000001111101011001",
			1944 => "0000000001111101011001",
			1945 => "0010110001001000001000",
			1946 => "0000100110010000000100",
			1947 => "0000000001111101011001",
			1948 => "0000000001111101011001",
			1949 => "0000000001111101011001",
			1950 => "0001101000010000010000",
			1951 => "0000111101000100000100",
			1952 => "0000000001111101011001",
			1953 => "0001001100001100000100",
			1954 => "0000000001111101011001",
			1955 => "0000011010011000000100",
			1956 => "0000000001111101011001",
			1957 => "0000000001111101011001",
			1958 => "0010110101110100010000",
			1959 => "0000010001000100001000",
			1960 => "0010101100011100000100",
			1961 => "0000000001111101011001",
			1962 => "0000000001111101011001",
			1963 => "0010000001110000000100",
			1964 => "0000000001111101011001",
			1965 => "0000001001111101011001",
			1966 => "0000011010011000001000",
			1967 => "0010001001101000000100",
			1968 => "1111111001111101011001",
			1969 => "0000000001111101011001",
			1970 => "0000000001111101011001",
			1971 => "0011100110010000101000",
			1972 => "0000011001111000011000",
			1973 => "0011000100000000001100",
			1974 => "0001011010111100000100",
			1975 => "0000000001111101011001",
			1976 => "0010110101101100000100",
			1977 => "0000001001111101011001",
			1978 => "0000000001111101011001",
			1979 => "0001000010010000001000",
			1980 => "0001110100000000000100",
			1981 => "0000000001111101011001",
			1982 => "1111111001111101011001",
			1983 => "0000000001111101011001",
			1984 => "0010001111000100001100",
			1985 => "0001101001100100000100",
			1986 => "0000000001111101011001",
			1987 => "0001000011111000000100",
			1988 => "0000001001111101011001",
			1989 => "0000000001111101011001",
			1990 => "0000000001111101011001",
			1991 => "0011100010110000001100",
			1992 => "0011010111010100001000",
			1993 => "0011001000000000000100",
			1994 => "0000000001111101011001",
			1995 => "1111111001111101011001",
			1996 => "0000000001111101011001",
			1997 => "0011011101101100001100",
			1998 => "0000011101111100000100",
			1999 => "0000000001111101011001",
			2000 => "0000010100111100000100",
			2001 => "0000000001111101011001",
			2002 => "0000000001111101011001",
			2003 => "0011000101110100000100",
			2004 => "0000000001111101011001",
			2005 => "0000000001111101011001",
			2006 => "0001101101011000101000",
			2007 => "0000010001000100010100",
			2008 => "0010001001000100010000",
			2009 => "0000000001110000000100",
			2010 => "1111111010000011000101",
			2011 => "0000011101011100001000",
			2012 => "0010010010001100000100",
			2013 => "0000000010000011000101",
			2014 => "0000001010000011000101",
			2015 => "1111111010000011000101",
			2016 => "1111111010000011000101",
			2017 => "0000111010000100010000",
			2018 => "0011010010011100001100",
			2019 => "0010010100101100001000",
			2020 => "0010110101100100000100",
			2021 => "1111111010000011000101",
			2022 => "0000000010000011000101",
			2023 => "0000001010000011000101",
			2024 => "0000010010000011000101",
			2025 => "1111111010000011000101",
			2026 => "0001010111111101100000",
			2027 => "0001101000010000110100",
			2028 => "0001001110000000011000",
			2029 => "0000010111100100001000",
			2030 => "0010111100101100000100",
			2031 => "0000000010000011000101",
			2032 => "1111111010000011000101",
			2033 => "0000000001110100001000",
			2034 => "0010100011101000000100",
			2035 => "0000001010000011000101",
			2036 => "0000000010000011000101",
			2037 => "0001101001100100000100",
			2038 => "0000000010000011000101",
			2039 => "0000001010000011000101",
			2040 => "0010111100101100001100",
			2041 => "0010110011011100000100",
			2042 => "1111111010000011000101",
			2043 => "0001111000111000000100",
			2044 => "0000001010000011000101",
			2045 => "0000000010000011000101",
			2046 => "0010001111001000001000",
			2047 => "0010101010110000000100",
			2048 => "0000000010000011000101",
			2049 => "0000001010000011000101",
			2050 => "0010011100011000000100",
			2051 => "1111111010000011000101",
			2052 => "0000000010000011000101",
			2053 => "0001000100001100011000",
			2054 => "0000001010101100001000",
			2055 => "0010110010001000000100",
			2056 => "1111111010000011000101",
			2057 => "0000001010000011000101",
			2058 => "0001111111011100001000",
			2059 => "0000011011101000000100",
			2060 => "0000000010000011000101",
			2061 => "0000001010000011000101",
			2062 => "0011111000110100000100",
			2063 => "1111111010000011000101",
			2064 => "0000001010000011000101",
			2065 => "0000010111100100001000",
			2066 => "0001101000010000000100",
			2067 => "0000001010000011000101",
			2068 => "0000001010000011000101",
			2069 => "0001001100111100001000",
			2070 => "0011001000000000000100",
			2071 => "0000000010000011000101",
			2072 => "1111111010000011000101",
			2073 => "1111111010000011000101",
			2074 => "0000001011000100101100",
			2075 => "0011011111010100011100",
			2076 => "0010010100101100001100",
			2077 => "0011001111011100001000",
			2078 => "0011011100000000000100",
			2079 => "0000000010000011000101",
			2080 => "0000001010000011000101",
			2081 => "0000000010000011000101",
			2082 => "0011010110111100001000",
			2083 => "0011111010110100000100",
			2084 => "1111111010000011000101",
			2085 => "0000001010000011000101",
			2086 => "0010101000010100000100",
			2087 => "0000010010000011000101",
			2088 => "1111111010000011000101",
			2089 => "0000000111000000000100",
			2090 => "0000010010000011000101",
			2091 => "0010010111101100000100",
			2092 => "0000001010000011000101",
			2093 => "0001101001111100000100",
			2094 => "1111111010000011000101",
			2095 => "0000000010000011000101",
			2096 => "1111111010000011000101",
			2097 => "0010010111101110000100",
			2098 => "0010001011010101000100",
			2099 => "0010101000010100100100",
			2100 => "0011000100011000010000",
			2101 => "0011011111010000001100",
			2102 => "0011000110000100000100",
			2103 => "0000000010001001011001",
			2104 => "0000011011101000000100",
			2105 => "0000000010001001011001",
			2106 => "0000000010001001011001",
			2107 => "1111111010001001011001",
			2108 => "0000001111001000001100",
			2109 => "0001110001101000000100",
			2110 => "0000000010001001011001",
			2111 => "0011001001110100000100",
			2112 => "0000000010001001011001",
			2113 => "0000000010001001011001",
			2114 => "0000111010000100000100",
			2115 => "0000000010001001011001",
			2116 => "0000000010001001011001",
			2117 => "0001000110111000001100",
			2118 => "0010111101111000001000",
			2119 => "0000010111100100000100",
			2120 => "0000000010001001011001",
			2121 => "0000000010001001011001",
			2122 => "0000000010001001011001",
			2123 => "0000111111101000001100",
			2124 => "0001111000111000000100",
			2125 => "0000000010001001011001",
			2126 => "0011000000101000000100",
			2127 => "0000000010001001011001",
			2128 => "1111111010001001011001",
			2129 => "0011101111101000000100",
			2130 => "0000000010001001011001",
			2131 => "0000000010001001011001",
			2132 => "0000011011101000100100",
			2133 => "0011001100110000100000",
			2134 => "0000111010011100010000",
			2135 => "0001111000111000001000",
			2136 => "0001101001100100000100",
			2137 => "0000000010001001011001",
			2138 => "0000000010001001011001",
			2139 => "0001000010010000000100",
			2140 => "1111111010001001011001",
			2141 => "0000000010001001011001",
			2142 => "0011100110100100001000",
			2143 => "0001111101100000000100",
			2144 => "0000001010001001011001",
			2145 => "0000000010001001011001",
			2146 => "0000110101110100000100",
			2147 => "0000000010001001011001",
			2148 => "0000000010001001011001",
			2149 => "1111111010001001011001",
			2150 => "0001011010010100001100",
			2151 => "0001000000100000001000",
			2152 => "0001101000010000000100",
			2153 => "0000000010001001011001",
			2154 => "0000001010001001011001",
			2155 => "0000000010001001011001",
			2156 => "0001010111100000000100",
			2157 => "1111111010001001011001",
			2158 => "0001000011110100000100",
			2159 => "0000000010001001011001",
			2160 => "0010100110011100000100",
			2161 => "0000001010001001011001",
			2162 => "0000000010001001011001",
			2163 => "0010011010100000100100",
			2164 => "0011101100010000000100",
			2165 => "0000000010001001011001",
			2166 => "0001000100001100011000",
			2167 => "0000000111000100001100",
			2168 => "0010100011101000001000",
			2169 => "0001110001101000000100",
			2170 => "0000000010001001011001",
			2171 => "0000000010001001011001",
			2172 => "0000000010001001011001",
			2173 => "0010100111110100000100",
			2174 => "0000000010001001011001",
			2175 => "0001111000011000000100",
			2176 => "0000001010001001011001",
			2177 => "0000000010001001011001",
			2178 => "0010101010110000000100",
			2179 => "0000000010001001011001",
			2180 => "0000000010001001011001",
			2181 => "0011100011010100100000",
			2182 => "0010111101000100011100",
			2183 => "0000010100110100001100",
			2184 => "0011101000110100001000",
			2185 => "0011010101110000000100",
			2186 => "0000000010001001011001",
			2187 => "0000000010001001011001",
			2188 => "0000000010001001011001",
			2189 => "0000011100011000001000",
			2190 => "0010000101000100000100",
			2191 => "0000000010001001011001",
			2192 => "0000001010001001011001",
			2193 => "0010110110100000000100",
			2194 => "0000000010001001011001",
			2195 => "0000000010001001011001",
			2196 => "1111111010001001011001",
			2197 => "0000000010001001011001",
			2198 => "0010001001000100011100",
			2199 => "0001110001101000011000",
			2200 => "0011001110001100000100",
			2201 => "0000000010001111000101",
			2202 => "0010111011011100010000",
			2203 => "0010000010101100000100",
			2204 => "0000000010001111000101",
			2205 => "0011010101110000001000",
			2206 => "0001010111100000000100",
			2207 => "0000000010001111000101",
			2208 => "0000000010001111000101",
			2209 => "0000000010001111000101",
			2210 => "0000000010001111000101",
			2211 => "0000000010001111000101",
			2212 => "0000000011010001010000",
			2213 => "0000010111100100100100",
			2214 => "0001111101100000011000",
			2215 => "0001010100011000010000",
			2216 => "0010110101101100001000",
			2217 => "0001000010110000000100",
			2218 => "0000000010001111000101",
			2219 => "0000000010001111000101",
			2220 => "0001111001110000000100",
			2221 => "0000000010001111000101",
			2222 => "0000000010001111000101",
			2223 => "0011001100001000000100",
			2224 => "0000000010001111000101",
			2225 => "1111111010001111000101",
			2226 => "0011000100000000000100",
			2227 => "0000000010001111000101",
			2228 => "0011110010011100000100",
			2229 => "0000000010001111000101",
			2230 => "0000000010001111000101",
			2231 => "0011010101100100010000",
			2232 => "0011110010000100001100",
			2233 => "0000010111100100000100",
			2234 => "0000000010001111000101",
			2235 => "0000001000101100000100",
			2236 => "0000000010001111000101",
			2237 => "0000001010001111000101",
			2238 => "0000000010001111000101",
			2239 => "0000011001011000001100",
			2240 => "0000011011101000000100",
			2241 => "0000000010001111000101",
			2242 => "0010111010111000000100",
			2243 => "0000000010001111000101",
			2244 => "1111111010001111000101",
			2245 => "0010010101010000001000",
			2246 => "0000001101010000000100",
			2247 => "0000000010001111000101",
			2248 => "0000000010001111000101",
			2249 => "0010101001000100000100",
			2250 => "0000000010001111000101",
			2251 => "0000000010001111000101",
			2252 => "0011001100110000101000",
			2253 => "0000110101110100011100",
			2254 => "0000101110110100001100",
			2255 => "0000111010011100001000",
			2256 => "0001001110111000000100",
			2257 => "0000000010001111000101",
			2258 => "0000000010001111000101",
			2259 => "0000001010001111000101",
			2260 => "0000000000111000001000",
			2261 => "0000000011010000000100",
			2262 => "0000000010001111000101",
			2263 => "1111111010001111000101",
			2264 => "0000110000011100000100",
			2265 => "0000000010001111000101",
			2266 => "0000000010001111000101",
			2267 => "0011111111100100001000",
			2268 => "0010001111001000000100",
			2269 => "0000000010001111000101",
			2270 => "0000001010001111000101",
			2271 => "0000000010001111000101",
			2272 => "0000000000111000001100",
			2273 => "0011001000011000001000",
			2274 => "0010000110001000000100",
			2275 => "0000000010001111000101",
			2276 => "0000000010001111000101",
			2277 => "0000000010001111000101",
			2278 => "0000110011011000010000",
			2279 => "0010000111000100001000",
			2280 => "0010000111000100000100",
			2281 => "0000000010001111000101",
			2282 => "0000000010001111000101",
			2283 => "0001001011100000000100",
			2284 => "0000000010001111000101",
			2285 => "1111111010001111000101",
			2286 => "0010001110111100000100",
			2287 => "0000000010001111000101",
			2288 => "0000000010001111000101",
			2289 => "0001011010111100001000",
			2290 => "0010000000101000000100",
			2291 => "1111111010010011011001",
			2292 => "0000000010010011011001",
			2293 => "0011000100000000011000",
			2294 => "0001000010111000001000",
			2295 => "0010010101011100000100",
			2296 => "0000000010010011011001",
			2297 => "0000000010010011011001",
			2298 => "0001011010111100000100",
			2299 => "0000000010010011011001",
			2300 => "0001101011001100001000",
			2301 => "0001101101011000000100",
			2302 => "0000000010010011011001",
			2303 => "0000000010010011011001",
			2304 => "0000001010010011011001",
			2305 => "0000110010000100111000",
			2306 => "0010000110001000100000",
			2307 => "0001000011000000010000",
			2308 => "0001101001100100001000",
			2309 => "0011000110000100000100",
			2310 => "0000000010010011011001",
			2311 => "0000000010010011011001",
			2312 => "0000101100010000000100",
			2313 => "0000000010010011011001",
			2314 => "0000000010010011011001",
			2315 => "0011110101110000001000",
			2316 => "0001111001110000000100",
			2317 => "0000000010010011011001",
			2318 => "0000000010010011011001",
			2319 => "0011000100000000000100",
			2320 => "0000000010010011011001",
			2321 => "1111111010010011011001",
			2322 => "0011000100000000001100",
			2323 => "0010001111001000000100",
			2324 => "0000000010010011011001",
			2325 => "0000110110100100000100",
			2326 => "0000000010010011011001",
			2327 => "1111111010010011011001",
			2328 => "0011001100110000001000",
			2329 => "0000111000011000000100",
			2330 => "0000000010010011011001",
			2331 => "0000000010010011011001",
			2332 => "1111111010010011011001",
			2333 => "0001010001000000010100",
			2334 => "0010000111000000010000",
			2335 => "0000101000101000001000",
			2336 => "0010011010100000000100",
			2337 => "0000000010010011011001",
			2338 => "0000000010010011011001",
			2339 => "0011111000101000000100",
			2340 => "0000000010010011011001",
			2341 => "0000001010010011011001",
			2342 => "0000000010010011011001",
			2343 => "0001011001010000010000",
			2344 => "0000010100110100001000",
			2345 => "0000110110111000000100",
			2346 => "1111111010010011011001",
			2347 => "0000000010010011011001",
			2348 => "0001010101001000000100",
			2349 => "0000000010010011011001",
			2350 => "0000000010010011011001",
			2351 => "0011000001011000001000",
			2352 => "0001000011101100000100",
			2353 => "0000000010010011011001",
			2354 => "0000000010010011011001",
			2355 => "0001011111100100000100",
			2356 => "1111111010010011011001",
			2357 => "0000000010010011011001",
			2358 => "0011011010111100001000",
			2359 => "0000100000010000000100",
			2360 => "1111111010011000000101",
			2361 => "0000000010011000000101",
			2362 => "0011110010011101001000",
			2363 => "0000110000011100110000",
			2364 => "0001001001001100010100",
			2365 => "0001110100000000001000",
			2366 => "0010110101101100000100",
			2367 => "0000000010011000000101",
			2368 => "0000000010011000000101",
			2369 => "0011111100100100001000",
			2370 => "0011010011100000000100",
			2371 => "0000000010011000000101",
			2372 => "0000000010011000000101",
			2373 => "1111111010011000000101",
			2374 => "0000101100010000001100",
			2375 => "0001101101011000000100",
			2376 => "0000000010011000000101",
			2377 => "0011001000111000000100",
			2378 => "0000001010011000000101",
			2379 => "0000000010011000000101",
			2380 => "0001101111000000001000",
			2381 => "0001111000111000000100",
			2382 => "0000000010011000000101",
			2383 => "1111111010011000000101",
			2384 => "0011001000111000000100",
			2385 => "0000001010011000000101",
			2386 => "0000000010011000000101",
			2387 => "0010101000010100010000",
			2388 => "0000101110000100001100",
			2389 => "0001110001111100000100",
			2390 => "0000000010011000000101",
			2391 => "0010111011000000000100",
			2392 => "0000000010011000000101",
			2393 => "0000000010011000000101",
			2394 => "0000000010011000000101",
			2395 => "0001000000101100000100",
			2396 => "0000001010011000000101",
			2397 => "0000000010011000000101",
			2398 => "0000111011011100001100",
			2399 => "0001101111000000000100",
			2400 => "1111111010011000000101",
			2401 => "0011111001011100000100",
			2402 => "0000001010011000000101",
			2403 => "0000000010011000000101",
			2404 => "0011000110100100100000",
			2405 => "0010110101110100010000",
			2406 => "0001101000010000001000",
			2407 => "0000101111010100000100",
			2408 => "0000000010011000000101",
			2409 => "0000000010011000000101",
			2410 => "0001001001000000000100",
			2411 => "0000001010011000000101",
			2412 => "0000000010011000000101",
			2413 => "0011011100010100001000",
			2414 => "0010011010100000000100",
			2415 => "1111110010011000000101",
			2416 => "0000000010011000000101",
			2417 => "0011011110110100000100",
			2418 => "0000000010011000000101",
			2419 => "1111111010011000000101",
			2420 => "0001101001111100001100",
			2421 => "0001001011110000000100",
			2422 => "0000000010011000000101",
			2423 => "0000011100011000000100",
			2424 => "0000001010011000000101",
			2425 => "0000000010011000000101",
			2426 => "0011100011010100001000",
			2427 => "0010111001011100000100",
			2428 => "1111111010011000000101",
			2429 => "0000000010011000000101",
			2430 => "0011011100111000000100",
			2431 => "0000001010011000000101",
			2432 => "0000000010011000000101",
			2433 => "0001101001100101100000",
			2434 => "0011110000010001010100",
			2435 => "0001101011001100100100",
			2436 => "0010010101010000010100",
			2437 => "0001101101011000001100",
			2438 => "0000010110101000000100",
			2439 => "1101001010011111000001",
			2440 => "0010011001011000000100",
			2441 => "1101011010011111000001",
			2442 => "1101001010011111000001",
			2443 => "0000110100000100000100",
			2444 => "1101001010011111000001",
			2445 => "1101010010011111000001",
			2446 => "0010100010101100001100",
			2447 => "0010111011011100001000",
			2448 => "0000101100000000000100",
			2449 => "1101010010011111000001",
			2450 => "1110010010011111000001",
			2451 => "1101001010011111000001",
			2452 => "1101001010011111000001",
			2453 => "0011000100000000011000",
			2454 => "0011010011100000001100",
			2455 => "0001010111001000000100",
			2456 => "1101001010011111000001",
			2457 => "0000011001111000000100",
			2458 => "1101110010011111000001",
			2459 => "1101001010011111000001",
			2460 => "0000101100010000001000",
			2461 => "0000110000011100000100",
			2462 => "1110000010011111000001",
			2463 => "1110110010011111000001",
			2464 => "1101001010011111000001",
			2465 => "0010100010101100001000",
			2466 => "0011000100011000000100",
			2467 => "1101101010011111000001",
			2468 => "1101001010011111000001",
			2469 => "0011001011000000001000",
			2470 => "0000101001010000000100",
			2471 => "1101010010011111000001",
			2472 => "1101001010011111000001",
			2473 => "0000111111010100000100",
			2474 => "1101100010011111000001",
			2475 => "1101001010011111000001",
			2476 => "0011000100011000000100",
			2477 => "1101111010011111000001",
			2478 => "0001001000101000000100",
			2479 => "1101001010011111000001",
			2480 => "1101100010011111000001",
			2481 => "0011001001110101010100",
			2482 => "0001100100111100101100",
			2483 => "0000101111010100011000",
			2484 => "0011001001110000001100",
			2485 => "0001011010111100000100",
			2486 => "1101010010011111000001",
			2487 => "0001101001100100000100",
			2488 => "1110011010011111000001",
			2489 => "1110110010011111000001",
			2490 => "0000010111100100001000",
			2491 => "0000010111100100000100",
			2492 => "1101010010011111000001",
			2493 => "1101001010011111000001",
			2494 => "1101101010011111000001",
			2495 => "0010111100101100000100",
			2496 => "1101110010011111000001",
			2497 => "0011111011101100001000",
			2498 => "0001000011000000000100",
			2499 => "1101001010011111000001",
			2500 => "1101001010011111000001",
			2501 => "0010000101000100000100",
			2502 => "1101010010011111000001",
			2503 => "1110011010011111000001",
			2504 => "0001010010011100011100",
			2505 => "0010000001010100001100",
			2506 => "0010111011011100000100",
			2507 => "1110001010011111000001",
			2508 => "0011010100101000000100",
			2509 => "1101011010011111000001",
			2510 => "1101001010011111000001",
			2511 => "0001001001000000001000",
			2512 => "0001101000010000000100",
			2513 => "1110011010011111000001",
			2514 => "1110110010011111000001",
			2515 => "0011001100110000000100",
			2516 => "1110011010011111000001",
			2517 => "1101001010011111000001",
			2518 => "0000100011110000001000",
			2519 => "0001101000010000000100",
			2520 => "1101100010011111000001",
			2521 => "1101001010011111000001",
			2522 => "1110000010011111000001",
			2523 => "0011000001101000010000",
			2524 => "0001100101010000001100",
			2525 => "0001100100111100001000",
			2526 => "0000011100011000000100",
			2527 => "1101101010011111000001",
			2528 => "1101001010011111000001",
			2529 => "1101001010011111000001",
			2530 => "1110001010011111000001",
			2531 => "0010011000010100010100",
			2532 => "0011011100010100000100",
			2533 => "1101100010011111000001",
			2534 => "0001101111000000001000",
			2535 => "0000011100011000000100",
			2536 => "1101011010011111000001",
			2537 => "1101001010011111000001",
			2538 => "0010110001001000000100",
			2539 => "1101001010011111000001",
			2540 => "1101001010011111000001",
			2541 => "0000111110111000000100",
			2542 => "1101001010011111000001",
			2543 => "1101111010011111000001",
			2544 => "0000101110000010100000",
			2545 => "0000100110111101000000",
			2546 => "0000110001101000010100",
			2547 => "0010100001010100001000",
			2548 => "0000010111100100000100",
			2549 => "1111111010100110000101",
			2550 => "0000000010100110000101",
			2551 => "0010001111000100001000",
			2552 => "0001011010111100000100",
			2553 => "0000000010100110000101",
			2554 => "0000000010100110000101",
			2555 => "0000000010100110000101",
			2556 => "0000001111000100011000",
			2557 => "0000010111100100001000",
			2558 => "0000101100010100000100",
			2559 => "0000000010100110000101",
			2560 => "1111111010100110000101",
			2561 => "0001010100000100001000",
			2562 => "0000011101101000000100",
			2563 => "0000000010100110000101",
			2564 => "0000000010100110000101",
			2565 => "0011000100011000000100",
			2566 => "0000000010100110000101",
			2567 => "0000000010100110000101",
			2568 => "0011100010001000010000",
			2569 => "0000100010000100001000",
			2570 => "0011001000111000000100",
			2571 => "0000000010100110000101",
			2572 => "1111111010100110000101",
			2573 => "0001101111000000000100",
			2574 => "0000000010100110000101",
			2575 => "0000000010100110000101",
			2576 => "0000001010100110000101",
			2577 => "0000010001111000111000",
			2578 => "0000000000111000011100",
			2579 => "0001001100001100010000",
			2580 => "0000100000010000001000",
			2581 => "0001010001101000000100",
			2582 => "0000000010100110000101",
			2583 => "1111111010100110000101",
			2584 => "0011101111100100000100",
			2585 => "0000000010100110000101",
			2586 => "0000000010100110000101",
			2587 => "0010111101111000000100",
			2588 => "0000000010100110000101",
			2589 => "0010101100011100000100",
			2590 => "1111111010100110000101",
			2591 => "0000000010100110000101",
			2592 => "0001100100111100001100",
			2593 => "0000101111010100001000",
			2594 => "0011000100000000000100",
			2595 => "0000000010100110000101",
			2596 => "0000000010100110000101",
			2597 => "1111111010100110000101",
			2598 => "0001110110000100001000",
			2599 => "0000101010000100000100",
			2600 => "0000000010100110000101",
			2601 => "0000001010100110000101",
			2602 => "0000111001011100000100",
			2603 => "1111111010100110000101",
			2604 => "0000000010100110000101",
			2605 => "0011001010111000001100",
			2606 => "0011101100010000000100",
			2607 => "0000000010100110000101",
			2608 => "0000010100110100000100",
			2609 => "0000001010100110000101",
			2610 => "0000000010100110000101",
			2611 => "0000001010101100001100",
			2612 => "0011101100111000001000",
			2613 => "0010000101000100000100",
			2614 => "0000000010100110000101",
			2615 => "0000000010100110000101",
			2616 => "0000000010100110000101",
			2617 => "0010110100010000001000",
			2618 => "0010000001010100000100",
			2619 => "0000000010100110000101",
			2620 => "0000001010100110000101",
			2621 => "0010110001001000000100",
			2622 => "0000000010100110000101",
			2623 => "0000000010100110000101",
			2624 => "0010100110011100101100",
			2625 => "0010110100010000001000",
			2626 => "0001010010110100000100",
			2627 => "0000000010100110000101",
			2628 => "0000001010100110000101",
			2629 => "0001000010100100011100",
			2630 => "0010110110100000010000",
			2631 => "0001010111111100001000",
			2632 => "0000100101000000000100",
			2633 => "0000000010100110000101",
			2634 => "0000000010100110000101",
			2635 => "0001110101110100000100",
			2636 => "1111111010100110000101",
			2637 => "0000000010100110000101",
			2638 => "0010001001101000001000",
			2639 => "0000111100001100000100",
			2640 => "0000000010100110000101",
			2641 => "0000000010100110000101",
			2642 => "0000000010100110000101",
			2643 => "0000000000111000000100",
			2644 => "0000001010100110000101",
			2645 => "0000000010100110000101",
			2646 => "0010100101000100000100",
			2647 => "1111111010100110000101",
			2648 => "0011000101100100010000",
			2649 => "0001010010011100001000",
			2650 => "0010110001101000000100",
			2651 => "0000000010100110000101",
			2652 => "1111111010100110000101",
			2653 => "0000010100110100000100",
			2654 => "0000000010100110000101",
			2655 => "0000001010100110000101",
			2656 => "0000000010100110000101",
			2657 => "0000111011000000010000",
			2658 => "0001101001100100000100",
			2659 => "1111111010101011111011",
			2660 => "0001000001001100000100",
			2661 => "0000000010101011111011",
			2662 => "0000101111100100000100",
			2663 => "0000001010101011111011",
			2664 => "0000000010101011111011",
			2665 => "0001100100111101100000",
			2666 => "0011001000111100100100",
			2667 => "0001101101011000000100",
			2668 => "1111111010101011111011",
			2669 => "0000100010000100010000",
			2670 => "0000101100010100001000",
			2671 => "0011100110100100000100",
			2672 => "0000001010101011111011",
			2673 => "1111111010101011111011",
			2674 => "0001010111001000000100",
			2675 => "0000000010101011111011",
			2676 => "0000001010101011111011",
			2677 => "0001101001100100001000",
			2678 => "0010110110000100000100",
			2679 => "0000000010101011111011",
			2680 => "1111110010101011111011",
			2681 => "0000010110101000000100",
			2682 => "0000000010101011111011",
			2683 => "0000001010101011111011",
			2684 => "0001001111101000011100",
			2685 => "0001101100011000001100",
			2686 => "0010010101011100001000",
			2687 => "0011001100110000000100",
			2688 => "0000000010101011111011",
			2689 => "0000001010101011111011",
			2690 => "1111111010101011111011",
			2691 => "0001101101011000001000",
			2692 => "0011000100011000000100",
			2693 => "0000000010101011111011",
			2694 => "0000001010101011111011",
			2695 => "0000001111001000000100",
			2696 => "0000000010101011111011",
			2697 => "0000001010101011111011",
			2698 => "0010111110001100010000",
			2699 => "0000110001011000001000",
			2700 => "0011111001010000000100",
			2701 => "0000000010101011111011",
			2702 => "1111111010101011111011",
			2703 => "0011111110010000000100",
			2704 => "0000001010101011111011",
			2705 => "0000000010101011111011",
			2706 => "0011100111010100001000",
			2707 => "0011001000111000000100",
			2708 => "0000000010101011111011",
			2709 => "1111111010101011111011",
			2710 => "0001011111010000000100",
			2711 => "0000000010101011111011",
			2712 => "1111111010101011111011",
			2713 => "0001010001000000011000",
			2714 => "0001000111011100001100",
			2715 => "0011100011001000001000",
			2716 => "0010110001111100000100",
			2717 => "0000001010101011111011",
			2718 => "0000000010101011111011",
			2719 => "0000001010101011111011",
			2720 => "0010010001000100000100",
			2721 => "0000001010101011111011",
			2722 => "0001001100111100000100",
			2723 => "0000000010101011111011",
			2724 => "1111111010101011111011",
			2725 => "0011111000000100011000",
			2726 => "0010010011101000010000",
			2727 => "0011111110000000001000",
			2728 => "0000011010011000000100",
			2729 => "1111111010101011111011",
			2730 => "0000000010101011111011",
			2731 => "0010110001001000000100",
			2732 => "0000000010101011111011",
			2733 => "0000000010101011111011",
			2734 => "0000111011110000000100",
			2735 => "0000001010101011111011",
			2736 => "1111111010101011111011",
			2737 => "0010000001010100010000",
			2738 => "0010110000110100001000",
			2739 => "0010010011101000000100",
			2740 => "0001111010101011111011",
			2741 => "0000000010101011111011",
			2742 => "0000111100001100000100",
			2743 => "1111111010101011111011",
			2744 => "0000011010101011111011",
			2745 => "0000001011000100001000",
			2746 => "0000011010011000000100",
			2747 => "0000001010101011111011",
			2748 => "0000000010101011111011",
			2749 => "1111111010101011111011",
			2750 => "0000111001110100100000",
			2751 => "0001000010010000001000",
			2752 => "0011011000011000000100",
			2753 => "1111111010101111001101",
			2754 => "0000000010101111001101",
			2755 => "0011101001110000010000",
			2756 => "0000100000010000000100",
			2757 => "1111111010101111001101",
			2758 => "0000100000010000001000",
			2759 => "0010101000110000000100",
			2760 => "0000000010101111001101",
			2761 => "0000000010101111001101",
			2762 => "0000000010101111001101",
			2763 => "0001010100011000000100",
			2764 => "0000001010101111001101",
			2765 => "0000000010101111001101",
			2766 => "0000100110010000101000",
			2767 => "0000011001111000001000",
			2768 => "0011101011000000000100",
			2769 => "0000001010101111001101",
			2770 => "0000000010101111001101",
			2771 => "0000110000011100001100",
			2772 => "0000000011010000000100",
			2773 => "1111111010101111001101",
			2774 => "0000111000011000000100",
			2775 => "1111111010101111001101",
			2776 => "0000000010101111001101",
			2777 => "0000001111000100010000",
			2778 => "0000010111100100001000",
			2779 => "0011000100000000000100",
			2780 => "0000000010101111001101",
			2781 => "1111111010101111001101",
			2782 => "0001001100010000000100",
			2783 => "0000000010101111001101",
			2784 => "0000001010101111001101",
			2785 => "0000001010101111001101",
			2786 => "0001011010111000001000",
			2787 => "0000100010000100000100",
			2788 => "0000000010101111001101",
			2789 => "1111111010101111001101",
			2790 => "0010001111000100011000",
			2791 => "0001010100011000001100",
			2792 => "0000000011111100000100",
			2793 => "1111111010101111001101",
			2794 => "0001101011001100000100",
			2795 => "0000000010101111001101",
			2796 => "0000001010101111001101",
			2797 => "0011011000000000000100",
			2798 => "1111111010101111001101",
			2799 => "0001000010111000000100",
			2800 => "0000000010101111001101",
			2801 => "0000000010101111001101",
			2802 => "1111111010101111001101",
			2803 => "0000111001110100100000",
			2804 => "0001101011001100001000",
			2805 => "0000010111100100000100",
			2806 => "1111111010110011010001",
			2807 => "0000000010110011010001",
			2808 => "0010011011101000010000",
			2809 => "0001010100001000000100",
			2810 => "0000000010110011010001",
			2811 => "0011110110100000001000",
			2812 => "0000000100011000000100",
			2813 => "0000001010110011010001",
			2814 => "0000000010110011010001",
			2815 => "0000000010110011010001",
			2816 => "0000011001111000000100",
			2817 => "1111111010110011010001",
			2818 => "0000000010110011010001",
			2819 => "0011110101001000100000",
			2820 => "0010001111001000010000",
			2821 => "0000110100000100000100",
			2822 => "1111111010110011010001",
			2823 => "0011110001000000001000",
			2824 => "0011111110101000000100",
			2825 => "0000000010110011010001",
			2826 => "0000001010110011010001",
			2827 => "0000000010110011010001",
			2828 => "0000110001101000001000",
			2829 => "0000011001111000000100",
			2830 => "0000001010110011010001",
			2831 => "1111111010110011010001",
			2832 => "0010111100101100000100",
			2833 => "0000001010110011010001",
			2834 => "0000000010110011010001",
			2835 => "0000110010001000100000",
			2836 => "0010111100101100010100",
			2837 => "0011111110010000010000",
			2838 => "0001101011001100001000",
			2839 => "0010110101101100000100",
			2840 => "0000000010110011010001",
			2841 => "1111111010110011010001",
			2842 => "0000110001011000000100",
			2843 => "0000000010110011010001",
			2844 => "0000001010110011010001",
			2845 => "1111111010110011010001",
			2846 => "0000101100010000000100",
			2847 => "1111110010110011010001",
			2848 => "0001101111000000000100",
			2849 => "1111111010110011010001",
			2850 => "0000000010110011010001",
			2851 => "0000010110101000001000",
			2852 => "0000001110111100000100",
			2853 => "1111111010110011010001",
			2854 => "0000000010110011010001",
			2855 => "0001011000000000001100",
			2856 => "0011110010000000001000",
			2857 => "0001010100011000000100",
			2858 => "0000000010110011010001",
			2859 => "0000001010110011010001",
			2860 => "0000000010110011010001",
			2861 => "0000010000111100001000",
			2862 => "0001101111000000000100",
			2863 => "0000000010110011010001",
			2864 => "0000000010110011010001",
			2865 => "0001001000001000000100",
			2866 => "0000000010110011010001",
			2867 => "0000000010110011010001",
			2868 => "0001111001110000110100",
			2869 => "0011110010011100100000",
			2870 => "0000110000011100011100",
			2871 => "0001000100001100001000",
			2872 => "0000111010001100000100",
			2873 => "1111111010110111001101",
			2874 => "0000000010110111001101",
			2875 => "0010110011011100001000",
			2876 => "0000111010111100000100",
			2877 => "0000000010110111001101",
			2878 => "0000000010110111001101",
			2879 => "0011110101001000001000",
			2880 => "0001101101011000000100",
			2881 => "0000000010110111001101",
			2882 => "0000001010110111001101",
			2883 => "0000000010110111001101",
			2884 => "0000001010110111001101",
			2885 => "0000110101110100010000",
			2886 => "0011100100000100001100",
			2887 => "0000011001111000001000",
			2888 => "0001000010100100000100",
			2889 => "0000000010110111001101",
			2890 => "0000000010110111001101",
			2891 => "0000000010110111001101",
			2892 => "1111111010110111001101",
			2893 => "0000000010110111001101",
			2894 => "0001111001110000010000",
			2895 => "0000111000011000001000",
			2896 => "0011001100001000000100",
			2897 => "0000000010110111001101",
			2898 => "0000000010110111001101",
			2899 => "0010001001101000000100",
			2900 => "0000000010110111001101",
			2901 => "0000001010110111001101",
			2902 => "0011011000000000001000",
			2903 => "0001000010010000000100",
			2904 => "1111111010110111001101",
			2905 => "0000000010110111001101",
			2906 => "0001011000000000010100",
			2907 => "0001101001100100001000",
			2908 => "0011000100000000000100",
			2909 => "0000000010110111001101",
			2910 => "0000000010110111001101",
			2911 => "0000000011111100001000",
			2912 => "0011111110010000000100",
			2913 => "0000000010110111001101",
			2914 => "0000000010110111001101",
			2915 => "0000001010110111001101",
			2916 => "0011001101010100010000",
			2917 => "0010101010110000001000",
			2918 => "0001001000000100000100",
			2919 => "0000000010110111001101",
			2920 => "1111111010110111001101",
			2921 => "0001110110000100000100",
			2922 => "0000000010110111001101",
			2923 => "0000000010110111001101",
			2924 => "0001000101010100001000",
			2925 => "0010000001110000000100",
			2926 => "0000000010110111001101",
			2927 => "0000000010110111001101",
			2928 => "0011111100001100000100",
			2929 => "0000000010110111001101",
			2930 => "0000000010110111001101",
			2931 => "0010110011011100001100",
			2932 => "0001000110110000000100",
			2933 => "1111111010111010001001",
			2934 => "0000000110000100000100",
			2935 => "0000000010111010001001",
			2936 => "0000000010111010001001",
			2937 => "0001111000111000010000",
			2938 => "0001101011001100000100",
			2939 => "0000000010111010001001",
			2940 => "0001111000111100001000",
			2941 => "0001110100000000000100",
			2942 => "0000000010111010001001",
			2943 => "0000000010111010001001",
			2944 => "0000001010111010001001",
			2945 => "0001111001110000001000",
			2946 => "0001001000000100000100",
			2947 => "0000000010111010001001",
			2948 => "1111111010111010001001",
			2949 => "0011010111111100011100",
			2950 => "0011101011101100010000",
			2951 => "0010101010110000001000",
			2952 => "0001001000000100000100",
			2953 => "0000000010111010001001",
			2954 => "1111111010111010001001",
			2955 => "0010011001011000000100",
			2956 => "0000000010111010001001",
			2957 => "0000000010111010001001",
			2958 => "0001010101001000001000",
			2959 => "0000010111101000000100",
			2960 => "0000000010111010001001",
			2961 => "0000001010111010001001",
			2962 => "0000000010111010001001",
			2963 => "0001011001010000010000",
			2964 => "0011011110010000001000",
			2965 => "0011101111101000000100",
			2966 => "0000000010111010001001",
			2967 => "0000000010111010001001",
			2968 => "0000111110000000000100",
			2969 => "1111111010111010001001",
			2970 => "0000000010111010001001",
			2971 => "0010000001010100001000",
			2972 => "0001110100010000000100",
			2973 => "0000000010111010001001",
			2974 => "0000000010111010001001",
			2975 => "0010110101110100000100",
			2976 => "0000000010111010001001",
			2977 => "0000000010111010001001",
			2978 => "0001010111001000010100",
			2979 => "0001000001101100001000",
			2980 => "0000111000011000000100",
			2981 => "1111111010111110011101",
			2982 => "0000000010111110011101",
			2983 => "0010110011011100001000",
			2984 => "0000110100001000000100",
			2985 => "0000000010111110011101",
			2986 => "0000000010111110011101",
			2987 => "0000000010111110011101",
			2988 => "0011111111010000110100",
			2989 => "0001111001110000011000",
			2990 => "0010101010110000001100",
			2991 => "0011000100000000000100",
			2992 => "1111111010111110011101",
			2993 => "0011000100000000000100",
			2994 => "0000001010111110011101",
			2995 => "0000000010111110011101",
			2996 => "0000111001110100000100",
			2997 => "0000000010111110011101",
			2998 => "0011000100000000000100",
			2999 => "0000001010111110011101",
			3000 => "0000000010111110011101",
			3001 => "0011101011011100010100",
			3002 => "0011111100100100001000",
			3003 => "0000000001110100000100",
			3004 => "0000000010111110011101",
			3005 => "1111111010111110011101",
			3006 => "0010101100011100000100",
			3007 => "0000000010111110011101",
			3008 => "0011001001110000000100",
			3009 => "0000000010111110011101",
			3010 => "0000000010111110011101",
			3011 => "0001100111101000000100",
			3012 => "0000000010111110011101",
			3013 => "0000001010111110011101",
			3014 => "0010011110010100101000",
			3015 => "0011100101110100011000",
			3016 => "0000110001011000001000",
			3017 => "0001101111000000000100",
			3018 => "1111111010111110011101",
			3019 => "0000000010111110011101",
			3020 => "0011010001101000001000",
			3021 => "0011111110010000000100",
			3022 => "0000000010111110011101",
			3023 => "0000000010111110011101",
			3024 => "0000110111110000000100",
			3025 => "1111111010111110011101",
			3026 => "0000000010111110011101",
			3027 => "0000110001001000000100",
			3028 => "1111111010111110011101",
			3029 => "0010111100101000000100",
			3030 => "0000000010111110011101",
			3031 => "0001100100111100000100",
			3032 => "0000000010111110011101",
			3033 => "1111111010111110011101",
			3034 => "0001011000011000001000",
			3035 => "0000001000110000000100",
			3036 => "0000000010111110011101",
			3037 => "0000001010111110011101",
			3038 => "0000110111100000000100",
			3039 => "1111111010111110011101",
			3040 => "0011011011101100001000",
			3041 => "0011111000110100000100",
			3042 => "0000000010111110011101",
			3043 => "0000000010111110011101",
			3044 => "0011100001101100000100",
			3045 => "1111111010111110011101",
			3046 => "0000000010111110011101",
			3047 => "0001011010111000100100",
			3048 => "0001001111100000001100",
			3049 => "0001111001110000000100",
			3050 => "1111111011000010111001",
			3051 => "0001111101100000000100",
			3052 => "0000000011000010111001",
			3053 => "0000000011000010111001",
			3054 => "0011010001111100000100",
			3055 => "1111111011000010111001",
			3056 => "0011111110000100010000",
			3057 => "0001101011001100001100",
			3058 => "0010100110011100001000",
			3059 => "0010101100011100000100",
			3060 => "0000000011000010111001",
			3061 => "0000000011000010111001",
			3062 => "0000000011000010111001",
			3063 => "0000001011000010111001",
			3064 => "1111111011000010111001",
			3065 => "0001010100011000100000",
			3066 => "0011011011000000010100",
			3067 => "0010110101101100001000",
			3068 => "0010011111001100000100",
			3069 => "0000000011000010111001",
			3070 => "1111111011000010111001",
			3071 => "0001111001110000001000",
			3072 => "0001101101011000000100",
			3073 => "0000000011000010111001",
			3074 => "0000001011000010111001",
			3075 => "0000000011000010111001",
			3076 => "0001101101011000000100",
			3077 => "0000000011000010111001",
			3078 => "0001111101100000000100",
			3079 => "0000001011000010111001",
			3080 => "0000000011000010111001",
			3081 => "0011011000000000011000",
			3082 => "0001000010100100010000",
			3083 => "0011110101110000001100",
			3084 => "0001111001110000000100",
			3085 => "0000000011000010111001",
			3086 => "0000011001111000000100",
			3087 => "0000000011000010111001",
			3088 => "1111111011000010111001",
			3089 => "1111111011000010111001",
			3090 => "0010111100101100000100",
			3091 => "0000000011000010111001",
			3092 => "0000000011000010111001",
			3093 => "0010111100101100010100",
			3094 => "0000000000111000010000",
			3095 => "0011011001001000001000",
			3096 => "0000010110101000000100",
			3097 => "0000000011000010111001",
			3098 => "1111111011000010111001",
			3099 => "0010111100101100000100",
			3100 => "0000000011000010111001",
			3101 => "0000001011000010111001",
			3102 => "0000001011000010111001",
			3103 => "0011100101100100010000",
			3104 => "0000000001110100001000",
			3105 => "0001111100101000000100",
			3106 => "0000000011000010111001",
			3107 => "0000000011000010111001",
			3108 => "0001101111000000000100",
			3109 => "1111111011000010111001",
			3110 => "0000000011000010111001",
			3111 => "0001111101100000001000",
			3112 => "0000010111100100000100",
			3113 => "0000000011000010111001",
			3114 => "0000001011000010111001",
			3115 => "0010011100011000000100",
			3116 => "0000000011000010111001",
			3117 => "0000000011000010111001",
			3118 => "0000000011010000110100",
			3119 => "0000010110101000001000",
			3120 => "0001000010110000000100",
			3121 => "1111111011000111011101",
			3122 => "0000000011000111011101",
			3123 => "0000000011010000101000",
			3124 => "0011000100000000001000",
			3125 => "0001101011001100000100",
			3126 => "0000000011000111011101",
			3127 => "0000001011000111011101",
			3128 => "0001110001111100010000",
			3129 => "0000101001100000001000",
			3130 => "0001001110000000000100",
			3131 => "0000000011000111011101",
			3132 => "0000000011000111011101",
			3133 => "0001101000010000000100",
			3134 => "0000000011000111011101",
			3135 => "0000000011000111011101",
			3136 => "0010001011010100001000",
			3137 => "0011011001011100000100",
			3138 => "0000000011000111011101",
			3139 => "0000000011000111011101",
			3140 => "0011000001101000000100",
			3141 => "0000001011000111011101",
			3142 => "0000000011000111011101",
			3143 => "1111111011000111011101",
			3144 => "0011001100110000111100",
			3145 => "0001101001100100011100",
			3146 => "0000101110110100010000",
			3147 => "0011101110110000001000",
			3148 => "0011100111001000000100",
			3149 => "0000000011000111011101",
			3150 => "0000000011000111011101",
			3151 => "0010101010110000000100",
			3152 => "0000000011000111011101",
			3153 => "0000001011000111011101",
			3154 => "0001000011011000001000",
			3155 => "0001110100000000000100",
			3156 => "0000000011000111011101",
			3157 => "1111111011000111011101",
			3158 => "0000000011000111011101",
			3159 => "0010101001101000011000",
			3160 => "0001100100111100010000",
			3161 => "0000101111010100001000",
			3162 => "0001001000001000000100",
			3163 => "0000000011000111011101",
			3164 => "0000000011000111011101",
			3165 => "0011110011001000000100",
			3166 => "0000000011000111011101",
			3167 => "0000000011000111011101",
			3168 => "0000000011010000000100",
			3169 => "0000000011000111011101",
			3170 => "0000001011000111011101",
			3171 => "0010101111001000000100",
			3172 => "0000000011000111011101",
			3173 => "0000000011000111011101",
			3174 => "0000000000111000001100",
			3175 => "0011001000011000001000",
			3176 => "0001101000010000000100",
			3177 => "0000000011000111011101",
			3178 => "0000000011000111011101",
			3179 => "0000000011000111011101",
			3180 => "0011100011010100010000",
			3181 => "0001000111011100001100",
			3182 => "0010000001110100001000",
			3183 => "0010000111000100000100",
			3184 => "0000000011000111011101",
			3185 => "0000000011000111011101",
			3186 => "0000000011000111011101",
			3187 => "1111111011000111011101",
			3188 => "0001111001010100000100",
			3189 => "0000000011000111011101",
			3190 => "0000000011000111011101",
			3191 => "0000111001110100010100",
			3192 => "0001101011001100001000",
			3193 => "0000010111100100000100",
			3194 => "1111111011001010110001",
			3195 => "0000000011001010110001",
			3196 => "0001111101100000001000",
			3197 => "0010111001110000000100",
			3198 => "0000000011001010110001",
			3199 => "0000001011001010110001",
			3200 => "1111111011001010110001",
			3201 => "0000001001110001010100",
			3202 => "0000000011010000100100",
			3203 => "0000110000011100001000",
			3204 => "0000000011111100000100",
			3205 => "1111111011001010110001",
			3206 => "1111110011001010110001",
			3207 => "0011111001010000001100",
			3208 => "0000000010011000001000",
			3209 => "0001110001111100000100",
			3210 => "0000000011001010110001",
			3211 => "0000001011001010110001",
			3212 => "0000001011001010110001",
			3213 => "0000010111100100001000",
			3214 => "0011110011001000000100",
			3215 => "0000000011001010110001",
			3216 => "1111111011001010110001",
			3217 => "0001010001101000000100",
			3218 => "0000001011001010110001",
			3219 => "0000000011001010110001",
			3220 => "0000001110111100010000",
			3221 => "0010101010110000000100",
			3222 => "1111111011001010110001",
			3223 => "0011001111011100001000",
			3224 => "0001101111000000000100",
			3225 => "0000000011001010110001",
			3226 => "0000001011001010110001",
			3227 => "1111111011001010110001",
			3228 => "0010100101000100010000",
			3229 => "0010000010101000001000",
			3230 => "0010100110011100000100",
			3231 => "1111111011001010110001",
			3232 => "0000000011001010110001",
			3233 => "0011110111111100000100",
			3234 => "0000000011001010110001",
			3235 => "1111111011001010110001",
			3236 => "0011000110000100001000",
			3237 => "0000001000111100000100",
			3238 => "0000001011001010110001",
			3239 => "0000000011001010110001",
			3240 => "0010111110101000000100",
			3241 => "1111111011001010110001",
			3242 => "0000001011001010110001",
			3243 => "1111111011001010110001",
			3244 => "0001111001110000111100",
			3245 => "0011110010011100100100",
			3246 => "0000110000011100100000",
			3247 => "0001000100001100001000",
			3248 => "0000111010001100000100",
			3249 => "1111111011001111110101",
			3250 => "0000000011001111110101",
			3251 => "0010110011011100001100",
			3252 => "0000100111011000001000",
			3253 => "0001111000111000000100",
			3254 => "0000000011001111110101",
			3255 => "0000000011001111110101",
			3256 => "0000000011001111110101",
			3257 => "0011110101001000001000",
			3258 => "0001101101011000000100",
			3259 => "0000000011001111110101",
			3260 => "0000001011001111110101",
			3261 => "0000000011001111110101",
			3262 => "0000001011001111110101",
			3263 => "0000110101110100010100",
			3264 => "0000010110101000010000",
			3265 => "0001111000111000001100",
			3266 => "0001001010110100000100",
			3267 => "0000000011001111110101",
			3268 => "0001000011010100000100",
			3269 => "0000000011001111110101",
			3270 => "0000000011001111110101",
			3271 => "0000000011001111110101",
			3272 => "1111111011001111110101",
			3273 => "0000000011001111110101",
			3274 => "0001111001110000011000",
			3275 => "0000000000110000001100",
			3276 => "0001101101011000000100",
			3277 => "0000000011001111110101",
			3278 => "0010111110001100000100",
			3279 => "0000001011001111110101",
			3280 => "0000000011001111110101",
			3281 => "0001010111001000001000",
			3282 => "0001011101010100000100",
			3283 => "0000000011001111110101",
			3284 => "0000000011001111110101",
			3285 => "0000000011001111110101",
			3286 => "0000111011011100011100",
			3287 => "0010100110011100001100",
			3288 => "0001111100101000001000",
			3289 => "0010110110000100000100",
			3290 => "0000000011001111110101",
			3291 => "1111111011001111110101",
			3292 => "0000000011001111110101",
			3293 => "0000111001110100001000",
			3294 => "0011010100011000000100",
			3295 => "0000000011001111110101",
			3296 => "0000000011001111110101",
			3297 => "0001111101100000000100",
			3298 => "0000000011001111110101",
			3299 => "0000000011001111110101",
			3300 => "0001011001110100010100",
			3301 => "0000000011111100001100",
			3302 => "0000010111100100000100",
			3303 => "0000000011001111110101",
			3304 => "0001101001100100000100",
			3305 => "0000000011001111110101",
			3306 => "0000001011001111110101",
			3307 => "0001000000010100000100",
			3308 => "0000001011001111110101",
			3309 => "0000000011001111110101",
			3310 => "0010111010111000010000",
			3311 => "0001101000010000001000",
			3312 => "0010110000001100000100",
			3313 => "0000000011001111110101",
			3314 => "1111111011001111110101",
			3315 => "0010110001111100000100",
			3316 => "0000000011001111110101",
			3317 => "0000000011001111110101",
			3318 => "0000000010011000001000",
			3319 => "0001010001000000000100",
			3320 => "0000000011001111110101",
			3321 => "0000000011001111110101",
			3322 => "0010101010110000000100",
			3323 => "1111111011001111110101",
			3324 => "0000000011001111110101",
			3325 => "0001100100111101011100",
			3326 => "0001110001101001010100",
			3327 => "0000011101101000111000",
			3328 => "0001010011100000100000",
			3329 => "0011011011000000010000",
			3330 => "0011001100001000001000",
			3331 => "0001011010111100000100",
			3332 => "0000000011010100011001",
			3333 => "0000000011010100011001",
			3334 => "0010000001110100000100",
			3335 => "1111111011010100011001",
			3336 => "0000000011010100011001",
			3337 => "0011000100000000001000",
			3338 => "0001111001110000000100",
			3339 => "1111111011010100011001",
			3340 => "0000000011010100011001",
			3341 => "0001111101100000000100",
			3342 => "0000001011010100011001",
			3343 => "0000000011010100011001",
			3344 => "0011000100000000001100",
			3345 => "0010101010110000001000",
			3346 => "0010010101011100000100",
			3347 => "0000000011010100011001",
			3348 => "0000000011010100011001",
			3349 => "0000000011010100011001",
			3350 => "0001101111000000001000",
			3351 => "0000010111100100000100",
			3352 => "1111111011010100011001",
			3353 => "0000000011010100011001",
			3354 => "0000000011010100011001",
			3355 => "0011100111010100010100",
			3356 => "0011000100011000001100",
			3357 => "0011101011011100000100",
			3358 => "0000000011010100011001",
			3359 => "0010011010100000000100",
			3360 => "0000000011010100011001",
			3361 => "0000000011010100011001",
			3362 => "0001010110100000000100",
			3363 => "0000000011010100011001",
			3364 => "0000000011010100011001",
			3365 => "0010101000100100000100",
			3366 => "0000000011010100011001",
			3367 => "0000000011010100011001",
			3368 => "0001110101100100000100",
			3369 => "1111111011010100011001",
			3370 => "0000000011010100011001",
			3371 => "0001011010011100001100",
			3372 => "0011000000101000000100",
			3373 => "0000000011010100011001",
			3374 => "0000101100000000000100",
			3375 => "0000000011010100011001",
			3376 => "0000001011010100011001",
			3377 => "0010011100011000001100",
			3378 => "0000110010000000000100",
			3379 => "1111111011010100011001",
			3380 => "0000011101101000000100",
			3381 => "0000000011010100011001",
			3382 => "0000000011010100011001",
			3383 => "0001011010010100001000",
			3384 => "0011000011011100000100",
			3385 => "0000000011010100011001",
			3386 => "0000001011010100011001",
			3387 => "0011101111100100001000",
			3388 => "0010010111101100000100",
			3389 => "1111111011010100011001",
			3390 => "0000000011010100011001",
			3391 => "0000001111000100001000",
			3392 => "0010101000100100000100",
			3393 => "0000000011010100011001",
			3394 => "0000000011010100011001",
			3395 => "0010100001010000000100",
			3396 => "1111111011010100011001",
			3397 => "0000000011010100011001",
			3398 => "0001101011001101010000",
			3399 => "0010011000010000110000",
			3400 => "0001101101011000010100",
			3401 => "0000010110101000000100",
			3402 => "1111111011011001100101",
			3403 => "0000000001110000000100",
			3404 => "1111111011011001100101",
			3405 => "0011110010000100001000",
			3406 => "0011001110001100000100",
			3407 => "0000000011011001100101",
			3408 => "0000101011011001100101",
			3409 => "1111111011011001100101",
			3410 => "0000111001110100000100",
			3411 => "1111111011011001100101",
			3412 => "0011110001000000001100",
			3413 => "0011001000111100001000",
			3414 => "0000000000111000000100",
			3415 => "0000001011011001100101",
			3416 => "0000011011011001100101",
			3417 => "0000000011011001100101",
			3418 => "0010011111000000001000",
			3419 => "0000101110110100000100",
			3420 => "0000000011011001100101",
			3421 => "1111111011011001100101",
			3422 => "0000011011011001100101",
			3423 => "0000100000010000011100",
			3424 => "0010101010100000000100",
			3425 => "0000010011011001100101",
			3426 => "0011100110010000001000",
			3427 => "0011110110010000000100",
			3428 => "0000001011011001100101",
			3429 => "1111111011011001100101",
			3430 => "0011011111010000001000",
			3431 => "0000010001111000000100",
			3432 => "0000010011011001100101",
			3433 => "1111111011011001100101",
			3434 => "0011000100011000000100",
			3435 => "0000000011011001100101",
			3436 => "1111111011011001100101",
			3437 => "0000010011011001100101",
			3438 => "0011000001101000110100",
			3439 => "0010101000010100011000",
			3440 => "0000011011111100000100",
			3441 => "0000010011011001100101",
			3442 => "0011010001000000001000",
			3443 => "0011100110111100000100",
			3444 => "1111111011011001100101",
			3445 => "0000000011011001100101",
			3446 => "0000001111001000000100",
			3447 => "1111111011011001100101",
			3448 => "0001000001011100000100",
			3449 => "0000101011011001100101",
			3450 => "0000000011011001100101",
			3451 => "0001000011111000010100",
			3452 => "0001011101010100001000",
			3453 => "0001001101110100000100",
			3454 => "1111111011011001100101",
			3455 => "0000001011011001100101",
			3456 => "0000001010101100000100",
			3457 => "0000000011011001100101",
			3458 => "0001010111111100000100",
			3459 => "0000001011011001100101",
			3460 => "0000000011011001100101",
			3461 => "0001101111000000000100",
			3462 => "1111111011011001100101",
			3463 => "0000001011011001100101",
			3464 => "0010011000010100011100",
			3465 => "0001010111111100001000",
			3466 => "0001010010011100000100",
			3467 => "1111111011011001100101",
			3468 => "0000001011011001100101",
			3469 => "0001101111000000000100",
			3470 => "0000001011011001100101",
			3471 => "0011010110111100001000",
			3472 => "0000010101011100000100",
			3473 => "0000000011011001100101",
			3474 => "1111111011011001100101",
			3475 => "0010101010110000000100",
			3476 => "0000000011011001100101",
			3477 => "1111111011011001100101",
			3478 => "0000110100001100000100",
			3479 => "1111111011011001100101",
			3480 => "0000010011011001100101",
			3481 => "0000111001110100011000",
			3482 => "0010100001010100001000",
			3483 => "0000010111100100000100",
			3484 => "1111111011011101010001",
			3485 => "0000000011011101010001",
			3486 => "0001111101100000001100",
			3487 => "0010111001110000001000",
			3488 => "0010110100000000000100",
			3489 => "1111111011011101010001",
			3490 => "0000000011011101010001",
			3491 => "0000001011011101010001",
			3492 => "1111111011011101010001",
			3493 => "0000001001110001011100",
			3494 => "0011010110111100111100",
			3495 => "0001010001000000011100",
			3496 => "0001110001101000010000",
			3497 => "0000000011010000001000",
			3498 => "0000110000011100000100",
			3499 => "1111111011011101010001",
			3500 => "0000000011011101010001",
			3501 => "0000001010000000000100",
			3502 => "0000000011011101010001",
			3503 => "0000000011011101010001",
			3504 => "0011111010000100000100",
			3505 => "1111111011011101010001",
			3506 => "0010111011011100000100",
			3507 => "0000001011011101010001",
			3508 => "0000000011011101010001",
			3509 => "0000110010010100010000",
			3510 => "0001010101110000001000",
			3511 => "0001111000011000000100",
			3512 => "0000000011011101010001",
			3513 => "1111111011011101010001",
			3514 => "0000011110010100000100",
			3515 => "0000000011011101010001",
			3516 => "1111111011011101010001",
			3517 => "0011101000101000001000",
			3518 => "0001001110000000000100",
			3519 => "0000000011011101010001",
			3520 => "0000001011011101010001",
			3521 => "0000110110111000000100",
			3522 => "1111111011011101010001",
			3523 => "0000000011011101010001",
			3524 => "0001110110110100001000",
			3525 => "0001111011011100000100",
			3526 => "0000001011011101010001",
			3527 => "0000010011011101010001",
			3528 => "0010010111101100001100",
			3529 => "0001011110110100000100",
			3530 => "0000000011011101010001",
			3531 => "0000000011010000000100",
			3532 => "0000001011011101010001",
			3533 => "0000000011011101010001",
			3534 => "0010111111010000001000",
			3535 => "0011001010001100000100",
			3536 => "0000000011011101010001",
			3537 => "1111111011011101010001",
			3538 => "0000001011011101010001",
			3539 => "1111111011011101010001",
			3540 => "0010001001000100011100",
			3541 => "0001110001101000011000",
			3542 => "0001111100101000000100",
			3543 => "0000000011100000101101",
			3544 => "0010111011011100010000",
			3545 => "0010000010101100000100",
			3546 => "0000000011100000101101",
			3547 => "0011010101110000001000",
			3548 => "0001010111100000000100",
			3549 => "0000000011100000101101",
			3550 => "0000000011100000101101",
			3551 => "0000000011100000101101",
			3552 => "0000000011100000101101",
			3553 => "0000000011100000101101",
			3554 => "0001101010011000000100",
			3555 => "1111111011100000101101",
			3556 => "0010111100110000010100",
			3557 => "0011011110110000010000",
			3558 => "0001111000111000001000",
			3559 => "0001111100001000000100",
			3560 => "0000000011100000101101",
			3561 => "0000000011100000101101",
			3562 => "0001111001110000000100",
			3563 => "0000000011100000101101",
			3564 => "0000000011100000101101",
			3565 => "0000001011100000101101",
			3566 => "0000110111110000011100",
			3567 => "0001000011110000001100",
			3568 => "0000010110101000000100",
			3569 => "1111111011100000101101",
			3570 => "0001001000000100000100",
			3571 => "1111111011100000101101",
			3572 => "0000000011100000101101",
			3573 => "0000111010011100001000",
			3574 => "0000100110111100000100",
			3575 => "0000000011100000101101",
			3576 => "0000000011100000101101",
			3577 => "0000100010000100000100",
			3578 => "0000001011100000101101",
			3579 => "0000000011100000101101",
			3580 => "0011110110010000010000",
			3581 => "0010110000001100001000",
			3582 => "0011101001010100000100",
			3583 => "0000001011100000101101",
			3584 => "0000000011100000101101",
			3585 => "0001110001111100000100",
			3586 => "0000000011100000101101",
			3587 => "0000000011100000101101",
			3588 => "0010000111000100001000",
			3589 => "0001000011101100000100",
			3590 => "0000000011100000101101",
			3591 => "0000000011100000101101",
			3592 => "0011100011010100000100",
			3593 => "0000000011100000101101",
			3594 => "0000000011100000101101",
			3595 => "0000110110111001111100",
			3596 => "0011011001011101011100",
			3597 => "0000111011111000111100",
			3598 => "0000100110010000011100",
			3599 => "0000101100010100010000",
			3600 => "0011100010001000001000",
			3601 => "0001101001011000000100",
			3602 => "0000000011100101111001",
			3603 => "0000000011100101111001",
			3604 => "0010111000000000000100",
			3605 => "0000000011100101111001",
			3606 => "0000000011100101111001",
			3607 => "0011000100010100000100",
			3608 => "0000000011100101111001",
			3609 => "0011000100000000000100",
			3610 => "0000001011100101111001",
			3611 => "0000000011100101111001",
			3612 => "0000000011010000010000",
			3613 => "0001110111001000001000",
			3614 => "0011001000111000000100",
			3615 => "0000000011100101111001",
			3616 => "1111111011100101111001",
			3617 => "0010001100011100000100",
			3618 => "0000000011100101111001",
			3619 => "0000000011100101111001",
			3620 => "0000000011010000001000",
			3621 => "0010101010110000000100",
			3622 => "0000000011100101111001",
			3623 => "0000001011100101111001",
			3624 => "0000111100010100000100",
			3625 => "0000000011100101111001",
			3626 => "0000000011100101111001",
			3627 => "0000000001110100010000",
			3628 => "0000111100111000001100",
			3629 => "0001000001011100000100",
			3630 => "0000000011100101111001",
			3631 => "0011001011000000000100",
			3632 => "0000000011100101111001",
			3633 => "0000000011100101111001",
			3634 => "0000000011100101111001",
			3635 => "0010010010101100001100",
			3636 => "0001101001111100001000",
			3637 => "0010110010001000000100",
			3638 => "0000001011100101111001",
			3639 => "0000000011100101111001",
			3640 => "0000000011100101111001",
			3641 => "0000000011100101111001",
			3642 => "0000100010010100010100",
			3643 => "0010110101110100001000",
			3644 => "0011001001110100000100",
			3645 => "0000000011100101111001",
			3646 => "0000000011100101111001",
			3647 => "0011000001101000001000",
			3648 => "0000001011010100000100",
			3649 => "0000000011100101111001",
			3650 => "0000000011100101111001",
			3651 => "0000000011100101111001",
			3652 => "0010010111101100000100",
			3653 => "0000000011100101111001",
			3654 => "0011011010001000000100",
			3655 => "0000000011100101111001",
			3656 => "1111111011100101111001",
			3657 => "0011011100111000100100",
			3658 => "0011111000110100001100",
			3659 => "0000000001110100000100",
			3660 => "0000000011100101111001",
			3661 => "0000110110111000000100",
			3662 => "0000000011100101111001",
			3663 => "0000000011100101111001",
			3664 => "0001110001101000000100",
			3665 => "0000000011100101111001",
			3666 => "0010101000100100000100",
			3667 => "0000000011100101111001",
			3668 => "0010010000001000001000",
			3669 => "0001101001111100000100",
			3670 => "0000000011100101111001",
			3671 => "0000000011100101111001",
			3672 => "0001100100111100000100",
			3673 => "0000000011100101111001",
			3674 => "0000000011100101111001",
			3675 => "0011000101110100000100",
			3676 => "0000000011100101111001",
			3677 => "0000000011100101111001",
			3678 => "0000010100110101110000",
			3679 => "0000100110010000110000",
			3680 => "0000101100010100010000",
			3681 => "0011100010001000001000",
			3682 => "0001101001011000000100",
			3683 => "0000000011101010111101",
			3684 => "0000000011101010111101",
			3685 => "0010111000000000000100",
			3686 => "0000000011101010111101",
			3687 => "0000000011101010111101",
			3688 => "0011000100010100000100",
			3689 => "0000000011101010111101",
			3690 => "0011000100000000001100",
			3691 => "0001101101011000000100",
			3692 => "0000000011101010111101",
			3693 => "0010110011011100000100",
			3694 => "0000000011101010111101",
			3695 => "0000001011101010111101",
			3696 => "0011001000111000001000",
			3697 => "0011011001110100000100",
			3698 => "0000000011101010111101",
			3699 => "0000000011101010111101",
			3700 => "0010011100011000000100",
			3701 => "0000000011101010111101",
			3702 => "0000000011101010111101",
			3703 => "0011011100010000101100",
			3704 => "0011011001011100011100",
			3705 => "0011011001010100010000",
			3706 => "0001111101100000001000",
			3707 => "0001000011110000000100",
			3708 => "0000000011101010111101",
			3709 => "0000000011101010111101",
			3710 => "0001101000010000000100",
			3711 => "1111111011101010111101",
			3712 => "0000000011101010111101",
			3713 => "0000011111001100000100",
			3714 => "0000000011101010111101",
			3715 => "0001000100001100000100",
			3716 => "0000000011101010111101",
			3717 => "0000000011101010111101",
			3718 => "0010010101010000001000",
			3719 => "0000010101011100000100",
			3720 => "0000000011101010111101",
			3721 => "0000000011101010111101",
			3722 => "0011101000110100000100",
			3723 => "1111111011101010111101",
			3724 => "0000000011101010111101",
			3725 => "0011010011000000010000",
			3726 => "0001101001111100001100",
			3727 => "0000010000111100000100",
			3728 => "0000000011101010111101",
			3729 => "0001011100010100000100",
			3730 => "0000000011101010111101",
			3731 => "0000000011101010111101",
			3732 => "0000000011101010111101",
			3733 => "0000000011101010111101",
			3734 => "0011000101100100110000",
			3735 => "0000011100011000001100",
			3736 => "0001110111010000001000",
			3737 => "0011101000101000000100",
			3738 => "0000001011101010111101",
			3739 => "0000000011101010111101",
			3740 => "0000000011101010111101",
			3741 => "0000011101011000010100",
			3742 => "0010000110001000010000",
			3743 => "0011111000110100001000",
			3744 => "0001111000011000000100",
			3745 => "0000000011101010111101",
			3746 => "0000000011101010111101",
			3747 => "0001110110110100000100",
			3748 => "0000000011101010111101",
			3749 => "0000000011101010111101",
			3750 => "0000000011101010111101",
			3751 => "0011111000011100000100",
			3752 => "0000000011101010111101",
			3753 => "0011101000000100000100",
			3754 => "0000000011101010111101",
			3755 => "0001101000010000000100",
			3756 => "0000000011101010111101",
			3757 => "0000000011101010111101",
			3758 => "0000000011101010111101",
			3759 => "0001011010111100001000",
			3760 => "0010000000101000000100",
			3761 => "1111111011101110110001",
			3762 => "0000000011101110110001",
			3763 => "0011000100000000010100",
			3764 => "0001000010111000001000",
			3765 => "0010010101011100000100",
			3766 => "0000000011101110110001",
			3767 => "0000000011101110110001",
			3768 => "0001011010111100000100",
			3769 => "0000000011101110110001",
			3770 => "0001101101011000000100",
			3771 => "0000000011101110110001",
			3772 => "0000001011101110110001",
			3773 => "0001000011000000101100",
			3774 => "0010110000011100010100",
			3775 => "0010101001000100010000",
			3776 => "0011000100011000001000",
			3777 => "0011100001111100000100",
			3778 => "0000000011101110110001",
			3779 => "0000000011101110110001",
			3780 => "0000000110001000000100",
			3781 => "0000000011101110110001",
			3782 => "0000000011101110110001",
			3783 => "0000000011101110110001",
			3784 => "0001010110100000001000",
			3785 => "0000011011111100000100",
			3786 => "0000000011101110110001",
			3787 => "0000001011101110110001",
			3788 => "0010100010101100001000",
			3789 => "0010010101010000000100",
			3790 => "0000000011101110110001",
			3791 => "0000000011101110110001",
			3792 => "0001001011101100000100",
			3793 => "0000000011101110110001",
			3794 => "0000000011101110110001",
			3795 => "0001100100111100011100",
			3796 => "0011001011000000010000",
			3797 => "0000000010011000001000",
			3798 => "0001001010110100000100",
			3799 => "1111111011101110110001",
			3800 => "0000000011101110110001",
			3801 => "0001111000111000000100",
			3802 => "0000000011101110110001",
			3803 => "0000000011101110110001",
			3804 => "0000011110010100000100",
			3805 => "0000000011101110110001",
			3806 => "0010000101000100000100",
			3807 => "0000000011101110110001",
			3808 => "0000000011101110110001",
			3809 => "0010111101111000001000",
			3810 => "0000011001111000000100",
			3811 => "0000000011101110110001",
			3812 => "0000001011101110110001",
			3813 => "0011000001011000001000",
			3814 => "0010011110010100000100",
			3815 => "0000000011101110110001",
			3816 => "0000000011101110110001",
			3817 => "0001011111100100000100",
			3818 => "1111111011101110110001",
			3819 => "0000000011101110110001",
			3820 => "0010110011011100001000",
			3821 => "0000100111011000000100",
			3822 => "1111111011110010111101",
			3823 => "0000000011110010111101",
			3824 => "0000000000111001000000",
			3825 => "0010001111001000110100",
			3826 => "0010101010110000100000",
			3827 => "0001001000001000010000",
			3828 => "0000010111101000001000",
			3829 => "0000010111101000000100",
			3830 => "0000000011110010111101",
			3831 => "1111111011110010111101",
			3832 => "0000001010101100000100",
			3833 => "0000000011110010111101",
			3834 => "0000000011110010111101",
			3835 => "0000101110100100001000",
			3836 => "0000001111000100000100",
			3837 => "0000000011110010111101",
			3838 => "1111111011110010111101",
			3839 => "0001001110111000000100",
			3840 => "0000000011110010111101",
			3841 => "0000000011110010111101",
			3842 => "0000000011111100001100",
			3843 => "0000011011101000000100",
			3844 => "0000000011110010111101",
			3845 => "0001010101110000000100",
			3846 => "0000001011110010111101",
			3847 => "0000000011110010111101",
			3848 => "0001101001111100000100",
			3849 => "0000001011110010111101",
			3850 => "0000000011110010111101",
			3851 => "0000011111001100000100",
			3852 => "1111111011110010111101",
			3853 => "0000010100110100000100",
			3854 => "0000000011110010111101",
			3855 => "0000000011110010111101",
			3856 => "0000101010110100110000",
			3857 => "0000000000110000010100",
			3858 => "0001001101001000001000",
			3859 => "0001101111000000000100",
			3860 => "1111111011110010111101",
			3861 => "0000000011110010111101",
			3862 => "0010011111001100000100",
			3863 => "0000000011110010111101",
			3864 => "0010101010110000000100",
			3865 => "0000000011110010111101",
			3866 => "0000001011110010111101",
			3867 => "0010101100011100001100",
			3868 => "0000100010000000001000",
			3869 => "0001000100001100000100",
			3870 => "0000000011110010111101",
			3871 => "0000000011110010111101",
			3872 => "1111111011110010111101",
			3873 => "0010000010101000001000",
			3874 => "0001101011001100000100",
			3875 => "0000000011110010111101",
			3876 => "0000001011110010111101",
			3877 => "0010100101000100000100",
			3878 => "0000000011110010111101",
			3879 => "0000000011110010111101",
			3880 => "0011100010100100001000",
			3881 => "0001100100101100000100",
			3882 => "0000000011110010111101",
			3883 => "1111111011110010111101",
			3884 => "0001100000001000000100",
			3885 => "0000001011110010111101",
			3886 => "0000000011110010111101",
			3887 => "0001001000000101000100",
			3888 => "0001001111100100011000",
			3889 => "0000111010000100010100",
			3890 => "0010100010101100010000",
			3891 => "0010110101100100001100",
			3892 => "0000011011111100000100",
			3893 => "0000000011111000101001",
			3894 => "0010110000011100000100",
			3895 => "0000000011111000101001",
			3896 => "0000000011111000101001",
			3897 => "0000000011111000101001",
			3898 => "0000000011111000101001",
			3899 => "0000000011111000101001",
			3900 => "0000111100111000011100",
			3901 => "0011001110001100010000",
			3902 => "0011001000111000001000",
			3903 => "0000110010001000000100",
			3904 => "0000000011111000101001",
			3905 => "0000000011111000101001",
			3906 => "0011001001110000000100",
			3907 => "0000000011111000101001",
			3908 => "0000000011111000101001",
			3909 => "0011001000000000001000",
			3910 => "0010010010101100000100",
			3911 => "0000000011111000101001",
			3912 => "0000000011111000101001",
			3913 => "0000000011111000101001",
			3914 => "0011001001001000001000",
			3915 => "0000100011000000000100",
			3916 => "0000000011111000101001",
			3917 => "0000000011111000101001",
			3918 => "0011000001101000000100",
			3919 => "0000000011111000101001",
			3920 => "0000000011111000101001",
			3921 => "0001001000110100001100",
			3922 => "0001101000010000001000",
			3923 => "0000000010011000000100",
			3924 => "1111111011111000101001",
			3925 => "0000000011111000101001",
			3926 => "0000000011111000101001",
			3927 => "0000101011110000111000",
			3928 => "0010111110001100011100",
			3929 => "0000110001011000010000",
			3930 => "0000011001111000001000",
			3931 => "0010110011011100000100",
			3932 => "0000000011111000101001",
			3933 => "0000000011111000101001",
			3934 => "0010111100110000000100",
			3935 => "0000000011111000101001",
			3936 => "0000000011111000101001",
			3937 => "0011111001011100000100",
			3938 => "0000001011111000101001",
			3939 => "0001101001100100000100",
			3940 => "0000000011111000101001",
			3941 => "0000000011111000101001",
			3942 => "0001001100001100001100",
			3943 => "0001100100111100000100",
			3944 => "0000000011111000101001",
			3945 => "0010101000010100000100",
			3946 => "0000000011111000101001",
			3947 => "0000000011111000101001",
			3948 => "0010101100011100001000",
			3949 => "0010010111101100000100",
			3950 => "1111111011111000101001",
			3951 => "0000000011111000101001",
			3952 => "0010111101010100000100",
			3953 => "0000000011111000101001",
			3954 => "0000000011111000101001",
			3955 => "0001100100101100011000",
			3956 => "0001000110001100001100",
			3957 => "0000111100001100001000",
			3958 => "0010111011110100000100",
			3959 => "0000000011111000101001",
			3960 => "0000000011111000101001",
			3961 => "0000000011111000101001",
			3962 => "0010100001110000001000",
			3963 => "0011100101010100000100",
			3964 => "0000000011111000101001",
			3965 => "0000000011111000101001",
			3966 => "0000000011111000101001",
			3967 => "0011100011010100010000",
			3968 => "0000101101001000001000",
			3969 => "0000010100110100000100",
			3970 => "0000000011111000101001",
			3971 => "0000000011111000101001",
			3972 => "0010000111000100000100",
			3973 => "0000000011111000101001",
			3974 => "1111111011111000101001",
			3975 => "0011011011101100000100",
			3976 => "0000000011111000101001",
			3977 => "0000000011111000101001",
			3978 => "0000001111000101011100",
			3979 => "0001111100101000010000",
			3980 => "0011001000111000001000",
			3981 => "0001101011001100000100",
			3982 => "0000000011111110111101",
			3983 => "0000000011111110111101",
			3984 => "0001111001110000000100",
			3985 => "0000000011111110111101",
			3986 => "0000000011111110111101",
			3987 => "0011011001011100100100",
			3988 => "0000000111000100010100",
			3989 => "0010100011101000001100",
			3990 => "0001010111100000001000",
			3991 => "0011001000000000000100",
			3992 => "0000000011111110111101",
			3993 => "0000000011111110111101",
			3994 => "0000000011111110111101",
			3995 => "0010000110011100000100",
			3996 => "0000000011111110111101",
			3997 => "0000000011111110111101",
			3998 => "0010011010100100001100",
			3999 => "0011001110001100000100",
			4000 => "0000000011111110111101",
			4001 => "0010100111110100000100",
			4002 => "0000000011111110111101",
			4003 => "0000000011111110111101",
			4004 => "0000000011111110111101",
			4005 => "0011001001001000001100",
			4006 => "0000001000101100001000",
			4007 => "0000111100111000000100",
			4008 => "0000000011111110111101",
			4009 => "1111111011111110111101",
			4010 => "0000000011111110111101",
			4011 => "0001101000010000001100",
			4012 => "0011011100010100000100",
			4013 => "0000000011111110111101",
			4014 => "0001010010000100000100",
			4015 => "0000000011111110111101",
			4016 => "0000000011111110111101",
			4017 => "0010001001101000001000",
			4018 => "0011011100010100000100",
			4019 => "0000000011111110111101",
			4020 => "0000000011111110111101",
			4021 => "0011101011110000000100",
			4022 => "0000000011111110111101",
			4023 => "0000000011111110111101",
			4024 => "0001011000000000101000",
			4025 => "0011011001001000100000",
			4026 => "0001111001110000010100",
			4027 => "0011111110010000010000",
			4028 => "0011011011000000001000",
			4029 => "0011001100001000000100",
			4030 => "0000000011111110111101",
			4031 => "0000000011111110111101",
			4032 => "0000111111011100000100",
			4033 => "0000000011111110111101",
			4034 => "0000000011111110111101",
			4035 => "0000000011111110111101",
			4036 => "0000110001011000001000",
			4037 => "0000100111010100000100",
			4038 => "0000000011111110111101",
			4039 => "0000000011111110111101",
			4040 => "0000000011111110111101",
			4041 => "0000110100000100000100",
			4042 => "0000000011111110111101",
			4043 => "0000001011111110111101",
			4044 => "0000101011110000100100",
			4045 => "0010100001010000001000",
			4046 => "0011100101100100000100",
			4047 => "0000000011111110111101",
			4048 => "1111111011111110111101",
			4049 => "0001110110000100010000",
			4050 => "0011000100000000001000",
			4051 => "0011010110100100000100",
			4052 => "0000000011111110111101",
			4053 => "0000000011111110111101",
			4054 => "0001101001100100000100",
			4055 => "0000000011111110111101",
			4056 => "0000000011111110111101",
			4057 => "0011101110110100001000",
			4058 => "0010111101111000000100",
			4059 => "0000000011111110111101",
			4060 => "1111111011111110111101",
			4061 => "0000000011111110111101",
			4062 => "0001100100101100011000",
			4063 => "0000101000001000001100",
			4064 => "0011001011000000000100",
			4065 => "0000000011111110111101",
			4066 => "0011101011110000000100",
			4067 => "0000000011111110111101",
			4068 => "0000000011111110111101",
			4069 => "0001110010001000001000",
			4070 => "0010000010101000000100",
			4071 => "0000000011111110111101",
			4072 => "0000000011111110111101",
			4073 => "0000000011111110111101",
			4074 => "0000101010110100000100",
			4075 => "0000000011111110111101",
			4076 => "0011101011100000000100",
			4077 => "1111111011111110111101",
			4078 => "0000000011111110111101",
			4079 => "0000110001101000111000",
			4080 => "0000111001110100101000",
			4081 => "0000111010111000011000",
			4082 => "0000110100001000000100",
			4083 => "1111111100000100111001",
			4084 => "0000100111011000001100",
			4085 => "0000100110010000000100",
			4086 => "1111111100000100111001",
			4087 => "0000100110010000000100",
			4088 => "0000000100000100111001",
			4089 => "1111111100000100111001",
			4090 => "0000100000010000000100",
			4091 => "0000001100000100111001",
			4092 => "1111111100000100111001",
			4093 => "0010100001110000001000",
			4094 => "0010111100101000000100",
			4095 => "1111111100000100111001",
			4096 => "0000001100000100111001",
			4097 => "0001111001110000000100",
			4098 => "0000010100000100111001",
			4099 => "1111111100000100111001",
			4100 => "0000000111111000000100",
			4101 => "1111111100000100111001",
			4102 => "0001111101100000001000",
			4103 => "0011111001010000000100",
			4104 => "0000011100000100111001",
			4105 => "1111111100000100111001",
			4106 => "1111111100000100111001",
			4107 => "0011000001101001101000",
			4108 => "0010101000100100110100",
			4109 => "0011110110111100011000",
			4110 => "0000111110101100001100",
			4111 => "0001110001111100000100",
			4112 => "1111111100000100111001",
			4113 => "0011110101110100000100",
			4114 => "1111111100000100111001",
			4115 => "0000101100000100111001",
			4116 => "0000010101011100000100",
			4117 => "1111111100000100111001",
			4118 => "0010001000100100000100",
			4119 => "0000010100000100111001",
			4120 => "1111111100000100111001",
			4121 => "0001010111100000010000",
			4122 => "0010011001111100001000",
			4123 => "0011000100011000000100",
			4124 => "0000010100000100111001",
			4125 => "0000100100000100111001",
			4126 => "0011010001000000000100",
			4127 => "1111111100000100111001",
			4128 => "0000001100000100111001",
			4129 => "0011011100010100000100",
			4130 => "1111111100000100111001",
			4131 => "0000010100110100000100",
			4132 => "0000011100000100111001",
			4133 => "1111111100000100111001",
			4134 => "0000110001011000011100",
			4135 => "0011001000111100010000",
			4136 => "0010101010110000001000",
			4137 => "0011011000000000000100",
			4138 => "1111111100000100111001",
			4139 => "0000000100000100111001",
			4140 => "0011011110110000000100",
			4141 => "1111111100000100111001",
			4142 => "0000010100000100111001",
			4143 => "0001111101100000001000",
			4144 => "0011111111010000000100",
			4145 => "0000010100000100111001",
			4146 => "1111111100000100111001",
			4147 => "1111111100000100111001",
			4148 => "0001010111111100010000",
			4149 => "0011100111010100001000",
			4150 => "0011001100110000000100",
			4151 => "0000010100000100111001",
			4152 => "0000000100000100111001",
			4153 => "0000001010101100000100",
			4154 => "0000001100000100111001",
			4155 => "0000010100000100111001",
			4156 => "0000000010111100000100",
			4157 => "1111111100000100111001",
			4158 => "0000010100000100111001",
			4159 => "0010011000010100011000",
			4160 => "0011011100010100000100",
			4161 => "0000001100000100111001",
			4162 => "0010110001001000001000",
			4163 => "0011001000011000000100",
			4164 => "0000010100000100111001",
			4165 => "1111111100000100111001",
			4166 => "0001011110010000000100",
			4167 => "0000000100000100111001",
			4168 => "0001110000011100000100",
			4169 => "0000000100000100111001",
			4170 => "1111111100000100111001",
			4171 => "0000000011010000000100",
			4172 => "1111111100000100111001",
			4173 => "0000010100000100111001",
			4174 => "0000010100110110001000",
			4175 => "0000100110111101000000",
			4176 => "0000110111110000100100",
			4177 => "0010100001010000001100",
			4178 => "0001010011100000000100",
			4179 => "0000000100001010011101",
			4180 => "0001001000101000000100",
			4181 => "0000000100001010011101",
			4182 => "1111111100001010011101",
			4183 => "0001111101100000001100",
			4184 => "0010010001000100001000",
			4185 => "0001111001110000000100",
			4186 => "0000000100001010011101",
			4187 => "0000000100001010011101",
			4188 => "0000000100001010011101",
			4189 => "0000110010001000001000",
			4190 => "0000010010001100000100",
			4191 => "0000000100001010011101",
			4192 => "0000000100001010011101",
			4193 => "0000000100001010011101",
			4194 => "0000111101000100001000",
			4195 => "0001100111101000000100",
			4196 => "0000000100001010011101",
			4197 => "0000001100001010011101",
			4198 => "0000100110111100010000",
			4199 => "0011001001001000001000",
			4200 => "0011001010111000000100",
			4201 => "0000000100001010011101",
			4202 => "0000000100001010011101",
			4203 => "0011001001110100000100",
			4204 => "0000000100001010011101",
			4205 => "0000000100001010011101",
			4206 => "0000000100001010011101",
			4207 => "0001101000010000110000",
			4208 => "0011001101010100011000",
			4209 => "0010101010110000001100",
			4210 => "0010010111101100001000",
			4211 => "0001000110111000000100",
			4212 => "0000000100001010011101",
			4213 => "1111111100001010011101",
			4214 => "0000000100001010011101",
			4215 => "0010000111000100000100",
			4216 => "0000001100001010011101",
			4217 => "0011111001011100000100",
			4218 => "0000000100001010011101",
			4219 => "0000000100001010011101",
			4220 => "0000011110010100001100",
			4221 => "0001101000010000001000",
			4222 => "0001101101011000000100",
			4223 => "0000000100001010011101",
			4224 => "0000000100001010011101",
			4225 => "0000000100001010011101",
			4226 => "0001111000011000001000",
			4227 => "0001110001101000000100",
			4228 => "0000000100001010011101",
			4229 => "0000000100001010011101",
			4230 => "1111111100001010011101",
			4231 => "0011000110000100001000",
			4232 => "0010101001101000000100",
			4233 => "0000000100001010011101",
			4234 => "0000000100001010011101",
			4235 => "0010000111000100001100",
			4236 => "0001111111011100000100",
			4237 => "0000000100001010011101",
			4238 => "0000100010110000000100",
			4239 => "1111111100001010011101",
			4240 => "0000000100001010011101",
			4241 => "1111111100001010011101",
			4242 => "0011000101100100101000",
			4243 => "0000011100011000001000",
			4244 => "0001110111010000000100",
			4245 => "0000000100001010011101",
			4246 => "0000000100001010011101",
			4247 => "0000011101011000011000",
			4248 => "0000111100001100010000",
			4249 => "0011111000110100001000",
			4250 => "0001111000011000000100",
			4251 => "0000000100001010011101",
			4252 => "0000000100001010011101",
			4253 => "0001110110110100000100",
			4254 => "0000000100001010011101",
			4255 => "0000000100001010011101",
			4256 => "0000011010011000000100",
			4257 => "0000000100001010011101",
			4258 => "0000000100001010011101",
			4259 => "0000111100001100000100",
			4260 => "0000000100001010011101",
			4261 => "0000000100001010011101",
			4262 => "0000000100001010011101",
			4263 => "0001001100001101001100",
			4264 => "0000000010111101000100",
			4265 => "0011000100011000011100",
			4266 => "0010101010110000011000",
			4267 => "0000001111000100010000",
			4268 => "0001000010010100001000",
			4269 => "0000000110001000000100",
			4270 => "0000000100001111101001",
			4271 => "0000000100001111101001",
			4272 => "0010010111101100000100",
			4273 => "0000000100001111101001",
			4274 => "0000000100001111101001",
			4275 => "0000110001011000000100",
			4276 => "0000000100001111101001",
			4277 => "0000000100001111101001",
			4278 => "1111111100001111101001",
			4279 => "0011000001101000010100",
			4280 => "0000011001011000000100",
			4281 => "0000000100001111101001",
			4282 => "0010011010100100001000",
			4283 => "0000100110111000000100",
			4284 => "0000000100001111101001",
			4285 => "0000000100001111101001",
			4286 => "0001001110000000000100",
			4287 => "0000000100001111101001",
			4288 => "0000000100001111101001",
			4289 => "0011111000110100001000",
			4290 => "0001010110010000000100",
			4291 => "0000000100001111101001",
			4292 => "0000000100001111101001",
			4293 => "0010000001010100000100",
			4294 => "0000000100001111101001",
			4295 => "0000001010101100000100",
			4296 => "0000000100001111101001",
			4297 => "0000000100001111101001",
			4298 => "0000110000011100000100",
			4299 => "0000000100001111101001",
			4300 => "0000001100001111101001",
			4301 => "0001000110001100010000",
			4302 => "0010101000010100000100",
			4303 => "0000000100001111101001",
			4304 => "0011001000111100000100",
			4305 => "0000000100001111101001",
			4306 => "0001001100001100000100",
			4307 => "0000000100001111101001",
			4308 => "1111111100001111101001",
			4309 => "0000001111000100010100",
			4310 => "0000110000010000000100",
			4311 => "0000000100001111101001",
			4312 => "0010010011101000001100",
			4313 => "0010101010110000001000",
			4314 => "0010000001010100000100",
			4315 => "0000000100001111101001",
			4316 => "0000000100001111101001",
			4317 => "0000000100001111101001",
			4318 => "0000000100001111101001",
			4319 => "0010101010110000011000",
			4320 => "0000101110100100001100",
			4321 => "0011100110111000001000",
			4322 => "0000001111000100000100",
			4323 => "0000000100001111101001",
			4324 => "1111111100001111101001",
			4325 => "0000000100001111101001",
			4326 => "0000011100011000001000",
			4327 => "0011101000001000000100",
			4328 => "0000000100001111101001",
			4329 => "0000000100001111101001",
			4330 => "0000000100001111101001",
			4331 => "0000101111010100010000",
			4332 => "0000111011011100001000",
			4333 => "0000101100010000000100",
			4334 => "0000000100001111101001",
			4335 => "0000000100001111101001",
			4336 => "0010101100011100000100",
			4337 => "0000001100001111101001",
			4338 => "0000000100001111101001",
			4339 => "0000000000111000001000",
			4340 => "0011100010000100000100",
			4341 => "0000000100001111101001",
			4342 => "0000000100001111101001",
			4343 => "0000000111111000000100",
			4344 => "0000000100001111101001",
			4345 => "0000000100001111101001",
			4346 => "0000111001110100010100",
			4347 => "0000010111100100010000",
			4348 => "0000110100001000000100",
			4349 => "1111111100010100011101",
			4350 => "0010001000110000000100",
			4351 => "1111111100010100011101",
			4352 => "0001111001110000000100",
			4353 => "0000010100010100011101",
			4354 => "1111111100010100011101",
			4355 => "0000001100010100011101",
			4356 => "0011000001101001100100",
			4357 => "0010000101000100101000",
			4358 => "0000001100000100001100",
			4359 => "0000010001000100001000",
			4360 => "0010001000010100000100",
			4361 => "1111111100010100011101",
			4362 => "0000000100010100011101",
			4363 => "0000010100010100011101",
			4364 => "0001001000001100001100",
			4365 => "0011011111010000001000",
			4366 => "0011000100001000000100",
			4367 => "1111111100010100011101",
			4368 => "0000011100010100011101",
			4369 => "1111111100010100011101",
			4370 => "0000111100010000001000",
			4371 => "0011000100011000000100",
			4372 => "1111111100010100011101",
			4373 => "0000000100010100011101",
			4374 => "0000000001110100000100",
			4375 => "0000000100010100011101",
			4376 => "0000011100010100011101",
			4377 => "0000110001011000100000",
			4378 => "0001001001001100010000",
			4379 => "0000110100000100001000",
			4380 => "0000111010001100000100",
			4381 => "1111111100010100011101",
			4382 => "0000000100010100011101",
			4383 => "0000101110110100000100",
			4384 => "0000010100010100011101",
			4385 => "1111111100010100011101",
			4386 => "0011111001010000001000",
			4387 => "0001111101100000000100",
			4388 => "0000010100010100011101",
			4389 => "1111111100010100011101",
			4390 => "0000110000011100000100",
			4391 => "1111111100010100011101",
			4392 => "0000001100010100011101",
			4393 => "0001000100001100010000",
			4394 => "0010000001110000001000",
			4395 => "0001001110000000000100",
			4396 => "0000010100010100011101",
			4397 => "0000000100010100011101",
			4398 => "0001110111010000000100",
			4399 => "0000010100010100011101",
			4400 => "1111111100010100011101",
			4401 => "0011001000111000000100",
			4402 => "0000010100010100011101",
			4403 => "0011111000001100000100",
			4404 => "1111111100010100011101",
			4405 => "0000001100010100011101",
			4406 => "0010011000010100011100",
			4407 => "0001010111111100001000",
			4408 => "0011101011111000000100",
			4409 => "1111111100010100011101",
			4410 => "0000010100010100011101",
			4411 => "0010000110001000010000",
			4412 => "0001000011110100001000",
			4413 => "0000010001000100000100",
			4414 => "0000110100010100011101",
			4415 => "1111111100010100011101",
			4416 => "0010000110001000000100",
			4417 => "0010001100010100011101",
			4418 => "0000011100010100011101",
			4419 => "1111111100010100011101",
			4420 => "0000110100001100000100",
			4421 => "1111111100010100011101",
			4422 => "0000011100010100011101",
			4423 => "0010110011011100001100",
			4424 => "0010101111001000000100",
			4425 => "1111111100011000001001",
			4426 => "0000000111010000000100",
			4427 => "0000001100011000001001",
			4428 => "0000000100011000001001",
			4429 => "0010101001101001100100",
			4430 => "0010001010110000101000",
			4431 => "0001001111100100010100",
			4432 => "0000111010000100010000",
			4433 => "0011110110111100001000",
			4434 => "0001010110100000000100",
			4435 => "0000000100011000001001",
			4436 => "0000000100011000001001",
			4437 => "0010111011011100000100",
			4438 => "0000001100011000001001",
			4439 => "0000000100011000001001",
			4440 => "1111111100011000001001",
			4441 => "0011001001110100010000",
			4442 => "0011000100011000001000",
			4443 => "0011001010111000000100",
			4444 => "0000000100011000001001",
			4445 => "0000000100011000001001",
			4446 => "0011001011000000000100",
			4447 => "0000010100011000001001",
			4448 => "0000001100011000001001",
			4449 => "0000000100011000001001",
			4450 => "0001000010100100100000",
			4451 => "0000110000011100010000",
			4452 => "0001000010111000001000",
			4453 => "0011111111010000000100",
			4454 => "1111111100011000001001",
			4455 => "1111110100011000001001",
			4456 => "0011000000101000000100",
			4457 => "0000001100011000001001",
			4458 => "0000000100011000001001",
			4459 => "0011110010011100001000",
			4460 => "0001111101100000000100",
			4461 => "0000001100011000001001",
			4462 => "0000000100011000001001",
			4463 => "0000110101110100000100",
			4464 => "0000000100011000001001",
			4465 => "0000000100011000001001",
			4466 => "0010110110000100001100",
			4467 => "0001011010111100000100",
			4468 => "0000000100011000001001",
			4469 => "0011001000111000000100",
			4470 => "0000001100011000001001",
			4471 => "0000000100011000001001",
			4472 => "0000111010001100001000",
			4473 => "0000111010011100000100",
			4474 => "1111111100011000001001",
			4475 => "0000000100011000001001",
			4476 => "0001001011100000000100",
			4477 => "0000001100011000001001",
			4478 => "0000000100011000001001",
			4479 => "0011001000111100000100",
			4480 => "0000001100011000001001",
			4481 => "1111111100011000001001",
			4482 => "0001101011001101100000",
			4483 => "0010011000010000111000",
			4484 => "0001101101011000011100",
			4485 => "0000010110101000000100",
			4486 => "1111111100011110010101",
			4487 => "0000000001110000001100",
			4488 => "0011010100010000001000",
			4489 => "0010110100011000000100",
			4490 => "1111111100011110010101",
			4491 => "0000010100011110010101",
			4492 => "1111111100011110010101",
			4493 => "0011110010000100001000",
			4494 => "0001111100101000000100",
			4495 => "1111111100011110010101",
			4496 => "0000011100011110010101",
			4497 => "1111111100011110010101",
			4498 => "0000111001110100000100",
			4499 => "1111111100011110010101",
			4500 => "0011110001000000001100",
			4501 => "0011001000111100001000",
			4502 => "0000110001101000000100",
			4503 => "0000001100011110010101",
			4504 => "0000011100011110010101",
			4505 => "0000000100011110010101",
			4506 => "0010011111000000001000",
			4507 => "0000101110110100000100",
			4508 => "0000000100011110010101",
			4509 => "1111111100011110010101",
			4510 => "0000010100011110010101",
			4511 => "0000101000001100011000",
			4512 => "0010101010100000000100",
			4513 => "0000010100011110010101",
			4514 => "0011000100011000010000",
			4515 => "0000111100000000001000",
			4516 => "0000101110110100000100",
			4517 => "0000000100011110010101",
			4518 => "1111111100011110010101",
			4519 => "0011010101001000000100",
			4520 => "0000011100011110010101",
			4521 => "0000000100011110010101",
			4522 => "1111111100011110010101",
			4523 => "0001101011001100001100",
			4524 => "0011001011000000000100",
			4525 => "0000011100011110010101",
			4526 => "0001101101011000000100",
			4527 => "1111111100011110010101",
			4528 => "0000001100011110010101",
			4529 => "1111111100011110010101",
			4530 => "0011000001101001000100",
			4531 => "0010101000010100011100",
			4532 => "0000011011111100000100",
			4533 => "0000010100011110010101",
			4534 => "0011101100010000001000",
			4535 => "0010100011101000000100",
			4536 => "0000001100011110010101",
			4537 => "1111111100011110010101",
			4538 => "0010110110110100001000",
			4539 => "0000010111101000000100",
			4540 => "0000100100011110010101",
			4541 => "0000001100011110010101",
			4542 => "0011011100010100000100",
			4543 => "1111111100011110010101",
			4544 => "0000001100011110010101",
			4545 => "0000001100101100100000",
			4546 => "0001101001100100010000",
			4547 => "0001110101101100001000",
			4548 => "0001011101010100000100",
			4549 => "1111111100011110010101",
			4550 => "0000001100011110010101",
			4551 => "0000100011000000000100",
			4552 => "1111111100011110010101",
			4553 => "0000000100011110010101",
			4554 => "0001110111010000001000",
			4555 => "0000001010101100000100",
			4556 => "0000000100011110010101",
			4557 => "0000001100011110010101",
			4558 => "0000110110001100000100",
			4559 => "1111111100011110010101",
			4560 => "0000001100011110010101",
			4561 => "0001101111000000000100",
			4562 => "1111111100011110010101",
			4563 => "0000000100011110010101",
			4564 => "0010011000010100011100",
			4565 => "0001010111111100001000",
			4566 => "0011111011110000000100",
			4567 => "1111111100011110010101",
			4568 => "0000001100011110010101",
			4569 => "0001101111000000000100",
			4570 => "0000001100011110010101",
			4571 => "0011010110111100001000",
			4572 => "0001110001011000000100",
			4573 => "0000000100011110010101",
			4574 => "1111111100011110010101",
			4575 => "0010101010110000000100",
			4576 => "0000000100011110010101",
			4577 => "1111111100011110010101",
			4578 => "0000110100001100000100",
			4579 => "1111111100011110010101",
			4580 => "0000010100011110010101",
			4581 => "0010010001111001010100",
			4582 => "0010111100101100101000",
			4583 => "0001101101011000000100",
			4584 => "1111111100100011010001",
			4585 => "0011001001110000100000",
			4586 => "0000101100000000010000",
			4587 => "0000110100000100001000",
			4588 => "0001000100001100000100",
			4589 => "0000000100100011010001",
			4590 => "0000000100100011010001",
			4591 => "0011100101110100000100",
			4592 => "0000001100100011010001",
			4593 => "0000000100100011010001",
			4594 => "0000100111011000001000",
			4595 => "0001111000111000000100",
			4596 => "0000000100100011010001",
			4597 => "1111111100100011010001",
			4598 => "0011011011000000000100",
			4599 => "0000000100100011010001",
			4600 => "0000000100100011010001",
			4601 => "1111111100100011010001",
			4602 => "0001101000010000100100",
			4603 => "0001000110001100011000",
			4604 => "0011001000111100001000",
			4605 => "0001101011001100000100",
			4606 => "0000000100100011010001",
			4607 => "0000000100100011010001",
			4608 => "0011000110000100001000",
			4609 => "0001011001001000000100",
			4610 => "0000000100100011010001",
			4611 => "1111111100100011010001",
			4612 => "0001100001000100000100",
			4613 => "0000000100100011010001",
			4614 => "0000000100100011010001",
			4615 => "0001010100011000000100",
			4616 => "0000000100100011010001",
			4617 => "0000110000110100000100",
			4618 => "1111111100100011010001",
			4619 => "0000000100100011010001",
			4620 => "0010011110010100000100",
			4621 => "0000000100100011010001",
			4622 => "0000000100100011010001",
			4623 => "0001011010011100000100",
			4624 => "0000001100100011010001",
			4625 => "0000110010000000010100",
			4626 => "0000000000111000001000",
			4627 => "0000101100010000000100",
			4628 => "0000000100100011010001",
			4629 => "1111111100100011010001",
			4630 => "0001001100111100001000",
			4631 => "0001111100101000000100",
			4632 => "0000001100100011010001",
			4633 => "0000000100100011010001",
			4634 => "0000000100100011010001",
			4635 => "0011011111010000100000",
			4636 => "0011000100011000010000",
			4637 => "0011111111010100001000",
			4638 => "0010000110011000000100",
			4639 => "0000000100100011010001",
			4640 => "0000000100100011010001",
			4641 => "0011111011110000000100",
			4642 => "0000001100100011010001",
			4643 => "0000000100100011010001",
			4644 => "0011000100011000001000",
			4645 => "0001011101000100000100",
			4646 => "1111111100100011010001",
			4647 => "0000000100100011010001",
			4648 => "0011001000000000000100",
			4649 => "0000000100100011010001",
			4650 => "0000000100100011010001",
			4651 => "0011000111001000000100",
			4652 => "1111111100100011010001",
			4653 => "0001101101011000001000",
			4654 => "0010011000010000000100",
			4655 => "0000000100100011010001",
			4656 => "0000000100100011010001",
			4657 => "0000111101101100000100",
			4658 => "0000000100100011010001",
			4659 => "0000000100100011010001",
			4660 => "0011101110101101100000",
			4661 => "0010111100101100111000",
			4662 => "0001001000000100001100",
			4663 => "0011000100000000000100",
			4664 => "0000000100101010101101",
			4665 => "0011011001110100000100",
			4666 => "1111111100101010101101",
			4667 => "0000000100101010101101",
			4668 => "0000110100000100011100",
			4669 => "0001001111100000010000",
			4670 => "0010110101101100001000",
			4671 => "0001101011001100000100",
			4672 => "0000000100101010101101",
			4673 => "0000000100101010101101",
			4674 => "0001111000111100000100",
			4675 => "0000000100101010101101",
			4676 => "1111111100101010101101",
			4677 => "0001010100001000000100",
			4678 => "0000000100101010101101",
			4679 => "0001111101100000000100",
			4680 => "0000000100101010101101",
			4681 => "0000000100101010101101",
			4682 => "0011111110010000001000",
			4683 => "0011011011000000000100",
			4684 => "0000000100101010101101",
			4685 => "0000001100101010101101",
			4686 => "0011010110100100000100",
			4687 => "1111111100101010101101",
			4688 => "0000000100101010101101",
			4689 => "0000100110010000010100",
			4690 => "0001001011110000001100",
			4691 => "0011110010110100000100",
			4692 => "0000000100101010101101",
			4693 => "0000001000101100000100",
			4694 => "0000000100101010101101",
			4695 => "0000000100101010101101",
			4696 => "0000000010111100000100",
			4697 => "0000000100101010101101",
			4698 => "0000000100101010101101",
			4699 => "0001101000010000001100",
			4700 => "0011000100000000000100",
			4701 => "0000000100101010101101",
			4702 => "0010010111101000000100",
			4703 => "1111111100101010101101",
			4704 => "0000000100101010101101",
			4705 => "0001011001110100000100",
			4706 => "0000000100101010101101",
			4707 => "0000000100101010101101",
			4708 => "0001010111100000111100",
			4709 => "0001100100111100101100",
			4710 => "0011000100001000010000",
			4711 => "0001000000010100001100",
			4712 => "0010110000001100000100",
			4713 => "0000000100101010101101",
			4714 => "0001110111001000000100",
			4715 => "1111111100101010101101",
			4716 => "0000000100101010101101",
			4717 => "0000000100101010101101",
			4718 => "0010010100101100001100",
			4719 => "0011010101110000001000",
			4720 => "0000001100000100000100",
			4721 => "0000000100101010101101",
			4722 => "0000000100101010101101",
			4723 => "0000000100101010101101",
			4724 => "0001001011101100001000",
			4725 => "0010110000011100000100",
			4726 => "0000000100101010101101",
			4727 => "0000000100101010101101",
			4728 => "0001001011110000000100",
			4729 => "0000000100101010101101",
			4730 => "0000000100101010101101",
			4731 => "0000000011010000001000",
			4732 => "0010011101111100000100",
			4733 => "0000000100101010101101",
			4734 => "0000001100101010101101",
			4735 => "0011000110000100000100",
			4736 => "0000000100101010101101",
			4737 => "0000000100101010101101",
			4738 => "0001010010011100100000",
			4739 => "0001111000011000010000",
			4740 => "0010000001010100001000",
			4741 => "0011001001110100000100",
			4742 => "0000000100101010101101",
			4743 => "0000000100101010101101",
			4744 => "0001001001001100000100",
			4745 => "0000000100101010101101",
			4746 => "0000000100101010101101",
			4747 => "0000110010010100001100",
			4748 => "0010110110110100000100",
			4749 => "0000000100101010101101",
			4750 => "0011010111111100000100",
			4751 => "0000000100101010101101",
			4752 => "1111111100101010101101",
			4753 => "0000000100101010101101",
			4754 => "0011101000101000010100",
			4755 => "0011010011001000000100",
			4756 => "0000000100101010101101",
			4757 => "0011000001101000001000",
			4758 => "0000001011010100000100",
			4759 => "0000000100101010101101",
			4760 => "0000001100101010101101",
			4761 => "0000110010010100000100",
			4762 => "0000000100101010101101",
			4763 => "0000000100101010101101",
			4764 => "0001010011001000010000",
			4765 => "0011101011110000001000",
			4766 => "0000110010010100000100",
			4767 => "0000000100101010101101",
			4768 => "1111111100101010101101",
			4769 => "0001011110010000000100",
			4770 => "0000000100101010101101",
			4771 => "0000000100101010101101",
			4772 => "0001110110110100001000",
			4773 => "0011011100000000000100",
			4774 => "0000000100101010101101",
			4775 => "0000000100101010101101",
			4776 => "0010011010100000000100",
			4777 => "0000000100101010101101",
			4778 => "0000000100101010101101",
			4779 => "0001010100001000001100",
			4780 => "0000001000011000000100",
			4781 => "1111111100101111111001",
			4782 => "0001000100100100000100",
			4783 => "0000000100101111111001",
			4784 => "0000000100101111111001",
			4785 => "0011110010011101001000",
			4786 => "0001101101011000010100",
			4787 => "0011101011011100001000",
			4788 => "0001101001011000000100",
			4789 => "0000000100101111111001",
			4790 => "1111111100101111111001",
			4791 => "0000011101101000000100",
			4792 => "0000000100101111111001",
			4793 => "0010000010101100000100",
			4794 => "0000000100101111111001",
			4795 => "0000001100101111111001",
			4796 => "0000101100010000011100",
			4797 => "0001001001001100010000",
			4798 => "0010110101101100001000",
			4799 => "0010100001010000000100",
			4800 => "0000000100101111111001",
			4801 => "1111111100101111111001",
			4802 => "0000000000110000000100",
			4803 => "0000000100101111111001",
			4804 => "0000000100101111111001",
			4805 => "0011001000111000001000",
			4806 => "0010110011011100000100",
			4807 => "0000000100101111111001",
			4808 => "0000001100101111111001",
			4809 => "0000000100101111111001",
			4810 => "0001101111000000010000",
			4811 => "0000010010001100001000",
			4812 => "0000100111011000000100",
			4813 => "0000000100101111111001",
			4814 => "0000000100101111111001",
			4815 => "0010011101011100000100",
			4816 => "1111111100101111111001",
			4817 => "0000000100101111111001",
			4818 => "0011001000111000000100",
			4819 => "0000001100101111111001",
			4820 => "0000000100101111111001",
			4821 => "0001001110100100101000",
			4822 => "0001101000010000011000",
			4823 => "0000010111100100001000",
			4824 => "0001001000110100000100",
			4825 => "1111111100101111111001",
			4826 => "0000000100101111111001",
			4827 => "0001010001101000001000",
			4828 => "0000001000110000000100",
			4829 => "0000000100101111111001",
			4830 => "0000001100101111111001",
			4831 => "0011000100001000000100",
			4832 => "1111111100101111111001",
			4833 => "0000000100101111111001",
			4834 => "0000000001110100000100",
			4835 => "0000000100101111111001",
			4836 => "0011001111011100001000",
			4837 => "0000011101011000000100",
			4838 => "0000001100101111111001",
			4839 => "0000000100101111111001",
			4840 => "0000000100101111111001",
			4841 => "0001101000010000011000",
			4842 => "0010111100101100001100",
			4843 => "0011011001001000001000",
			4844 => "0001000010111000000100",
			4845 => "1111111100101111111001",
			4846 => "0000000100101111111001",
			4847 => "0000001100101111111001",
			4848 => "0011001000111000000100",
			4849 => "1111111100101111111001",
			4850 => "0000011011111100000100",
			4851 => "0000000100101111111001",
			4852 => "1111111100101111111001",
			4853 => "0010111010111100000100",
			4854 => "0000001100101111111001",
			4855 => "0000101011110000001000",
			4856 => "0001101000010000000100",
			4857 => "1111111100101111111001",
			4858 => "0000000100101111111001",
			4859 => "0000001111000100000100",
			4860 => "0000000100101111111001",
			4861 => "0000000100101111111001",
			4862 => "0000111011000000001100",
			4863 => "0001101001100100000100",
			4864 => "1111111100110100111101",
			4865 => "0001111000111000000100",
			4866 => "0000001100110100111101",
			4867 => "1111111100110100111101",
			4868 => "0001100100111101001100",
			4869 => "0001110101101100100100",
			4870 => "0001101101011000000100",
			4871 => "1111111100110100111101",
			4872 => "0000100010000100010000",
			4873 => "0000110100000100001000",
			4874 => "0001001111100000000100",
			4875 => "0000000100110100111101",
			4876 => "0000001100110100111101",
			4877 => "0000101100010100000100",
			4878 => "0000000100110100111101",
			4879 => "0000001100110100111101",
			4880 => "0001101001100100001000",
			4881 => "0010011011101000000100",
			4882 => "0000001100110100111101",
			4883 => "1111111100110100111101",
			4884 => "0011110111111100000100",
			4885 => "0000001100110100111101",
			4886 => "0000000100110100111101",
			4887 => "0010101001000100011100",
			4888 => "0010110110110100010000",
			4889 => "0011101100010000001000",
			4890 => "0010001010110000000100",
			4891 => "0000000100110100111101",
			4892 => "0000000100110100111101",
			4893 => "0010100010101100000100",
			4894 => "0000010100110100111101",
			4895 => "0000000100110100111101",
			4896 => "0010010100101100001000",
			4897 => "0011111011101100000100",
			4898 => "1111111100110100111101",
			4899 => "0000001100110100111101",
			4900 => "1111111100110100111101",
			4901 => "0010101001000100000100",
			4902 => "1111110100110100111101",
			4903 => "0010101001000100000100",
			4904 => "0000001100110100111101",
			4905 => "1111111100110100111101",
			4906 => "0001010001000000011100",
			4907 => "0001000111011100010000",
			4908 => "0011100011001000001000",
			4909 => "0001110110000100000100",
			4910 => "0000001100110100111101",
			4911 => "0000000100110100111101",
			4912 => "0010000001010100000100",
			4913 => "0000000100110100111101",
			4914 => "0000001100110100111101",
			4915 => "0010010001000100000100",
			4916 => "0000001100110100111101",
			4917 => "0001001100111100000100",
			4918 => "0000000100110100111101",
			4919 => "1111111100110100111101",
			4920 => "0011111000000100010100",
			4921 => "0001111000011000000100",
			4922 => "0000000100110100111101",
			4923 => "0010000101000100001000",
			4924 => "0001101000010000000100",
			4925 => "0000000100110100111101",
			4926 => "0000001100110100111101",
			4927 => "0011111110000000000100",
			4928 => "1111111100110100111101",
			4929 => "0000000100110100111101",
			4930 => "0000110110001100010000",
			4931 => "0010000001010100001000",
			4932 => "0000110101000000000100",
			4933 => "0000000100110100111101",
			4934 => "0000011100110100111101",
			4935 => "0000000000110000000100",
			4936 => "0000001100110100111101",
			4937 => "1111111100110100111101",
			4938 => "0000001011000100001000",
			4939 => "0011100010110000000100",
			4940 => "1111111100110100111101",
			4941 => "0000000100110100111101",
			4942 => "1111111100110100111101",
			4943 => "0001101101011000110100",
			4944 => "0000000110001000100100",
			4945 => "0000000101000100000100",
			4946 => "1111111100111011011001",
			4947 => "0010110101100100010000",
			4948 => "0011001011000000001100",
			4949 => "0011001110001100000100",
			4950 => "1111111100111011011001",
			4951 => "0011011110101100000100",
			4952 => "0000010100111011011001",
			4953 => "0000000100111011011001",
			4954 => "0000011100111011011001",
			4955 => "0000101000001100001000",
			4956 => "0011011111010000000100",
			4957 => "0000000100111011011001",
			4958 => "1111111100111011011001",
			4959 => "0010111011110100000100",
			4960 => "0000010100111011011001",
			4961 => "1111111100111011011001",
			4962 => "0000111010001100000100",
			4963 => "1111111100111011011001",
			4964 => "0011111111010000001000",
			4965 => "0011110111100000000100",
			4966 => "1111111100111011011001",
			4967 => "0000001100111011011001",
			4968 => "1111111100111011011001",
			4969 => "0011001000011001110100",
			4970 => "0001101111000001000000",
			4971 => "0000101100000000100000",
			4972 => "0010111100101100010000",
			4973 => "0000110001101000001000",
			4974 => "0001001111100000000100",
			4975 => "1111111100111011011001",
			4976 => "0000001100111011011001",
			4977 => "0011010100011000000100",
			4978 => "0000000100111011011001",
			4979 => "0000001100111011011001",
			4980 => "0001000010010100001000",
			4981 => "0001101001100100000100",
			4982 => "1111111100111011011001",
			4983 => "0000001100111011011001",
			4984 => "0000000010011000000100",
			4985 => "1111110100111011011001",
			4986 => "0000000100111011011001",
			4987 => "0000111100010000010000",
			4988 => "0011001000111100001000",
			4989 => "0000101010000100000100",
			4990 => "0000000100111011011001",
			4991 => "1111111100111011011001",
			4992 => "0011110110100000000100",
			4993 => "0000000100111011011001",
			4994 => "1111111100111011011001",
			4995 => "0011111010000100001000",
			4996 => "0011100010000100000100",
			4997 => "0000000100111011011001",
			4998 => "0000010100111011011001",
			4999 => "0000001011010100000100",
			5000 => "1111111100111011011001",
			5001 => "0000000100111011011001",
			5002 => "0010000001110000011000",
			5003 => "0001111000011000001100",
			5004 => "0001001000011100001000",
			5005 => "0000000111000100000100",
			5006 => "1111111100111011011001",
			5007 => "0000001100111011011001",
			5008 => "0000000100111011011001",
			5009 => "0001010001000000000100",
			5010 => "0000001100111011011001",
			5011 => "0010111010010100000100",
			5012 => "1111111100111011011001",
			5013 => "0000000100111011011001",
			5014 => "0011100001011100010000",
			5015 => "0001110110000100001000",
			5016 => "0011011011000000000100",
			5017 => "0000000100111011011001",
			5018 => "0000001100111011011001",
			5019 => "0000111110010000000100",
			5020 => "0000000100111011011001",
			5021 => "0000001100111011011001",
			5022 => "0001101000010000000100",
			5023 => "0000010100111011011001",
			5024 => "0010111011110100000100",
			5025 => "0000001100111011011001",
			5026 => "0000000100111011011001",
			5027 => "0011010110111100010000",
			5028 => "0011000001011000001000",
			5029 => "0001101111000000000100",
			5030 => "0000000100111011011001",
			5031 => "1111111100111011011001",
			5032 => "0000111000110100000100",
			5033 => "0000010100111011011001",
			5034 => "0000000100111011011001",
			5035 => "0000000111000000001000",
			5036 => "0011101110000000000100",
			5037 => "0000000100111011011001",
			5038 => "0001001100111011011001",
			5039 => "0000001011000100001100",
			5040 => "0001001010110100000100",
			5041 => "1111111100111011011001",
			5042 => "0010100001010000000100",
			5043 => "0000010100111011011001",
			5044 => "0000000100111011011001",
			5045 => "1111111100111011011001",
			5046 => "0001101101011000111100",
			5047 => "0010010101010000100000",
			5048 => "0000010111100100001100",
			5049 => "0000111010001100000100",
			5050 => "1111111101000001110101",
			5051 => "0000110100000100000100",
			5052 => "0000000101000001110101",
			5053 => "1111111101000001110101",
			5054 => "0001110011100000010000",
			5055 => "0011001110001100000100",
			5056 => "1111111101000001110101",
			5057 => "0000000001110000000100",
			5058 => "1111111101000001110101",
			5059 => "0000001101010000000100",
			5060 => "0000010101000001110101",
			5061 => "0000000101000001110101",
			5062 => "1111111101000001110101",
			5063 => "0010101010100100001000",
			5064 => "0010110101100100000100",
			5065 => "0000010101000001110101",
			5066 => "0000000101000001110101",
			5067 => "0010110000011100000100",
			5068 => "1111111101000001110101",
			5069 => "0000011110010100001100",
			5070 => "0001110110100100000100",
			5071 => "0000001101000001110101",
			5072 => "0000010001000100000100",
			5073 => "0000000101000001110101",
			5074 => "1111111101000001110101",
			5075 => "0000001101000001110101",
			5076 => "0010110000110101101000",
			5077 => "0001101111000000111000",
			5078 => "0010111100101100011000",
			5079 => "0011111110010000010000",
			5080 => "0000110001011000001000",
			5081 => "0011111001010000000100",
			5082 => "0000001101000001110101",
			5083 => "1111111101000001110101",
			5084 => "0001001000000100000100",
			5085 => "0000001101000001110101",
			5086 => "0000001101000001110101",
			5087 => "0000110111110000000100",
			5088 => "1111111101000001110101",
			5089 => "0000000101000001110101",
			5090 => "0001000110111000010000",
			5091 => "0010101000100100001000",
			5092 => "0011111010000100000100",
			5093 => "0000001101000001110101",
			5094 => "0000000101000001110101",
			5095 => "0000011101101000000100",
			5096 => "0000001101000001110101",
			5097 => "0000010101000001110101",
			5098 => "0010111010001100001000",
			5099 => "0000001111000100000100",
			5100 => "1111111101000001110101",
			5101 => "0000000101000001110101",
			5102 => "0000010111101000000100",
			5103 => "0000001101000001110101",
			5104 => "1111111101000001110101",
			5105 => "0011100110111000100000",
			5106 => "0001010001000000010000",
			5107 => "0011101111100100001000",
			5108 => "0001110110000100000100",
			5109 => "0000001101000001110101",
			5110 => "0000000101000001110101",
			5111 => "0010010010101100000100",
			5112 => "0000001101000001110101",
			5113 => "0000000101000001110101",
			5114 => "0001111000011000001000",
			5115 => "0001001011110000000100",
			5116 => "0000000101000001110101",
			5117 => "0000001101000001110101",
			5118 => "0000111111101000000100",
			5119 => "1111111101000001110101",
			5120 => "0000000101000001110101",
			5121 => "0001101000010000000100",
			5122 => "0000100101000001110101",
			5123 => "0001010011001000001000",
			5124 => "0011001001110100000100",
			5125 => "0000001101000001110101",
			5126 => "0000000101000001110101",
			5127 => "1111111101000001110101",
			5128 => "0000001011000100101000",
			5129 => "0010011010100000010100",
			5130 => "0001101001111100001100",
			5131 => "0010010000001000001000",
			5132 => "0001010110010000000100",
			5133 => "0000000101000001110101",
			5134 => "0000001101000001110101",
			5135 => "0000010101000001110101",
			5136 => "0000010111101000000100",
			5137 => "0000001101000001110101",
			5138 => "1111111101000001110101",
			5139 => "0001001011100000010000",
			5140 => "0010110110100000001000",
			5141 => "0011000100000100000100",
			5142 => "1111111101000001110101",
			5143 => "0000000101000001110101",
			5144 => "0000001010101100000100",
			5145 => "0000011101000001110101",
			5146 => "1111111101000001110101",
			5147 => "0000001101000001110101",
			5148 => "1111111101000001110101",
			5149 => "0001000011000001000000",
			5150 => "0011000100011000100100",
			5151 => "0001110110100100011000",
			5152 => "0000011101101000000100",
			5153 => "0000000101001000001001",
			5154 => "0000011110010100001100",
			5155 => "0010000010101100000100",
			5156 => "0000000101001000001001",
			5157 => "0011000100011000000100",
			5158 => "0000000101001000001001",
			5159 => "0000000101001000001001",
			5160 => "0011101100010000000100",
			5161 => "0000000101001000001001",
			5162 => "0000000101001000001001",
			5163 => "0000100000010000000100",
			5164 => "0000000101001000001001",
			5165 => "0010001100011100000100",
			5166 => "0000000101001000001001",
			5167 => "0000000101001000001001",
			5168 => "0001111000011000011000",
			5169 => "0010001010110000010000",
			5170 => "0001001100010000000100",
			5171 => "0000000101001000001001",
			5172 => "0010111011011100001000",
			5173 => "0000000101000100000100",
			5174 => "0000000101001000001001",
			5175 => "0000000101001000001001",
			5176 => "0000000101001000001001",
			5177 => "0010000110011100000100",
			5178 => "0000000101001000001001",
			5179 => "0000000101001000001001",
			5180 => "0000000101001000001001",
			5181 => "0000000000111000111100",
			5182 => "0010000111000100111000",
			5183 => "0000111111101000011100",
			5184 => "0011001001110000010000",
			5185 => "0000010110101000001000",
			5186 => "0010111100101100000100",
			5187 => "0000000101001000001001",
			5188 => "1111111101001000001001",
			5189 => "0000000011010000000100",
			5190 => "0000000101001000001001",
			5191 => "0000000101001000001001",
			5192 => "0000011001011000000100",
			5193 => "1111111101001000001001",
			5194 => "0001111000011000000100",
			5195 => "0000000101001000001001",
			5196 => "0000000101001000001001",
			5197 => "0000010100110100001100",
			5198 => "0011000100011000000100",
			5199 => "0000000101001000001001",
			5200 => "0010101010110000000100",
			5201 => "0000000101001000001001",
			5202 => "0000000101001000001001",
			5203 => "0010101000010100001000",
			5204 => "0011001010001100000100",
			5205 => "0000000101001000001001",
			5206 => "0000000101001000001001",
			5207 => "0011001001110100000100",
			5208 => "0000000101001000001001",
			5209 => "0000000101001000001001",
			5210 => "1111111101001000001001",
			5211 => "0000001010000000100000",
			5212 => "0001011110110100011100",
			5213 => "0001001101001000010000",
			5214 => "0000000000111000001000",
			5215 => "0010001111001000000100",
			5216 => "0000000101001000001001",
			5217 => "0000000101001000001001",
			5218 => "0000000000110000000100",
			5219 => "0000000101001000001001",
			5220 => "0000000101001000001001",
			5221 => "0010011111001100000100",
			5222 => "0000000101001000001001",
			5223 => "0011001000000000000100",
			5224 => "0000001101001000001001",
			5225 => "0000000101001000001001",
			5226 => "0000000101001000001001",
			5227 => "0010100101000100010100",
			5228 => "0000011001111000001100",
			5229 => "0001010111001000000100",
			5230 => "0000000101001000001001",
			5231 => "0000101100010000000100",
			5232 => "0000000101001000001001",
			5233 => "0000000101001000001001",
			5234 => "0001001010110100000100",
			5235 => "0000000101001000001001",
			5236 => "1111111101001000001001",
			5237 => "0010001111000100010000",
			5238 => "0011000011011100001000",
			5239 => "0000011001111000000100",
			5240 => "0000000101001000001001",
			5241 => "0000001101001000001001",
			5242 => "0000110101010100000100",
			5243 => "0000000101001000001001",
			5244 => "0000000101001000001001",
			5245 => "0001000001001100000100",
			5246 => "0000000101001000001001",
			5247 => "0001010000001100000100",
			5248 => "0000000101001000001001",
			5249 => "0000000101001000001001",
			5250 => "0001101101011000110100",
			5251 => "0000010101011100010100",
			5252 => "0001101001011000001000",
			5253 => "0000001100000100000100",
			5254 => "0000000101001111011111",
			5255 => "0000000101001111011111",
			5256 => "0001000101110000001000",
			5257 => "0010000010101100000100",
			5258 => "0000000101001111011111",
			5259 => "0000000101001111011111",
			5260 => "1111111101001111011111",
			5261 => "0000111010000100011000",
			5262 => "0011001011000000010000",
			5263 => "0001000111010100000100",
			5264 => "1111111101001111011111",
			5265 => "0010100010101100000100",
			5266 => "0000001101001111011111",
			5267 => "0011101001011100000100",
			5268 => "0000000101001111011111",
			5269 => "0000000101001111011111",
			5270 => "0010010101010000000100",
			5271 => "0000000101001111011111",
			5272 => "0000001101001111011111",
			5273 => "0000010101011100000100",
			5274 => "0000000101001111011111",
			5275 => "1111111101001111011111",
			5276 => "0001101000010001110000",
			5277 => "0011111001011100111100",
			5278 => "0000111000011000011100",
			5279 => "0011000000101000001100",
			5280 => "0001110100000000000100",
			5281 => "1111111101001111011111",
			5282 => "0001001110111000000100",
			5283 => "0000000101001111011111",
			5284 => "0000001101001111011111",
			5285 => "0011100111001000001000",
			5286 => "0011011110110000000100",
			5287 => "1111111101001111011111",
			5288 => "0000000101001111011111",
			5289 => "0011101011000000000100",
			5290 => "1111111101001111011111",
			5291 => "0000000101001111011111",
			5292 => "0000000011111100010000",
			5293 => "0000110000011100001000",
			5294 => "0000000010111100000100",
			5295 => "1111111101001111011111",
			5296 => "1111110101001111011111",
			5297 => "0011000100000000000100",
			5298 => "0000001101001111011111",
			5299 => "0000000101001111011111",
			5300 => "0001111001110000001000",
			5301 => "0011110001000000000100",
			5302 => "0000001101001111011111",
			5303 => "0000001101001111011111",
			5304 => "0001101001100100000100",
			5305 => "1111111101001111011111",
			5306 => "0000001101001111011111",
			5307 => "0001001100001100010100",
			5308 => "0000000010111100010000",
			5309 => "0000011101101000001000",
			5310 => "0011101001010100000100",
			5311 => "1111110101001111011111",
			5312 => "1111111101001111011111",
			5313 => "0001010001101000000100",
			5314 => "0000001101001111011111",
			5315 => "0000000101001111011111",
			5316 => "0000001101001111011111",
			5317 => "0001000010111000010000",
			5318 => "0001100100111100001000",
			5319 => "0000000011111100000100",
			5320 => "1111111101001111011111",
			5321 => "0000000101001111011111",
			5322 => "0011111000011100000100",
			5323 => "1111110101001111011111",
			5324 => "0000000101001111011111",
			5325 => "0001101001100100001000",
			5326 => "0000001111000100000100",
			5327 => "0000000101001111011111",
			5328 => "1111111101001111011111",
			5329 => "0010010000111100000100",
			5330 => "1111111101001111011111",
			5331 => "0000000101001111011111",
			5332 => "0011011010001000100000",
			5333 => "0010000110001000001100",
			5334 => "0000001010101100000100",
			5335 => "0000000101001111011111",
			5336 => "0001001001001100000100",
			5337 => "0000001101001111011111",
			5338 => "0000000101001111011111",
			5339 => "0001110110000100001000",
			5340 => "0010011100011000000100",
			5341 => "0000001101001111011111",
			5342 => "0000000101001111011111",
			5343 => "0010011010011000000100",
			5344 => "1111111101001111011111",
			5345 => "0001111110110000000100",
			5346 => "0000001101001111011111",
			5347 => "0000000101001111011111",
			5348 => "0011111000000100001100",
			5349 => "0011110110111000001000",
			5350 => "0011110010010100000100",
			5351 => "0000000101001111011111",
			5352 => "0000000101001111011111",
			5353 => "1111111101001111011111",
			5354 => "0000000111000000001100",
			5355 => "0011111000110100000100",
			5356 => "0000000101001111011111",
			5357 => "0001110100010000000100",
			5358 => "0000001101001111011111",
			5359 => "0000000101001111011111",
			5360 => "0000111000000100001000",
			5361 => "0000111011110000000100",
			5362 => "0000000101001111011111",
			5363 => "0000001101001111011111",
			5364 => "0011011110110100000100",
			5365 => "0000001101001111011111",
			5366 => "0000000101001111011111",
			5367 => "0000111001110100100100",
			5368 => "0010100001010100001000",
			5369 => "0010110100001000000100",
			5370 => "1111111101010011000001",
			5371 => "0000000101010011000001",
			5372 => "0010101001101000001100",
			5373 => "0001011010111100000100",
			5374 => "0000000101010011000001",
			5375 => "0001101001100100000100",
			5376 => "0000000101010011000001",
			5377 => "0000001101010011000001",
			5378 => "0000100000010000000100",
			5379 => "1111111101010011000001",
			5380 => "0000100110101100001000",
			5381 => "0011100111000000000100",
			5382 => "0000000101010011000001",
			5383 => "0000000101010011000001",
			5384 => "0000000101010011000001",
			5385 => "0011111100100100011000",
			5386 => "0010011111001100001000",
			5387 => "0010000111000100000100",
			5388 => "0000000101010011000001",
			5389 => "0000001101010011000001",
			5390 => "0000110001101000000100",
			5391 => "1111111101010011000001",
			5392 => "0000000110011000000100",
			5393 => "0000000101010011000001",
			5394 => "0001111000111000000100",
			5395 => "0000000101010011000001",
			5396 => "0000001101010011000001",
			5397 => "0001011010111000010000",
			5398 => "0011111111010000001100",
			5399 => "0000111010011100001000",
			5400 => "0011101000000000000100",
			5401 => "1111111101010011000001",
			5402 => "0000000101010011000001",
			5403 => "0000001101010011000001",
			5404 => "1111111101010011000001",
			5405 => "0001111000111000001100",
			5406 => "0000000010011000000100",
			5407 => "1111111101010011000001",
			5408 => "0011011011000000000100",
			5409 => "0000000101010011000001",
			5410 => "0000001101010011000001",
			5411 => "0011011000000000010000",
			5412 => "0000000000110000001000",
			5413 => "0000101001100000000100",
			5414 => "0000000101010011000001",
			5415 => "1111111101010011000001",
			5416 => "0010100110011100000100",
			5417 => "0000000101010011000001",
			5418 => "0000000101010011000001",
			5419 => "0010001111000100001000",
			5420 => "0001011000000000000100",
			5421 => "0000000101010011000001",
			5422 => "0000000101010011000001",
			5423 => "1111111101010011000001",
			5424 => "0000111001110100100100",
			5425 => "0001000010010000001000",
			5426 => "0011011000011000000100",
			5427 => "1111111101010111000101",
			5428 => "0000000101010111000101",
			5429 => "0000110100001000010000",
			5430 => "0000100000010000000100",
			5431 => "1111111101010111000101",
			5432 => "0000100000010000001000",
			5433 => "0010110011100000000100",
			5434 => "0000000101010111000101",
			5435 => "0000000101010111000101",
			5436 => "0000000101010111000101",
			5437 => "0001000101001100001000",
			5438 => "0001111101100000000100",
			5439 => "0000001101010111000101",
			5440 => "0000000101010111000101",
			5441 => "0000000101010111000101",
			5442 => "0011111100100100011100",
			5443 => "0000011001111000001000",
			5444 => "0010000111000100000100",
			5445 => "0000000101010111000101",
			5446 => "0000001101010111000101",
			5447 => "0011011011000000000100",
			5448 => "1111111101010111000101",
			5449 => "0011110000110100000100",
			5450 => "0000000101010111000101",
			5451 => "0011000100000000000100",
			5452 => "0000000101010111000101",
			5453 => "0011101000000000000100",
			5454 => "0000000101010111000101",
			5455 => "0000001101010111000101",
			5456 => "0011011011000000010000",
			5457 => "0011111111010000001000",
			5458 => "0001101011001100000100",
			5459 => "1111111101010111000101",
			5460 => "0000000101010111000101",
			5461 => "0000110000011100000100",
			5462 => "1111111101010111000101",
			5463 => "0000000101010111000101",
			5464 => "0011110101110000011000",
			5465 => "0001111001110000001000",
			5466 => "0000110100000100000100",
			5467 => "0000000101010111000101",
			5468 => "0000001101010111000101",
			5469 => "0000110010001000001000",
			5470 => "0010000001110100000100",
			5471 => "1111111101010111000101",
			5472 => "0000000101010111000101",
			5473 => "0001101010011000000100",
			5474 => "0000000101010111000101",
			5475 => "0000001101010111000101",
			5476 => "0000010111100100010000",
			5477 => "0000000010011000001000",
			5478 => "0011010110100100000100",
			5479 => "1111111101010111000101",
			5480 => "0000000101010111000101",
			5481 => "0011111001100000000100",
			5482 => "0000000101010111000101",
			5483 => "1111111101010111000101",
			5484 => "0010110000001100000100",
			5485 => "0000001101010111000101",
			5486 => "0000010000111100000100",
			5487 => "0000000101010111000101",
			5488 => "0000000101010111000101",
			5489 => "0001111001110000110100",
			5490 => "0011100100000100101000",
			5491 => "0000110000011100100000",
			5492 => "0001000100001100001000",
			5493 => "0011011011000000000100",
			5494 => "1111111101011011001001",
			5495 => "0000000101011011001001",
			5496 => "0000101100010000010000",
			5497 => "0010110011011100001000",
			5498 => "0000100010000100000100",
			5499 => "0000000101011011001001",
			5500 => "0000000101011011001001",
			5501 => "0011000100000000000100",
			5502 => "0000001101011011001001",
			5503 => "0000000101011011001001",
			5504 => "0001101111000000000100",
			5505 => "1111111101011011001001",
			5506 => "0000000101011011001001",
			5507 => "0010011001011000000100",
			5508 => "0000000101011011001001",
			5509 => "0000001101011011001001",
			5510 => "0000110101110100001000",
			5511 => "0001101001100100000100",
			5512 => "0000000101011011001001",
			5513 => "1111111101011011001001",
			5514 => "0000000101011011001001",
			5515 => "0001111001110000010100",
			5516 => "0011001000111100001100",
			5517 => "0001101101011000000100",
			5518 => "0000000101011011001001",
			5519 => "0011011110110000000100",
			5520 => "0000000101011011001001",
			5521 => "0000001101011011001001",
			5522 => "0001111001110000000100",
			5523 => "0000000101011011001001",
			5524 => "0000000101011011001001",
			5525 => "0011011000000000001000",
			5526 => "0001000010010000000100",
			5527 => "1111111101011011001001",
			5528 => "0000000101011011001001",
			5529 => "0010110000001100011000",
			5530 => "0001101001100100001000",
			5531 => "0010011101011100000100",
			5532 => "0000000101011011001001",
			5533 => "1111111101011011001001",
			5534 => "0000000011111100001000",
			5535 => "0000010111100100000100",
			5536 => "0000000101011011001001",
			5537 => "0000001101011011001001",
			5538 => "0001110110000100000100",
			5539 => "0000001101011011001001",
			5540 => "0000000101011011001001",
			5541 => "0001111110001100001100",
			5542 => "0001101000010000001000",
			5543 => "0001111101100000000100",
			5544 => "0000000101011011001001",
			5545 => "1111111101011011001001",
			5546 => "0000000101011011001001",
			5547 => "0000000010011000001000",
			5548 => "0000111010000100000100",
			5549 => "0000000101011011001001",
			5550 => "0000000101011011001001",
			5551 => "0010101010110000000100",
			5552 => "1111111101011011001001",
			5553 => "0000000101011011001001",
			5554 => "0000111001110100011000",
			5555 => "0010100001010100001000",
			5556 => "0000010111100100000100",
			5557 => "1111111101011110010101",
			5558 => "0000000101011110010101",
			5559 => "0001111101100000001100",
			5560 => "0010111001110000001000",
			5561 => "0010110100000000000100",
			5562 => "1111111101011110010101",
			5563 => "0000000101011110010101",
			5564 => "0000001101011110010101",
			5565 => "1111111101011110010101",
			5566 => "0000001001110001001100",
			5567 => "0000000011010000011100",
			5568 => "0000110000011100001000",
			5569 => "0000000011111100000100",
			5570 => "1111111101011110010101",
			5571 => "1111110101011110010101",
			5572 => "0001010100011000000100",
			5573 => "0000001101011110010101",
			5574 => "0000010111100100001000",
			5575 => "0000010111100100000100",
			5576 => "0000000101011110010101",
			5577 => "1111110101011110010101",
			5578 => "0001010001101000000100",
			5579 => "0000001101011110010101",
			5580 => "0000000101011110010101",
			5581 => "0000001110111100010000",
			5582 => "0010101010110000000100",
			5583 => "1111111101011110010101",
			5584 => "0011001111011100001000",
			5585 => "0010010000111100000100",
			5586 => "0000000101011110010101",
			5587 => "0000001101011110010101",
			5588 => "1111111101011110010101",
			5589 => "0010100101000100010000",
			5590 => "0011111001011100001000",
			5591 => "0010100110011100000100",
			5592 => "1111111101011110010101",
			5593 => "0000000101011110010101",
			5594 => "0000000111111000000100",
			5595 => "0000000101011110010101",
			5596 => "1111111101011110010101",
			5597 => "0011000110000100001000",
			5598 => "0001000010010000000100",
			5599 => "0000001101011110010101",
			5600 => "0000000101011110010101",
			5601 => "0010111110101000000100",
			5602 => "1111111101011110010101",
			5603 => "0000001101011110010101",
			5604 => "1111111101011110010101",
			5605 => "0000111001110100011100",
			5606 => "0001101011001100001000",
			5607 => "0000010111100100000100",
			5608 => "1111111101100010101001",
			5609 => "0000000101100010101001",
			5610 => "0011100001111100010000",
			5611 => "0000111101010100001000",
			5612 => "0000100111011000000100",
			5613 => "1111111101100010101001",
			5614 => "0000000101100010101001",
			5615 => "0010110101101100000100",
			5616 => "0000001101100010101001",
			5617 => "0000000101100010101001",
			5618 => "1111111101100010101001",
			5619 => "0011110101110000110100",
			5620 => "0001111001110000011100",
			5621 => "0011010100011000001100",
			5622 => "0011111110101000001000",
			5623 => "0001001000000100000100",
			5624 => "0000000101100010101001",
			5625 => "0000000101100010101001",
			5626 => "1111111101100010101001",
			5627 => "0000101100010100000100",
			5628 => "0000000101100010101001",
			5629 => "0011101110110000000100",
			5630 => "0000000101100010101001",
			5631 => "0001101101011000000100",
			5632 => "0000000101100010101001",
			5633 => "0000001101100010101001",
			5634 => "0000110100000100001000",
			5635 => "0001001011100000000100",
			5636 => "1111111101100010101001",
			5637 => "0000000101100010101001",
			5638 => "0001010110110100001100",
			5639 => "0011110010011100001000",
			5640 => "0011110000110100000100",
			5641 => "0000000101100010101001",
			5642 => "0000001101100010101001",
			5643 => "0000000101100010101001",
			5644 => "0000000101100010101001",
			5645 => "0000110001001000100000",
			5646 => "0011100111110000011100",
			5647 => "0001111001110000001100",
			5648 => "0000110101110100001000",
			5649 => "0001000010111000000100",
			5650 => "1111111101100010101001",
			5651 => "0000000101100010101001",
			5652 => "0000001101100010101001",
			5653 => "0011001000111000001000",
			5654 => "0001101001100100000100",
			5655 => "0000000101100010101001",
			5656 => "0000001101100010101001",
			5657 => "0001101111000000000100",
			5658 => "0000000101100010101001",
			5659 => "0000001101100010101001",
			5660 => "1111111101100010101001",
			5661 => "0011011101101100011000",
			5662 => "0010110000001100001000",
			5663 => "0001101111000000000100",
			5664 => "0000000101100010101001",
			5665 => "0000001101100010101001",
			5666 => "0000111001011100001000",
			5667 => "0001010001101000000100",
			5668 => "0000000101100010101001",
			5669 => "1111111101100010101001",
			5670 => "0001110100001000000100",
			5671 => "0000001101100010101001",
			5672 => "0000000101100010101001",
			5673 => "1111111101100010101001",
			5674 => "0001101101011000101100",
			5675 => "0000010001000100010100",
			5676 => "0010001001000100010000",
			5677 => "0001010110110100001100",
			5678 => "0001111100101000000100",
			5679 => "1111111101100110100101",
			5680 => "0010000000001000000100",
			5681 => "0000000101100110100101",
			5682 => "0000001101100110100101",
			5683 => "1111111101100110100101",
			5684 => "1111111101100110100101",
			5685 => "0000111010000100010100",
			5686 => "0000100110111100010000",
			5687 => "0000010111101000001100",
			5688 => "0010101010100000000100",
			5689 => "0000001101100110100101",
			5690 => "0011010101001000000100",
			5691 => "0000000101100110100101",
			5692 => "1111111101100110100101",
			5693 => "0000001101100110100101",
			5694 => "0000010101100110100101",
			5695 => "1111111101100110100101",
			5696 => "0010101011010101001100",
			5697 => "0001101000010000101100",
			5698 => "0001000010010100011000",
			5699 => "0011001000000000001100",
			5700 => "0010011011111100000100",
			5701 => "1111111101100110100101",
			5702 => "0010011001111100000100",
			5703 => "0000001101100110100101",
			5704 => "0000000101100110100101",
			5705 => "0010000001010000001000",
			5706 => "0000100111010100000100",
			5707 => "0000000101100110100101",
			5708 => "0000001101100110100101",
			5709 => "1111111101100110100101",
			5710 => "0001101011001100000100",
			5711 => "1111111101100110100101",
			5712 => "0011111001010000001000",
			5713 => "0001111101100000000100",
			5714 => "0000001101100110100101",
			5715 => "1111111101100110100101",
			5716 => "0000110001011000000100",
			5717 => "1111111101100110100101",
			5718 => "0000000101100110100101",
			5719 => "0001111111011100010000",
			5720 => "0001000111011100001100",
			5721 => "0010011010011000000100",
			5722 => "0000000101100110100101",
			5723 => "0010001100000100000100",
			5724 => "0000000101100110100101",
			5725 => "0000001101100110100101",
			5726 => "0000000101100110100101",
			5727 => "0011100011010100001100",
			5728 => "0010010111110100001000",
			5729 => "0011110110001100000100",
			5730 => "0000000101100110100101",
			5731 => "0000001101100110100101",
			5732 => "1111111101100110100101",
			5733 => "0000001101100110100101",
			5734 => "0001010100011000000100",
			5735 => "0000000101100110100101",
			5736 => "1111111101100110100101",
			5737 => "0001111001110000101100",
			5738 => "0001101001100100100000",
			5739 => "0011100100000100011000",
			5740 => "0011010100011000000100",
			5741 => "0000000101101011011001",
			5742 => "0011000100000000001000",
			5743 => "0001101001100100000100",
			5744 => "0000000101101011011001",
			5745 => "0000000101101011011001",
			5746 => "0000101100010000001000",
			5747 => "0001101101011000000100",
			5748 => "0000000101101011011001",
			5749 => "0000000101101011011001",
			5750 => "0000000101101011011001",
			5751 => "0010001011010100000100",
			5752 => "0000000101101011011001",
			5753 => "1111111101101011011001",
			5754 => "0011011000000000001000",
			5755 => "0001111000111000000100",
			5756 => "0000000101101011011001",
			5757 => "0000000101101011011001",
			5758 => "0000000101101011011001",
			5759 => "0000101111010100101000",
			5760 => "0001101011001100011000",
			5761 => "0011001110001100001000",
			5762 => "0010110101101100000100",
			5763 => "0000000101101011011001",
			5764 => "0000000101101011011001",
			5765 => "0010110101100100001100",
			5766 => "0011101011011100000100",
			5767 => "0000000101101011011001",
			5768 => "0000010001111000000100",
			5769 => "0000000101101011011001",
			5770 => "0000000101101011011001",
			5771 => "0000000101101011011001",
			5772 => "0010100111110100000100",
			5773 => "0000000101101011011001",
			5774 => "0011010011100000000100",
			5775 => "0000000101101011011001",
			5776 => "0011100001101000000100",
			5777 => "0000000101101011011001",
			5778 => "0000001101101011011001",
			5779 => "0010111011110100100100",
			5780 => "0010000010101000011100",
			5781 => "0000101000000100010000",
			5782 => "0000000011010000001000",
			5783 => "0000011001011000000100",
			5784 => "0000000101101011011001",
			5785 => "0000000101101011011001",
			5786 => "0001111101111000000100",
			5787 => "0000000101101011011001",
			5788 => "0000000101101011011001",
			5789 => "0011110011001100001000",
			5790 => "0011001001110100000100",
			5791 => "0000001101101011011001",
			5792 => "0000000101101011011001",
			5793 => "0000000101101011011001",
			5794 => "0000011101101000000100",
			5795 => "0000000101101011011001",
			5796 => "0000000101101011011001",
			5797 => "0011100011110100011100",
			5798 => "0000010001111000001100",
			5799 => "0001110000011100000100",
			5800 => "0000000101101011011001",
			5801 => "0011101011101100000100",
			5802 => "0000000101101011011001",
			5803 => "0000000101101011011001",
			5804 => "0001101000010000001000",
			5805 => "0000001010101100000100",
			5806 => "0000000101101011011001",
			5807 => "0000000101101011011001",
			5808 => "0000001010101100000100",
			5809 => "0000000101101011011001",
			5810 => "0000000101101011011001",
			5811 => "0001100000001000000100",
			5812 => "0000000101101011011001",
			5813 => "0000000101101011011001",
			5814 => "0001011010111000100100",
			5815 => "0001001111100000001100",
			5816 => "0001111001110000000100",
			5817 => "1111111101110000001101",
			5818 => "0001111101100000000100",
			5819 => "0000000101110000001101",
			5820 => "0000000101110000001101",
			5821 => "0011010001111100000100",
			5822 => "1111111101110000001101",
			5823 => "0011000000101000001000",
			5824 => "0001101011001100000100",
			5825 => "0000000101110000001101",
			5826 => "0000001101110000001101",
			5827 => "0001101001100100001000",
			5828 => "0001000111011100000100",
			5829 => "1111111101110000001101",
			5830 => "0000000101110000001101",
			5831 => "0000001101110000001101",
			5832 => "0001010100011000100000",
			5833 => "0011011011000000010100",
			5834 => "0000000011010000000100",
			5835 => "1111111101110000001101",
			5836 => "0000101100010000001000",
			5837 => "0001101101011000000100",
			5838 => "0000000101110000001101",
			5839 => "0000001101110000001101",
			5840 => "0010011101011100000100",
			5841 => "0000000101110000001101",
			5842 => "0000000101110000001101",
			5843 => "0001101101011000000100",
			5844 => "0000000101110000001101",
			5845 => "0001111101100000000100",
			5846 => "0000001101110000001101",
			5847 => "0000000101110000001101",
			5848 => "0011011000000000011100",
			5849 => "0001000010100100010000",
			5850 => "0001111000111000000100",
			5851 => "0000000101110000001101",
			5852 => "0000011001111000000100",
			5853 => "0000000101110000001101",
			5854 => "0000000011111100000100",
			5855 => "0000000101110000001101",
			5856 => "1111111101110000001101",
			5857 => "0000100111010100001000",
			5858 => "0011001100110000000100",
			5859 => "0000001101110000001101",
			5860 => "0000000101110000001101",
			5861 => "0000000101110000001101",
			5862 => "0000100010000100011100",
			5863 => "0010100001010000010000",
			5864 => "0000110111110000001000",
			5865 => "0001000011000000000100",
			5866 => "0000000101110000001101",
			5867 => "1111111101110000001101",
			5868 => "0000011101101000000100",
			5869 => "0000000101110000001101",
			5870 => "0000001101110000001101",
			5871 => "0011001001110000001000",
			5872 => "0001011000000000000100",
			5873 => "0000001101110000001101",
			5874 => "0000000101110000001101",
			5875 => "0000000101110000001101",
			5876 => "0011100101100100010000",
			5877 => "0001101001100100001000",
			5878 => "0011101000000000000100",
			5879 => "0000000101110000001101",
			5880 => "1111111101110000001101",
			5881 => "0011010001101000000100",
			5882 => "0000001101110000001101",
			5883 => "1111111101110000001101",
			5884 => "0011011100111000001000",
			5885 => "0000110110111000000100",
			5886 => "0000000101110000001101",
			5887 => "0000000101110000001101",
			5888 => "0011000101110100000100",
			5889 => "1111111101110000001101",
			5890 => "0000000101110000001101",
			5891 => "0000110111110001010100",
			5892 => "0010100001010000100000",
			5893 => "0011111001010000010100",
			5894 => "0011101010001100001000",
			5895 => "0001101001011000000100",
			5896 => "0000000101110101101001",
			5897 => "0000000101110101101001",
			5898 => "0000010111100100000100",
			5899 => "0000000101110101101001",
			5900 => "0010000000001000000100",
			5901 => "0000000101110101101001",
			5902 => "0000000101110101101001",
			5903 => "0011001100001000000100",
			5904 => "0000000101110101101001",
			5905 => "0011010001101000000100",
			5906 => "1111111101110101101001",
			5907 => "0000000101110101101001",
			5908 => "0001000101000000001000",
			5909 => "0000110000011100000100",
			5910 => "0000000101110101101001",
			5911 => "0000001101110101101001",
			5912 => "0001000011001100010000",
			5913 => "0001110100000000000100",
			5914 => "0000000101110101101001",
			5915 => "0000010110101000001000",
			5916 => "0011000000101000000100",
			5917 => "0000000101110101101001",
			5918 => "1111111101110101101001",
			5919 => "0000000101110101101001",
			5920 => "0001101001100100010000",
			5921 => "0000101110110100001000",
			5922 => "0000111001110100000100",
			5923 => "0000000101110101101001",
			5924 => "0000000101110101101001",
			5925 => "0001110100000000000100",
			5926 => "0000000101110101101001",
			5927 => "1111111101110101101001",
			5928 => "0011010001101000001000",
			5929 => "0000100110101100000100",
			5930 => "0000000101110101101001",
			5931 => "0000000101110101101001",
			5932 => "0000000101110101101001",
			5933 => "0011111100010000100000",
			5934 => "0011011110000100011100",
			5935 => "0001001101001000010100",
			5936 => "0000010111100100001000",
			5937 => "0011001000111000000100",
			5938 => "0000000101110101101001",
			5939 => "0000000101110101101001",
			5940 => "0010011001111100001000",
			5941 => "0010000010101100000100",
			5942 => "0000000101110101101001",
			5943 => "0000000101110101101001",
			5944 => "0000000101110101101001",
			5945 => "0001110101101100000100",
			5946 => "0000000101110101101001",
			5947 => "0000000101110101101001",
			5948 => "0000000101110101101001",
			5949 => "0010011100011000010000",
			5950 => "0000101111101000001000",
			5951 => "0011010111010000000100",
			5952 => "0000000101110101101001",
			5953 => "1111111101110101101001",
			5954 => "0000001011000100000100",
			5955 => "0000000101110101101001",
			5956 => "0000000101110101101001",
			5957 => "0011011110101100001100",
			5958 => "0011000011011100000100",
			5959 => "0000000101110101101001",
			5960 => "0000101000100000000100",
			5961 => "0000000101110101101001",
			5962 => "0000001101110101101001",
			5963 => "0000010111101000010000",
			5964 => "0011111000110100001000",
			5965 => "0001100100111100000100",
			5966 => "0000000101110101101001",
			5967 => "1111111101110101101001",
			5968 => "0000000000111000000100",
			5969 => "0000000101110101101001",
			5970 => "0000000101110101101001",
			5971 => "0001001000001000001000",
			5972 => "0010101000100100000100",
			5973 => "0000000101110101101001",
			5974 => "0000000101110101101001",
			5975 => "0011110101000000000100",
			5976 => "0000000101110101101001",
			5977 => "0000000101110101101001",
			5978 => "0000110010001001000000",
			5979 => "0010111100101100110100",
			5980 => "0000000011010000010100",
			5981 => "0011011000000000001100",
			5982 => "0010001001101000000100",
			5983 => "0000000101111010011101",
			5984 => "0001000010110000000100",
			5985 => "1111111101111010011101",
			5986 => "0000000101111010011101",
			5987 => "0001001000110100000100",
			5988 => "0000000101111010011101",
			5989 => "0000000101111010011101",
			5990 => "0011111110010000011100",
			5991 => "0000111010011100010000",
			5992 => "0001000100001100001000",
			5993 => "0000110001101000000100",
			5994 => "1111111101111010011101",
			5995 => "0000000101111010011101",
			5996 => "0010110101101100000100",
			5997 => "0000000101111010011101",
			5998 => "0000000101111010011101",
			5999 => "0000101100010000000100",
			6000 => "0000001101111010011101",
			6001 => "0000110001011000000100",
			6002 => "0000000101111010011101",
			6003 => "0000000101111010011101",
			6004 => "1111111101111010011101",
			6005 => "0011111111010000000100",
			6006 => "0000000101111010011101",
			6007 => "0000100111010100000100",
			6008 => "1111111101111010011101",
			6009 => "0000000101111010011101",
			6010 => "0001011001001000001100",
			6011 => "0000010110101000000100",
			6012 => "0000000101111010011101",
			6013 => "0000001101010000000100",
			6014 => "0000000101111010011101",
			6015 => "0000001101111010011101",
			6016 => "0010110111001000011100",
			6017 => "0001101000010000010100",
			6018 => "0001111101100000001000",
			6019 => "0010111110001100000100",
			6020 => "0000000101111010011101",
			6021 => "0000000101111010011101",
			6022 => "0000000000111000001000",
			6023 => "0000011111001100000100",
			6024 => "1111111101111010011101",
			6025 => "0000000101111010011101",
			6026 => "0000000101111010011101",
			6027 => "0010111010111100000100",
			6028 => "0000001101111010011101",
			6029 => "0000000101111010011101",
			6030 => "0010111011000000010100",
			6031 => "0001111101111000001000",
			6032 => "0000100011000000000100",
			6033 => "0000000101111010011101",
			6034 => "0000000101111010011101",
			6035 => "0000111001010100000100",
			6036 => "0000000101111010011101",
			6037 => "0001000000100000000100",
			6038 => "0000001101111010011101",
			6039 => "0000000101111010011101",
			6040 => "0000001111000100010000",
			6041 => "0011110110111100001000",
			6042 => "0001010110110100000100",
			6043 => "0000000101111010011101",
			6044 => "0000000101111010011101",
			6045 => "0001111001001000000100",
			6046 => "0000000101111010011101",
			6047 => "0000000101111010011101",
			6048 => "0010001001101000001000",
			6049 => "0000110110111000000100",
			6050 => "1111111101111010011101",
			6051 => "0000000101111010011101",
			6052 => "0000100011110100000100",
			6053 => "0000000101111010011101",
			6054 => "0000000101111010011101",
			6055 => "0010110011011100011000",
			6056 => "0000100111011000010000",
			6057 => "0001011101010100000100",
			6058 => "1111111101111110011001",
			6059 => "0010110011011100000100",
			6060 => "0000000101111110011001",
			6061 => "0001011101010100000100",
			6062 => "0000000101111110011001",
			6063 => "0000000101111110011001",
			6064 => "0010001111000100000100",
			6065 => "1111111101111110011001",
			6066 => "0000001101111110011001",
			6067 => "0010101011010101100000",
			6068 => "0001101000010000111000",
			6069 => "0011000100000000011000",
			6070 => "0001101011001100001100",
			6071 => "0011111100100100001000",
			6072 => "0010101010110000000100",
			6073 => "1111111101111110011001",
			6074 => "0000001101111110011001",
			6075 => "1111111101111110011001",
			6076 => "0000101100000000000100",
			6077 => "0000001101111110011001",
			6078 => "0011011000000000000100",
			6079 => "1111111101111110011001",
			6080 => "0000001101111110011001",
			6081 => "0000111000011000010000",
			6082 => "0010111100110000001000",
			6083 => "0001101011001100000100",
			6084 => "1111111101111110011001",
			6085 => "0000001101111110011001",
			6086 => "0010001000110000000100",
			6087 => "1111111101111110011001",
			6088 => "0000000101111110011001",
			6089 => "0011100110100100001000",
			6090 => "0010111100101100000100",
			6091 => "0000001101111110011001",
			6092 => "1111111101111110011001",
			6093 => "0000110000011100000100",
			6094 => "1111111101111110011001",
			6095 => "0000000101111110011001",
			6096 => "0011010111111100010000",
			6097 => "0010000110001000000100",
			6098 => "0000001101111110011001",
			6099 => "0010111010111100000100",
			6100 => "0000001101111110011001",
			6101 => "0000011111001100000100",
			6102 => "1111111101111110011001",
			6103 => "0000000101111110011001",
			6104 => "0011111000000100001100",
			6105 => "0010110010001000000100",
			6106 => "0000000101111110011001",
			6107 => "0011101100111000000100",
			6108 => "0000000101111110011001",
			6109 => "1111111101111110011001",
			6110 => "0011000100011000000100",
			6111 => "1111111101111110011001",
			6112 => "0010111011110100000100",
			6113 => "0000001101111110011001",
			6114 => "0000000101111110011001",
			6115 => "0011001000111100000100",
			6116 => "0000000101111110011001",
			6117 => "1111111101111110011001",
			6118 => "0011011110110000010100",
			6119 => "0001000000101100000100",
			6120 => "1111111110000010110101",
			6121 => "0000000011011100001000",
			6122 => "0010100001010100000100",
			6123 => "0000000110000010110101",
			6124 => "0000000110000010110101",
			6125 => "0000100111010100000100",
			6126 => "0000000110000010110101",
			6127 => "0000000110000010110101",
			6128 => "0001001000001000110000",
			6129 => "0000010110101000001100",
			6130 => "0001000110001100000100",
			6131 => "1111111110000010110101",
			6132 => "0001011110110000000100",
			6133 => "0000000110000010110101",
			6134 => "0000000110000010110101",
			6135 => "0011000100000000001000",
			6136 => "0000110010001000000100",
			6137 => "0000000110000010110101",
			6138 => "0000001110000010110101",
			6139 => "0011000100011000001100",
			6140 => "0001111000111000000100",
			6141 => "0000001110000010110101",
			6142 => "0001010001000000000100",
			6143 => "0000000110000010110101",
			6144 => "1111111110000010110101",
			6145 => "0010010101010000001000",
			6146 => "0001110101100100000100",
			6147 => "1111111110000010110101",
			6148 => "0000000110000010110101",
			6149 => "0010011010100100000100",
			6150 => "0000001110000010110101",
			6151 => "0000000110000010110101",
			6152 => "0001111100101000011000",
			6153 => "0010101010110000000100",
			6154 => "1111111110000010110101",
			6155 => "0000111001011100010000",
			6156 => "0000101111010100001000",
			6157 => "0000111011011100000100",
			6158 => "0000000110000010110101",
			6159 => "0000001110000010110101",
			6160 => "0010100101000100000100",
			6161 => "0000000110000010110101",
			6162 => "0000000110000010110101",
			6163 => "0000001110000010110101",
			6164 => "0000101000000100010100",
			6165 => "0010101100011100001100",
			6166 => "0001000000010100000100",
			6167 => "1111111110000010110101",
			6168 => "0010101001000100000100",
			6169 => "0000000110000010110101",
			6170 => "0000000110000010110101",
			6171 => "0001001001000000000100",
			6172 => "0000000110000010110101",
			6173 => "0000000110000010110101",
			6174 => "0010000001110100010000",
			6175 => "0011000001101000001000",
			6176 => "0010100001010000000100",
			6177 => "0000000110000010110101",
			6178 => "0000001110000010110101",
			6179 => "0001011110110100000100",
			6180 => "1111111110000010110101",
			6181 => "0000000110000010110101",
			6182 => "0011100010100100001000",
			6183 => "0000101101001000000100",
			6184 => "0000000110000010110101",
			6185 => "1111111110000010110101",
			6186 => "0011011100111000000100",
			6187 => "0000000110000010110101",
			6188 => "0000000110000010110101",
			6189 => "0010110011011100011000",
			6190 => "0000100111011000010000",
			6191 => "0001011101010100000100",
			6192 => "1111111110000110111001",
			6193 => "0010110011011100000100",
			6194 => "0000000110000110111001",
			6195 => "0001011101010100000100",
			6196 => "0000000110000110111001",
			6197 => "0000000110000110111001",
			6198 => "0010001111000100000100",
			6199 => "1111111110000110111001",
			6200 => "0000001110000110111001",
			6201 => "0010101011010101100100",
			6202 => "0001101000010000110100",
			6203 => "0011000100000000011000",
			6204 => "0001000010111000001100",
			6205 => "0000010110101000001000",
			6206 => "0011110101110000000100",
			6207 => "0000000110000110111001",
			6208 => "1111110110000110111001",
			6209 => "0000001110000110111001",
			6210 => "0001010111001000001000",
			6211 => "0011110110100000000100",
			6212 => "0000001110000110111001",
			6213 => "1111111110000110111001",
			6214 => "0000001110000110111001",
			6215 => "0011011011000000001100",
			6216 => "0011000100000000000100",
			6217 => "1111110110000110111001",
			6218 => "0001000010100100000100",
			6219 => "1111111110000110111001",
			6220 => "0000000110000110111001",
			6221 => "0010110110000100001000",
			6222 => "0001101011001100000100",
			6223 => "0000000110000110111001",
			6224 => "0000001110000110111001",
			6225 => "0001001100001100000100",
			6226 => "0000000110000110111001",
			6227 => "0000000110000110111001",
			6228 => "0011010111111100010100",
			6229 => "0010000110001000000100",
			6230 => "0000001110000110111001",
			6231 => "0011000110000100001000",
			6232 => "0010001111001000000100",
			6233 => "0000000110000110111001",
			6234 => "0000001110000110111001",
			6235 => "0000010101011100000100",
			6236 => "1111111110000110111001",
			6237 => "0000000110000110111001",
			6238 => "0011111000000100001100",
			6239 => "0010110010001000000100",
			6240 => "0000000110000110111001",
			6241 => "0011101100111000000100",
			6242 => "0000000110000110111001",
			6243 => "1111111110000110111001",
			6244 => "0000000111000000001000",
			6245 => "0011111000110100000100",
			6246 => "0000000110000110111001",
			6247 => "0000001110000110111001",
			6248 => "0010101001000100000100",
			6249 => "1111111110000110111001",
			6250 => "0000000110000110111001",
			6251 => "0001010100011000000100",
			6252 => "0000000110000110111001",
			6253 => "1111111110000110111001",
			6254 => "0001001000000101001000",
			6255 => "0001001111100100011000",
			6256 => "0000111010000100010100",
			6257 => "0010100010101100010000",
			6258 => "0010110101100100001100",
			6259 => "0000011011111100000100",
			6260 => "0000000110001100001101",
			6261 => "0010110000011100000100",
			6262 => "0000000110001100001101",
			6263 => "0000000110001100001101",
			6264 => "0000000110001100001101",
			6265 => "0000000110001100001101",
			6266 => "0000000110001100001101",
			6267 => "0000111100111000100000",
			6268 => "0001111100101000010000",
			6269 => "0011001001110000001100",
			6270 => "0000111011011100000100",
			6271 => "0000000110001100001101",
			6272 => "0001110101101100000100",
			6273 => "0000000110001100001101",
			6274 => "0000000110001100001101",
			6275 => "0000000110001100001101",
			6276 => "0011001000000000001100",
			6277 => "0010011010100100001000",
			6278 => "0010010111101100000100",
			6279 => "0000001110001100001101",
			6280 => "0000000110001100001101",
			6281 => "0000000110001100001101",
			6282 => "0000000110001100001101",
			6283 => "0011001001001000001000",
			6284 => "0000100011000000000100",
			6285 => "0000000110001100001101",
			6286 => "0000000110001100001101",
			6287 => "0011000001101000000100",
			6288 => "0000000110001100001101",
			6289 => "0000000110001100001101",
			6290 => "0001001000110100001100",
			6291 => "0000010001111000001000",
			6292 => "0000000010011000000100",
			6293 => "1111111110001100001101",
			6294 => "0000000110001100001101",
			6295 => "0000000110001100001101",
			6296 => "0011111110000000111100",
			6297 => "0001110101101100011100",
			6298 => "0000110000011100010000",
			6299 => "0010110101101100001000",
			6300 => "0001001001001100000100",
			6301 => "0000000110001100001101",
			6302 => "0000000110001100001101",
			6303 => "0000100010000000000100",
			6304 => "0000000110001100001101",
			6305 => "0000000110001100001101",
			6306 => "0010100001010000000100",
			6307 => "0000000110001100001101",
			6308 => "0000101100000000000100",
			6309 => "0000001110001100001101",
			6310 => "0000000110001100001101",
			6311 => "0010100101000100010000",
			6312 => "0010010111101100001000",
			6313 => "0010101000100100000100",
			6314 => "0000000110001100001101",
			6315 => "1111111110001100001101",
			6316 => "0010110101110100000100",
			6317 => "0000000110001100001101",
			6318 => "0000000110001100001101",
			6319 => "0010100001110000001000",
			6320 => "0011101011011100000100",
			6321 => "0000000110001100001101",
			6322 => "0000000110001100001101",
			6323 => "0001110101101100000100",
			6324 => "0000000110001100001101",
			6325 => "0000000110001100001101",
			6326 => "0010100110011100010000",
			6327 => "0000001010101100000100",
			6328 => "0000000110001100001101",
			6329 => "0001110111010000000100",
			6330 => "0000000110001100001101",
			6331 => "0001110000011100000100",
			6332 => "0000000110001100001101",
			6333 => "0000000110001100001101",
			6334 => "0011100010100100001000",
			6335 => "0000101101001000000100",
			6336 => "0000000110001100001101",
			6337 => "1111111110001100001101",
			6338 => "0000000110001100001101",
			6339 => "0001101001100101001000",
			6340 => "0001010111001000000100",
			6341 => "1111111110010000111001",
			6342 => "0011111110000100011100",
			6343 => "0001101101011000001100",
			6344 => "0000100110100000001000",
			6345 => "0000000110011000000100",
			6346 => "0000000110010000111001",
			6347 => "0000000110010000111001",
			6348 => "1111111110010000111001",
			6349 => "0001000010111000000100",
			6350 => "0000000110010000111001",
			6351 => "0000111001110100000100",
			6352 => "0000000110010000111001",
			6353 => "0011001001110000000100",
			6354 => "0000001110010000111001",
			6355 => "0000000110010000111001",
			6356 => "0001001000000100010100",
			6357 => "0010011110010100001000",
			6358 => "0001001011110000000100",
			6359 => "0000000110010000111001",
			6360 => "0000001110010000111001",
			6361 => "0010011000010000000100",
			6362 => "1111111110010000111001",
			6363 => "0011001011000000000100",
			6364 => "0000000110010000111001",
			6365 => "0000000110010000111001",
			6366 => "0000101100010000001100",
			6367 => "0000100110010000000100",
			6368 => "0000000110010000111001",
			6369 => "0011001000111000000100",
			6370 => "0000000110010000111001",
			6371 => "0000000110010000111001",
			6372 => "0011000111001000000100",
			6373 => "1111111110010000111001",
			6374 => "0000000110010000111001",
			6375 => "0001111101100000011100",
			6376 => "0010111100101100011000",
			6377 => "0011111110010000010100",
			6378 => "0011001000111100010000",
			6379 => "0011011110110000001000",
			6380 => "0000100010000100000100",
			6381 => "0000000110010000111001",
			6382 => "0000000110010000111001",
			6383 => "0010011111001100000100",
			6384 => "0000000110010000111001",
			6385 => "0000001110010000111001",
			6386 => "0000000110010000111001",
			6387 => "0000000110010000111001",
			6388 => "0000001110010000111001",
			6389 => "0011000100000000001000",
			6390 => "0010001011010100000100",
			6391 => "0000000110010000111001",
			6392 => "1111111110010000111001",
			6393 => "0000000111111000011100",
			6394 => "0010101100011100010000",
			6395 => "0010000111000100001000",
			6396 => "0010000110001000000100",
			6397 => "0000000110010000111001",
			6398 => "0000000110010000111001",
			6399 => "0011110110010000000100",
			6400 => "0000000110010000111001",
			6401 => "1111111110010000111001",
			6402 => "0011001000000000000100",
			6403 => "0000001110010000111001",
			6404 => "0011110000010100000100",
			6405 => "1111111110010000111001",
			6406 => "0000000110010000111001",
			6407 => "0001111101100000000100",
			6408 => "0000000110010000111001",
			6409 => "0000110011011000000100",
			6410 => "1111111110010000111001",
			6411 => "0010100010101000000100",
			6412 => "0000000110010000111001",
			6413 => "0000000110010000111001",
			6414 => "0000111011000000010100",
			6415 => "0001101001100100000100",
			6416 => "1111111110010101111101",
			6417 => "0010110011011100000100",
			6418 => "0000000110010101111101",
			6419 => "0000100111011000000100",
			6420 => "0000001110010101111101",
			6421 => "0010101111001000000100",
			6422 => "0000000110010101111101",
			6423 => "0000000110010101111101",
			6424 => "0001100100111101000100",
			6425 => "0010110110110100110000",
			6426 => "0001101100011000010000",
			6427 => "0010010101011100001100",
			6428 => "0000010110101000000100",
			6429 => "1111111110010101111101",
			6430 => "0000001010100000000100",
			6431 => "0000000110010101111101",
			6432 => "0000001110010101111101",
			6433 => "1111111110010101111101",
			6434 => "0001000011000000010000",
			6435 => "0010010111101100001000",
			6436 => "0010011011111100000100",
			6437 => "1111111110010101111101",
			6438 => "0000001110010101111101",
			6439 => "0010100111110100000100",
			6440 => "1111111110010101111101",
			6441 => "0000001110010101111101",
			6442 => "0011111001010000001000",
			6443 => "0001001111100000000100",
			6444 => "0000000110010101111101",
			6445 => "0000001110010101111101",
			6446 => "0011011000000000000100",
			6447 => "1111111110010101111101",
			6448 => "0000000110010101111101",
			6449 => "0000011110010100001100",
			6450 => "0011111011101100000100",
			6451 => "1111111110010101111101",
			6452 => "0000010101011100000100",
			6453 => "0000000110010101111101",
			6454 => "0000001110010101111101",
			6455 => "0010000001010100000100",
			6456 => "1111111110010101111101",
			6457 => "1111110110010101111101",
			6458 => "0001010001000000011100",
			6459 => "0001000111011100010000",
			6460 => "0011100011001000001000",
			6461 => "0010110001111100000100",
			6462 => "0000001110010101111101",
			6463 => "0000000110010101111101",
			6464 => "0010000001010100000100",
			6465 => "0000000110010101111101",
			6466 => "0000001110010101111101",
			6467 => "0010010001000100000100",
			6468 => "0000001110010101111101",
			6469 => "0001100101010000000100",
			6470 => "1111111110010101111101",
			6471 => "0000000110010101111101",
			6472 => "0011111000000100010100",
			6473 => "0010010011101000001100",
			6474 => "0011010111111100000100",
			6475 => "0000000110010101111101",
			6476 => "0011111110000000000100",
			6477 => "1111111110010101111101",
			6478 => "0000000110010101111101",
			6479 => "0011110110111000000100",
			6480 => "0000001110010101111101",
			6481 => "1111111110010101111101",
			6482 => "0001000000010100010000",
			6483 => "0000011101011000001000",
			6484 => "0011111000110100000100",
			6485 => "0000000110010101111101",
			6486 => "0000001110010101111101",
			6487 => "0011011110110100000100",
			6488 => "0000000110010101111101",
			6489 => "1111111110010101111101",
			6490 => "0000001011000100001000",
			6491 => "0001000011101100000100",
			6492 => "0000000110010101111101",
			6493 => "0000000110010101111101",
			6494 => "1111111110010101111101",
			6495 => "0010110011011100001000",
			6496 => "0000100111011000000100",
			6497 => "1111111110011001110001",
			6498 => "0000000110011001110001",
			6499 => "0011001100001000010100",
			6500 => "0001000010110000001000",
			6501 => "0000110101110100000100",
			6502 => "1111111110011001110001",
			6503 => "0000000110011001110001",
			6504 => "0001011010111100000100",
			6505 => "0000000110011001110001",
			6506 => "0001101011001100000100",
			6507 => "0000000110011001110001",
			6508 => "0000001110011001110001",
			6509 => "0001001000000100100100",
			6510 => "0001011000000000001000",
			6511 => "0001101011001100000100",
			6512 => "0000000110011001110001",
			6513 => "0000001110011001110001",
			6514 => "0000110001001000001100",
			6515 => "0011110010110100001000",
			6516 => "0011000110000100000100",
			6517 => "0000000110011001110001",
			6518 => "0000000110011001110001",
			6519 => "1111111110011001110001",
			6520 => "0000000111000100001000",
			6521 => "0000101000100000000100",
			6522 => "0000000110011001110001",
			6523 => "1111111110011001110001",
			6524 => "0001011100100100000100",
			6525 => "0000000110011001110001",
			6526 => "0000000110011001110001",
			6527 => "0001100100111100011100",
			6528 => "0010110110000100001100",
			6529 => "0011011110110000000100",
			6530 => "0000000110011001110001",
			6531 => "0000100111011000000100",
			6532 => "0000001110011001110001",
			6533 => "0000000110011001110001",
			6534 => "0001000110001100001000",
			6535 => "0000000010111100000100",
			6536 => "1111111110011001110001",
			6537 => "0000000110011001110001",
			6538 => "0000111001010100000100",
			6539 => "0000000110011001110001",
			6540 => "0000000110011001110001",
			6541 => "0011000110000100010000",
			6542 => "0000000011010000001000",
			6543 => "0001010001101000000100",
			6544 => "0000000110011001110001",
			6545 => "0000000110011001110001",
			6546 => "0010110110000100000100",
			6547 => "0000000110011001110001",
			6548 => "0000001110011001110001",
			6549 => "0011101011101100001000",
			6550 => "0001001000001000000100",
			6551 => "0000000110011001110001",
			6552 => "1111111110011001110001",
			6553 => "0011011010001000000100",
			6554 => "0000000110011001110001",
			6555 => "0000000110011001110001",
			6556 => "0001010111100010001000",
			6557 => "0001111110110001001100",
			6558 => "0010000110001000011000",
			6559 => "0011000100000000001000",
			6560 => "0001101011001100000100",
			6561 => "0000000110100000011101",
			6562 => "0000000110100000011101",
			6563 => "0011111001010000000100",
			6564 => "0000000110100000011101",
			6565 => "0000101100010100000100",
			6566 => "0000000110100000011101",
			6567 => "0001101000010000000100",
			6568 => "1111111110100000011101",
			6569 => "0000000110100000011101",
			6570 => "0000111011011100011100",
			6571 => "0011111111010000010000",
			6572 => "0000111001110100001000",
			6573 => "0011110110100000000100",
			6574 => "0000000110100000011101",
			6575 => "0000000110100000011101",
			6576 => "0000010110101000000100",
			6577 => "0000000110100000011101",
			6578 => "0000000110100000011101",
			6579 => "0001111000111000000100",
			6580 => "0000000110100000011101",
			6581 => "0001101111000000000100",
			6582 => "1111111110100000011101",
			6583 => "0000000110100000011101",
			6584 => "0000100110111100001000",
			6585 => "0000000000111000000100",
			6586 => "0000001110100000011101",
			6587 => "0000000110100000011101",
			6588 => "0010101100011100001000",
			6589 => "0011001000111100000100",
			6590 => "0000000110100000011101",
			6591 => "0000000110100000011101",
			6592 => "0010001101010000000100",
			6593 => "0000000110100000011101",
			6594 => "0000000110100000011101",
			6595 => "0011111111010100011000",
			6596 => "0011001010111000010000",
			6597 => "0010100011101000001100",
			6598 => "0001111001001000001000",
			6599 => "0000010111101000000100",
			6600 => "0000000110100000011101",
			6601 => "0000000110100000011101",
			6602 => "0000000110100000011101",
			6603 => "0000000110100000011101",
			6604 => "0001111000011000000100",
			6605 => "0000000110100000011101",
			6606 => "0000000110100000011101",
			6607 => "0001110001101000011000",
			6608 => "0001111001001000001100",
			6609 => "0011000100011000001000",
			6610 => "0011000100001000000100",
			6611 => "0000000110100000011101",
			6612 => "0000000110100000011101",
			6613 => "0000000110100000011101",
			6614 => "0011111010000100000100",
			6615 => "0000000110100000011101",
			6616 => "0001110110100100000100",
			6617 => "0000000110100000011101",
			6618 => "0000000110100000011101",
			6619 => "0011000111001000000100",
			6620 => "0000000110100000011101",
			6621 => "0011011110000100000100",
			6622 => "0000000110100000011101",
			6623 => "0000000110100000011101",
			6624 => "0000110110111000011000",
			6625 => "0000010100110100001100",
			6626 => "0001110101100100001000",
			6627 => "0010011010100100000100",
			6628 => "1111111110100000011101",
			6629 => "0000000110100000011101",
			6630 => "0000000110100000011101",
			6631 => "0001111000011000000100",
			6632 => "0000000110100000011101",
			6633 => "0001111111011100000100",
			6634 => "0000000110100000011101",
			6635 => "0000000110100000011101",
			6636 => "0011011100010100001100",
			6637 => "0011000100011000000100",
			6638 => "0000000110100000011101",
			6639 => "0011111000011100000100",
			6640 => "0000000110100000011101",
			6641 => "0000000110100000011101",
			6642 => "0011100010110000011000",
			6643 => "0001101000010000001100",
			6644 => "0011001111011100000100",
			6645 => "0000000110100000011101",
			6646 => "0001111011011100000100",
			6647 => "0000000110100000011101",
			6648 => "0000000110100000011101",
			6649 => "0010101000010100000100",
			6650 => "0000000110100000011101",
			6651 => "0001011100010000000100",
			6652 => "1111111110100000011101",
			6653 => "0000000110100000011101",
			6654 => "0011011101101100001100",
			6655 => "0000011101111100000100",
			6656 => "0000000110100000011101",
			6657 => "0000101101001000000100",
			6658 => "0000000110100000011101",
			6659 => "0000000110100000011101",
			6660 => "0011000101110100000100",
			6661 => "0000000110100000011101",
			6662 => "0000000110100000011101",
			6663 => "0001011010111100010100",
			6664 => "0000101100000000000100",
			6665 => "1111111110100100001001",
			6666 => "0001000000101100000100",
			6667 => "0000000110100100001001",
			6668 => "0000100000010000001000",
			6669 => "0000000100000000000100",
			6670 => "0000000110100100001001",
			6671 => "0000000110100100001001",
			6672 => "0000000110100100001001",
			6673 => "0011011101101101100000",
			6674 => "0001000011001100111100",
			6675 => "0000010101011100011100",
			6676 => "0000101100000000010000",
			6677 => "0000000010011000001000",
			6678 => "0000010111100100000100",
			6679 => "1111111110100100001001",
			6680 => "0000000110100100001001",
			6681 => "0011001001110000000100",
			6682 => "0000000110100100001001",
			6683 => "1111111110100100001001",
			6684 => "0010000111000100001000",
			6685 => "0010101010110000000100",
			6686 => "1111111110100100001001",
			6687 => "0000000110100100001001",
			6688 => "1111111110100100001001",
			6689 => "0001010111100000010000",
			6690 => "0011000100011000001000",
			6691 => "0000100000010000000100",
			6692 => "0000000110100100001001",
			6693 => "0000000110100100001001",
			6694 => "0010111011011100000100",
			6695 => "0000001110100100001001",
			6696 => "0000000110100100001001",
			6697 => "0000010100110100001000",
			6698 => "0000010101011100000100",
			6699 => "0000001110100100001001",
			6700 => "0000000110100100001001",
			6701 => "0001110110110100000100",
			6702 => "0000000110100100001001",
			6703 => "0000000110100100001001",
			6704 => "0011000000101000001000",
			6705 => "0001101011001100000100",
			6706 => "0000000110100100001001",
			6707 => "0000001110100100001001",
			6708 => "0011100011100000001100",
			6709 => "0001111101100000001000",
			6710 => "0001000010100100000100",
			6711 => "0000000110100100001001",
			6712 => "0000001110100100001001",
			6713 => "1111111110100100001001",
			6714 => "0011001100110000001000",
			6715 => "0001011010111000000100",
			6716 => "0000000110100100001001",
			6717 => "0000001110100100001001",
			6718 => "0000101000000100000100",
			6719 => "1111111110100100001001",
			6720 => "0000000110100100001001",
			6721 => "1111111110100100001001",
			6722 => "0010011011111101010000",
			6723 => "0001111000111000100000",
			6724 => "0001101101011000000100",
			6725 => "1111111110101001111101",
			6726 => "0000111001110100010000",
			6727 => "0001111000111000001100",
			6728 => "0010111000111100000100",
			6729 => "0000000110101001111101",
			6730 => "0001101001100100000100",
			6731 => "0000000110101001111101",
			6732 => "0000001110101001111101",
			6733 => "0000000110101001111101",
			6734 => "0000101111010100001000",
			6735 => "0001111000111100000100",
			6736 => "0000000110101001111101",
			6737 => "0000001110101001111101",
			6738 => "0000000110101001111101",
			6739 => "0001000010010000100000",
			6740 => "0011110010000000011000",
			6741 => "0001100100111100010000",
			6742 => "0000101100000000001000",
			6743 => "0011001001110000000100",
			6744 => "0000000110101001111101",
			6745 => "1111111110101001111101",
			6746 => "0011011001001000000100",
			6747 => "1111111110101001111101",
			6748 => "0000000110101001111101",
			6749 => "0001100100111100000100",
			6750 => "0000001110101001111101",
			6751 => "0000000110101001111101",
			6752 => "0001101000010000000100",
			6753 => "1111111110101001111101",
			6754 => "0000000110101001111101",
			6755 => "0011000011011100001100",
			6756 => "0001101001100100000100",
			6757 => "0000000110101001111101",
			6758 => "0001000000000100000100",
			6759 => "0000001110101001111101",
			6760 => "0000000110101001111101",
			6761 => "0000000110101001111101",
			6762 => "0011111111100100110000",
			6763 => "0010111011011100101100",
			6764 => "0010110000011100011000",
			6765 => "0010000101000100001100",
			6766 => "0000110101110100000100",
			6767 => "0000000110101001111101",
			6768 => "0011110000010000000100",
			6769 => "1111111110101001111101",
			6770 => "0000000110101001111101",
			6771 => "0011110000010000001000",
			6772 => "0001010001101000000100",
			6773 => "0000000110101001111101",
			6774 => "0000000110101001111101",
			6775 => "0000001110101001111101",
			6776 => "0001111001001000000100",
			6777 => "0000000110101001111101",
			6778 => "0001110110100100001000",
			6779 => "0000101000001100000100",
			6780 => "0000001110101001111101",
			6781 => "0000000110101001111101",
			6782 => "0001110110100100000100",
			6783 => "0000000110101001111101",
			6784 => "0000000110101001111101",
			6785 => "0000000110101001111101",
			6786 => "0010010100111100001100",
			6787 => "0001111100101000000100",
			6788 => "0000000110101001111101",
			6789 => "0000000010111100000100",
			6790 => "0000000110101001111101",
			6791 => "1111111110101001111101",
			6792 => "0001011110101000010000",
			6793 => "0000000001110100000100",
			6794 => "0000000110101001111101",
			6795 => "0011111110000000001000",
			6796 => "0010011010100000000100",
			6797 => "0000001110101001111101",
			6798 => "0000000110101001111101",
			6799 => "0000000110101001111101",
			6800 => "0001010010011100010000",
			6801 => "0000110110111000001000",
			6802 => "0001001101001000000100",
			6803 => "0000000110101001111101",
			6804 => "1111111110101001111101",
			6805 => "0011110011001100000100",
			6806 => "0000001110101001111101",
			6807 => "0000000110101001111101",
			6808 => "0010111011110100001000",
			6809 => "0010110101110100000100",
			6810 => "0000000110101001111101",
			6811 => "0000001110101001111101",
			6812 => "0011001001110100000100",
			6813 => "1111111110101001111101",
			6814 => "0000000110101001111101",
			6815 => "0001101011001101011000",
			6816 => "0000010101011100110000",
			6817 => "0001101011001100011100",
			6818 => "0001101001011000001000",
			6819 => "0011001100110000000100",
			6820 => "1111111110110000011001",
			6821 => "0000010110110000011001",
			6822 => "0000111010001100000100",
			6823 => "1111111110110000011001",
			6824 => "0011100110100100001000",
			6825 => "0001101101011000000100",
			6826 => "1111111110110000011001",
			6827 => "0000010110110000011001",
			6828 => "0011010100010000000100",
			6829 => "0000000110110000011001",
			6830 => "1111111110110000011001",
			6831 => "0000100010000100010000",
			6832 => "0011101010111000000100",
			6833 => "1111111110110000011001",
			6834 => "0010101010110000001000",
			6835 => "0000000010011000000100",
			6836 => "0000000110110000011001",
			6837 => "1111111110110000011001",
			6838 => "0000010110110000011001",
			6839 => "1111111110110000011001",
			6840 => "0000111100000000001000",
			6841 => "0000010101011100000100",
			6842 => "0000000110110000011001",
			6843 => "1111111110110000011001",
			6844 => "0000001001101000010000",
			6845 => "0001110110100100000100",
			6846 => "0000001110110000011001",
			6847 => "0000010111101000001000",
			6848 => "0010110101100100000100",
			6849 => "0000000110110000011001",
			6850 => "1111111110110000011001",
			6851 => "0000001110110000011001",
			6852 => "0010100011101000001100",
			6853 => "0000011110010100000100",
			6854 => "0000100110110000011001",
			6855 => "0011011001010000000100",
			6856 => "0000010110110000011001",
			6857 => "0000000110110000011001",
			6858 => "1111111110110000011001",
			6859 => "0010110001001001001100",
			6860 => "0010000001010100100100",
			6861 => "0001001000000100011100",
			6862 => "0000000001110100010000",
			6863 => "0001011101000100001000",
			6864 => "0011101111010100000100",
			6865 => "0000000110110000011001",
			6866 => "0000010110110000011001",
			6867 => "0000101000101000000100",
			6868 => "1111111110110000011001",
			6869 => "0000001110110000011001",
			6870 => "0000000010101000001000",
			6871 => "0011100111010100000100",
			6872 => "0000000110110000011001",
			6873 => "0000010110110000011001",
			6874 => "0000001110110000011001",
			6875 => "0001010111111100000100",
			6876 => "1111111110110000011001",
			6877 => "0000000110110000011001",
			6878 => "0001000100001100010000",
			6879 => "0011011110110000000100",
			6880 => "1111111110110000011001",
			6881 => "0001110101100100001000",
			6882 => "0000001010101100000100",
			6883 => "0000000110110000011001",
			6884 => "0000001110110000011001",
			6885 => "0000100110110000011001",
			6886 => "0011001000111000001100",
			6887 => "0001010100001000000100",
			6888 => "1111111110110000011001",
			6889 => "0001001110001000000100",
			6890 => "0000001110110000011001",
			6891 => "0000000110110000011001",
			6892 => "0001101111000000000100",
			6893 => "1111111110110000011001",
			6894 => "0001111100101000000100",
			6895 => "0000001110110000011001",
			6896 => "1111111110110000011001",
			6897 => "0000011111000000100100",
			6898 => "0001110101100100001100",
			6899 => "0000100011001100001000",
			6900 => "0010110000110100000100",
			6901 => "0000001110110000011001",
			6902 => "1111111110110000011001",
			6903 => "0000001110110000011001",
			6904 => "0000010001111000001100",
			6905 => "0010101010110000001000",
			6906 => "0011010111010100000100",
			6907 => "0000001110110000011001",
			6908 => "0001000110110000011001",
			6909 => "1111111110110000011001",
			6910 => "0011011010000100000100",
			6911 => "1111111110110000011001",
			6912 => "0001011110110100000100",
			6913 => "0000100110110000011001",
			6914 => "1111111110110000011001",
			6915 => "0000100011110100000100",
			6916 => "1111111110110000011001",
			6917 => "0000001110110000011001",
			6918 => "0011101110101101101100",
			6919 => "0010111110001101001000",
			6920 => "0011011001001000110000",
			6921 => "0001000011001100010100",
			6922 => "0000101100010100001000",
			6923 => "0000110100000100000100",
			6924 => "0000000110110111011101",
			6925 => "0000000110110111011101",
			6926 => "0010001001101000000100",
			6927 => "0000000110110111011101",
			6928 => "0000000011010000000100",
			6929 => "1111111110110111011101",
			6930 => "0000000110110111011101",
			6931 => "0000111001110100001100",
			6932 => "0010100001010100000100",
			6933 => "1111111110110111011101",
			6934 => "0010111001110000000100",
			6935 => "0000000110110111011101",
			6936 => "0000000110110111011101",
			6937 => "0011000100000000001000",
			6938 => "0011011110110000000100",
			6939 => "0000000110110111011101",
			6940 => "0000000110110111011101",
			6941 => "0010001010101100000100",
			6942 => "0000000110110111011101",
			6943 => "0000000110110111011101",
			6944 => "0000000011010000001000",
			6945 => "0001101011001100000100",
			6946 => "0000000110110111011101",
			6947 => "0000001110110111011101",
			6948 => "0011100100000100001000",
			6949 => "0000110100000100000100",
			6950 => "0000000110110111011101",
			6951 => "0000001110110111011101",
			6952 => "0001100100111100000100",
			6953 => "1111111110110111011101",
			6954 => "0000000110110111011101",
			6955 => "0000000011010000010000",
			6956 => "0011000100000000000100",
			6957 => "0000000110110111011101",
			6958 => "0000110001001000001000",
			6959 => "0001001000101000000100",
			6960 => "0000000110110111011101",
			6961 => "1111111110110111011101",
			6962 => "0000000110110111011101",
			6963 => "0011010001101000001000",
			6964 => "0000110010001000000100",
			6965 => "0000000110110111011101",
			6966 => "0000001110110111011101",
			6967 => "0010100110011100000100",
			6968 => "1111111110110111011101",
			6969 => "0000110010110100000100",
			6970 => "0000000110110111011101",
			6971 => "0000000110110111011101",
			6972 => "0001001000001001000000",
			6973 => "0001100100111100100000",
			6974 => "0011000000001100001000",
			6975 => "0001010001101000000100",
			6976 => "0000000110110111011101",
			6977 => "1111111110110111011101",
			6978 => "0010011010100100001100",
			6979 => "0010000101000100001000",
			6980 => "0010010101010000000100",
			6981 => "0000000110110111011101",
			6982 => "0000000110110111011101",
			6983 => "0000001110110111011101",
			6984 => "0001000110111000000100",
			6985 => "0000000110110111011101",
			6986 => "0010011010100100000100",
			6987 => "0000000110110111011101",
			6988 => "0000000110110111011101",
			6989 => "0011010111111100000100",
			6990 => "0000001110110111011101",
			6991 => "0011111000110100001100",
			6992 => "0000100011000000000100",
			6993 => "0000000110110111011101",
			6994 => "0010110100010000000100",
			6995 => "0000000110110111011101",
			6996 => "0000000110110111011101",
			6997 => "0010111110101100001000",
			6998 => "0010010011101000000100",
			6999 => "0000001110110111011101",
			7000 => "0000000110110111011101",
			7001 => "0010010011101000000100",
			7002 => "0000000110110111011101",
			7003 => "0000000110110111011101",
			7004 => "0010001011010100011100",
			7005 => "0000110010010100001100",
			7006 => "0001100100111100000100",
			7007 => "0000000110110111011101",
			7008 => "0011100110111000000100",
			7009 => "1111111110110111011101",
			7010 => "0000000110110111011101",
			7011 => "0001011110010000001000",
			7012 => "0000001101010000000100",
			7013 => "0000000110110111011101",
			7014 => "0000000110110111011101",
			7015 => "0010010100101100000100",
			7016 => "0000000110110111011101",
			7017 => "0000000110110111011101",
			7018 => "0011000011011100000100",
			7019 => "0000000110110111011101",
			7020 => "0011000000001100001000",
			7021 => "0001000010111000000100",
			7022 => "0000000110110111011101",
			7023 => "0000001110110111011101",
			7024 => "0011100011010100001000",
			7025 => "0010001111001000000100",
			7026 => "0000000110110111011101",
			7027 => "0000000110110111011101",
			7028 => "0000001100001000000100",
			7029 => "0000001110110111011101",
			7030 => "0000000110110111011101",
			7031 => "0010110011011100010100",
			7032 => "0000100111011000000100",
			7033 => "1111111110111100010001",
			7034 => "0000100000010000001100",
			7035 => "0010011101101000001000",
			7036 => "0010011100110100000100",
			7037 => "0000000110111100010001",
			7038 => "0000000110111100010001",
			7039 => "0000000110111100010001",
			7040 => "0000000110111100010001",
			7041 => "0001111000111000100100",
			7042 => "0011110101001000010100",
			7043 => "0000101100010100000100",
			7044 => "0000000110111100010001",
			7045 => "0011001000111000001100",
			7046 => "0010110011011100000100",
			7047 => "0000000110111100010001",
			7048 => "0010100001010000000100",
			7049 => "0000000110111100010001",
			7050 => "0000001110111100010001",
			7051 => "0000000110111100010001",
			7052 => "0000101111010100001100",
			7053 => "0000110000011100000100",
			7054 => "0000000110111100010001",
			7055 => "0000000010011000000100",
			7056 => "0000000110111100010001",
			7057 => "0000001110111100010001",
			7058 => "1111111110111100010001",
			7059 => "0010010111101001000000",
			7060 => "0000100010000000100000",
			7061 => "0000100011001000010000",
			7062 => "0010011011111100001000",
			7063 => "0010101010100000000100",
			7064 => "0000000110111100010001",
			7065 => "0000000110111100010001",
			7066 => "0001011000011000000100",
			7067 => "0000000110111100010001",
			7068 => "0000000110111100010001",
			7069 => "0001111001110000001000",
			7070 => "0000111001110100000100",
			7071 => "0000000110111100010001",
			7072 => "0000001110111100010001",
			7073 => "0001010111010000000100",
			7074 => "0000000110111100010001",
			7075 => "0000000110111100010001",
			7076 => "0001011001001000010000",
			7077 => "0011011001001000001000",
			7078 => "0001001110111000000100",
			7079 => "1111111110111100010001",
			7080 => "0000000110111100010001",
			7081 => "0000000010111100000100",
			7082 => "1111111110111100010001",
			7083 => "0000000110111100010001",
			7084 => "0000101010000100001000",
			7085 => "0011010110100100000100",
			7086 => "0000000110111100010001",
			7087 => "1111111110111100010001",
			7088 => "0011001001110000000100",
			7089 => "0000000110111100010001",
			7090 => "0000000110111100010001",
			7091 => "0001011010011100001000",
			7092 => "0011100010011100000100",
			7093 => "0000001110111100010001",
			7094 => "0000000110111100010001",
			7095 => "0000111001011100001100",
			7096 => "0000101101000100001000",
			7097 => "0011110101110100000100",
			7098 => "0000000110111100010001",
			7099 => "0000000110111100010001",
			7100 => "1111111110111100010001",
			7101 => "0001111100101000001000",
			7102 => "0000000011111100000100",
			7103 => "0000000110111100010001",
			7104 => "0000001110111100010001",
			7105 => "0001110111001000000100",
			7106 => "1111111110111100010001",
			7107 => "0000000110111100010001",
			7108 => "0001101001100101010000",
			7109 => "0001010111001000000100",
			7110 => "1111111111000001101101",
			7111 => "0000011001111000010000",
			7112 => "0011110001000000001100",
			7113 => "0010000111000100000100",
			7114 => "0000000111000001101101",
			7115 => "0000111001110100000100",
			7116 => "0000000111000001101101",
			7117 => "0000001111000001101101",
			7118 => "0000000111000001101101",
			7119 => "0010001010110000011100",
			7120 => "0001001011101100010000",
			7121 => "0011011111010000001000",
			7122 => "0000001011010100000100",
			7123 => "0000000111000001101101",
			7124 => "0000000111000001101101",
			7125 => "0011010100101000000100",
			7126 => "1111111111000001101101",
			7127 => "0000000111000001101101",
			7128 => "0001101101011000000100",
			7129 => "0000000111000001101101",
			7130 => "0000111111010100000100",
			7131 => "0000000111000001101101",
			7132 => "0000001111000001101101",
			7133 => "0011110101110000010000",
			7134 => "0011101010001100001000",
			7135 => "0010011101011100000100",
			7136 => "0000000111000001101101",
			7137 => "0000000111000001101101",
			7138 => "0001000110111000000100",
			7139 => "0000000111000001101101",
			7140 => "0000000111000001101101",
			7141 => "0011001010111000001000",
			7142 => "0011000100000000000100",
			7143 => "0000000111000001101101",
			7144 => "1111111111000001101101",
			7145 => "0011010010011100000100",
			7146 => "0000000111000001101101",
			7147 => "0000000111000001101101",
			7148 => "0011010110100100110000",
			7149 => "0010111100101100100100",
			7150 => "0011011001001000011100",
			7151 => "0010110101101100010000",
			7152 => "0010011111001100001000",
			7153 => "0010111000111000000100",
			7154 => "0000000111000001101101",
			7155 => "0000001111000001101101",
			7156 => "0000000000110000000100",
			7157 => "0000000111000001101101",
			7158 => "1111111111000001101101",
			7159 => "0011011000000000001000",
			7160 => "0001010100011000000100",
			7161 => "0000000111000001101101",
			7162 => "1111111111000001101101",
			7163 => "0000000111000001101101",
			7164 => "0000000010111100000100",
			7165 => "0000000111000001101101",
			7166 => "0000001111000001101101",
			7167 => "0000000010011000000100",
			7168 => "0000000111000001101101",
			7169 => "0011111110000100000100",
			7170 => "0000000111000001101101",
			7171 => "0000001111000001101101",
			7172 => "0010011011111100010000",
			7173 => "0010101100011100000100",
			7174 => "1111111111000001101101",
			7175 => "0011011000011000001000",
			7176 => "0000110101110100000100",
			7177 => "0000000111000001101101",
			7178 => "0000000111000001101101",
			7179 => "0000000111000001101101",
			7180 => "0001010001101000001000",
			7181 => "0001101111000000000100",
			7182 => "0000000111000001101101",
			7183 => "0000001111000001101101",
			7184 => "0011101110101000001000",
			7185 => "0001101001100100000100",
			7186 => "0000000111000001101101",
			7187 => "1111111111000001101101",
			7188 => "0011000110000100001000",
			7189 => "0010001111001000000100",
			7190 => "0000000111000001101101",
			7191 => "0000001111000001101101",
			7192 => "0001001000001000000100",
			7193 => "0000000111000001101101",
			7194 => "0000000111000001101101",
			7195 => "0010110011011100010000",
			7196 => "0000100111011000000100",
			7197 => "1111111111000110110001",
			7198 => "0011010001111100000100",
			7199 => "1111111111000110110001",
			7200 => "0011011101010100000100",
			7201 => "0000000111000110110001",
			7202 => "0000000111000110110001",
			7203 => "0001000011000001000000",
			7204 => "0000100111010100100000",
			7205 => "0011111010000100011100",
			7206 => "0011111111010100001100",
			7207 => "0010101001000100001000",
			7208 => "0011011111010000000100",
			7209 => "0000000111000110110001",
			7210 => "1111111111000110110001",
			7211 => "0000001111000110110001",
			7212 => "0000101111010100001000",
			7213 => "0000111010000100000100",
			7214 => "0000001111000110110001",
			7215 => "0000000111000110110001",
			7216 => "0011001011000000000100",
			7217 => "0000000111000110110001",
			7218 => "0000000111000110110001",
			7219 => "1111111111000110110001",
			7220 => "0011100111010100001100",
			7221 => "0011111000001100000100",
			7222 => "0000000111000110110001",
			7223 => "0001110001101000000100",
			7224 => "0000001111000110110001",
			7225 => "0000010111000110110001",
			7226 => "0000100110101100001100",
			7227 => "0001110001101000000100",
			7228 => "1111111111000110110001",
			7229 => "0000010001111000000100",
			7230 => "0000000111000110110001",
			7231 => "0000000111000110110001",
			7232 => "0010100011101000000100",
			7233 => "0000001111000110110001",
			7234 => "0000000111000110110001",
			7235 => "0011001000111100100100",
			7236 => "0000001111000100001100",
			7237 => "0000001111000100001000",
			7238 => "0010001001101000000100",
			7239 => "0000000111000110110001",
			7240 => "0000000111000110110001",
			7241 => "1111110111000110110001",
			7242 => "0001001011100000010000",
			7243 => "0000110001101000001000",
			7244 => "0011000000101000000100",
			7245 => "0000000111000110110001",
			7246 => "1111111111000110110001",
			7247 => "0000100010000100000100",
			7248 => "0000001111000110110001",
			7249 => "0000000111000110110001",
			7250 => "0001111101100000000100",
			7251 => "0000001111000110110001",
			7252 => "0000000111000110110001",
			7253 => "0000110010000000011100",
			7254 => "0010000110001000010000",
			7255 => "0000001000101100001000",
			7256 => "0010101000100100000100",
			7257 => "0000000111000110110001",
			7258 => "0000001111000110110001",
			7259 => "0000000010111100000100",
			7260 => "1111111111000110110001",
			7261 => "0000000111000110110001",
			7262 => "0001001100001100000100",
			7263 => "0000001111000110110001",
			7264 => "0011001100110000000100",
			7265 => "0000000111000110110001",
			7266 => "1111111111000110110001",
			7267 => "0001110001111100000100",
			7268 => "0000001111000110110001",
			7269 => "0000001111000100001000",
			7270 => "0000000111000100000100",
			7271 => "0000000111000110110001",
			7272 => "0000000111000110110001",
			7273 => "0010001001101000000100",
			7274 => "1111110111000110110001",
			7275 => "0000000111000110110001",
			7276 => "0001010111100010001000",
			7277 => "0001111110110001001100",
			7278 => "0010000110001000011000",
			7279 => "0011000100000000001000",
			7280 => "0001101011001100000100",
			7281 => "0000000111001101011101",
			7282 => "0000000111001101011101",
			7283 => "0011011000000000000100",
			7284 => "0000000111001101011101",
			7285 => "0010001001000100000100",
			7286 => "0000000111001101011101",
			7287 => "0001101000010000000100",
			7288 => "0000000111001101011101",
			7289 => "0000000111001101011101",
			7290 => "0000111011011100011100",
			7291 => "0011111111010000010000",
			7292 => "0000111001110100001000",
			7293 => "0011110110100000000100",
			7294 => "0000000111001101011101",
			7295 => "0000000111001101011101",
			7296 => "0000010110101000000100",
			7297 => "0000000111001101011101",
			7298 => "0000000111001101011101",
			7299 => "0001111000111000000100",
			7300 => "0000000111001101011101",
			7301 => "0001101111000000000100",
			7302 => "1111111111001101011101",
			7303 => "0000000111001101011101",
			7304 => "0011111001011100001000",
			7305 => "0001010110100100000100",
			7306 => "0000001111001101011101",
			7307 => "0000000111001101011101",
			7308 => "0001100100111100001000",
			7309 => "0000101100000000000100",
			7310 => "0000000111001101011101",
			7311 => "0000000111001101011101",
			7312 => "0000100101000000000100",
			7313 => "0000000111001101011101",
			7314 => "0000000111001101011101",
			7315 => "0011110110111100010100",
			7316 => "0011001010111000010000",
			7317 => "0000101110110100001100",
			7318 => "0011010111100000001000",
			7319 => "0011111110101000000100",
			7320 => "0000000111001101011101",
			7321 => "0000000111001101011101",
			7322 => "0000000111001101011101",
			7323 => "0000000111001101011101",
			7324 => "0000000111001101011101",
			7325 => "0001110001101000011000",
			7326 => "0001111001001000001100",
			7327 => "0011000100011000001000",
			7328 => "0011000100001000000100",
			7329 => "0000000111001101011101",
			7330 => "0000000111001101011101",
			7331 => "0000000111001101011101",
			7332 => "0011111010000100000100",
			7333 => "0000000111001101011101",
			7334 => "0001110110100100000100",
			7335 => "0000000111001101011101",
			7336 => "0000000111001101011101",
			7337 => "0011111010000100000100",
			7338 => "0000000111001101011101",
			7339 => "0010110101100100000100",
			7340 => "0000000111001101011101",
			7341 => "0010110010001000000100",
			7342 => "0000000111001101011101",
			7343 => "0000000111001101011101",
			7344 => "0000110110111000011000",
			7345 => "0000010100110100001100",
			7346 => "0001110101100100001000",
			7347 => "0010011010100100000100",
			7348 => "1111111111001101011101",
			7349 => "0000000111001101011101",
			7350 => "0000000111001101011101",
			7351 => "0001111000011000000100",
			7352 => "0000000111001101011101",
			7353 => "0001111111011100000100",
			7354 => "0000000111001101011101",
			7355 => "0000000111001101011101",
			7356 => "0001010111111100001000",
			7357 => "0000010100110100000100",
			7358 => "0000000111001101011101",
			7359 => "0000000111001101011101",
			7360 => "0000110010111000011000",
			7361 => "0001101000010000001100",
			7362 => "0011001111011100000100",
			7363 => "0000000111001101011101",
			7364 => "0001111011011100000100",
			7365 => "0000000111001101011101",
			7366 => "0000000111001101011101",
			7367 => "0010101000010100000100",
			7368 => "0000000111001101011101",
			7369 => "0001011100010000000100",
			7370 => "1111111111001101011101",
			7371 => "0000000111001101011101",
			7372 => "0011000111010000001100",
			7373 => "0000011010011000000100",
			7374 => "0000000111001101011101",
			7375 => "0010001001101000000100",
			7376 => "0000000111001101011101",
			7377 => "0000000111001101011101",
			7378 => "0001110000110100000100",
			7379 => "0000000111001101011101",
			7380 => "0001100100101100000100",
			7381 => "0000000111001101011101",
			7382 => "0000000111001101011101",
			7383 => "0011101110101101101100",
			7384 => "0011111001010000110100",
			7385 => "0000111010001100100100",
			7386 => "0000101110110100001100",
			7387 => "0001001110111000001000",
			7388 => "0011010111010000000100",
			7389 => "1111111111010100110001",
			7390 => "0000000111010100110001",
			7391 => "0000000111010100110001",
			7392 => "0001101011001100001100",
			7393 => "0000010010001100001000",
			7394 => "0001011010111000000100",
			7395 => "0000000111010100110001",
			7396 => "0000000111010100110001",
			7397 => "0000000111010100110001",
			7398 => "0000111001110100001000",
			7399 => "0001011110110000000100",
			7400 => "0000000111010100110001",
			7401 => "0000000111010100110001",
			7402 => "0000001111010100110001",
			7403 => "0000101100010100000100",
			7404 => "0000000111010100110001",
			7405 => "0011000100000000000100",
			7406 => "0000000111010100110001",
			7407 => "0000001100001000000100",
			7408 => "0000001111010100110001",
			7409 => "0000000111010100110001",
			7410 => "0001000010111000011000",
			7411 => "0011000100000000001000",
			7412 => "0001101001100100000100",
			7413 => "0000000111010100110001",
			7414 => "0000000111010100110001",
			7415 => "0000010111100100001000",
			7416 => "0001101011001100000100",
			7417 => "0000000111010100110001",
			7418 => "1111111111010100110001",
			7419 => "0001101001100100000100",
			7420 => "0000000111010100110001",
			7421 => "0000000111010100110001",
			7422 => "0000000000110000001100",
			7423 => "0001101001100100000100",
			7424 => "0000000111010100110001",
			7425 => "0001010110100100000100",
			7426 => "0000001111010100110001",
			7427 => "0000000111010100110001",
			7428 => "0001101111000000001000",
			7429 => "0010100001010100000100",
			7430 => "1111111111010100110001",
			7431 => "0000000111010100110001",
			7432 => "0010101100000100001000",
			7433 => "0000110010001000000100",
			7434 => "0000000111010100110001",
			7435 => "0000000111010100110001",
			7436 => "0000000111010100110001",
			7437 => "0001010111100000110100",
			7438 => "0000110010000100011100",
			7439 => "0011111111100100011000",
			7440 => "0010100001010000001100",
			7441 => "0000100111011000001000",
			7442 => "0011100101001000000100",
			7443 => "0000000111010100110001",
			7444 => "0000000111010100110001",
			7445 => "1111111111010100110001",
			7446 => "0010010001111000000100",
			7447 => "0000000111010100110001",
			7448 => "0011100111111100000100",
			7449 => "0000001111010100110001",
			7450 => "0000000111010100110001",
			7451 => "1111111111010100110001",
			7452 => "0010000111000000010100",
			7453 => "0000101000101000010000",
			7454 => "0010010111101100001000",
			7455 => "0011110110111100000100",
			7456 => "0000000111010100110001",
			7457 => "0000000111010100110001",
			7458 => "0000010001111000000100",
			7459 => "0000000111010100110001",
			7460 => "0000000111010100110001",
			7461 => "0000001111010100110001",
			7462 => "0000000111010100110001",
			7463 => "0001010010011100011000",
			7464 => "0001011111010000001100",
			7465 => "0000001010101100000100",
			7466 => "0000000111010100110001",
			7467 => "0001001001001100000100",
			7468 => "0000001111010100110001",
			7469 => "0000000111010100110001",
			7470 => "0010010010101100001000",
			7471 => "0000110110111000000100",
			7472 => "1111111111010100110001",
			7473 => "0000000111010100110001",
			7474 => "0000000111010100110001",
			7475 => "0011101000101000010100",
			7476 => "0011010011001000000100",
			7477 => "0000000111010100110001",
			7478 => "0011000001101000001000",
			7479 => "0000001011010100000100",
			7480 => "0000000111010100110001",
			7481 => "0000001111010100110001",
			7482 => "0000010101011100000100",
			7483 => "0000000111010100110001",
			7484 => "0000000111010100110001",
			7485 => "0001010011001000010000",
			7486 => "0011101011110000001000",
			7487 => "0000110010010100000100",
			7488 => "0000000111010100110001",
			7489 => "1111111111010100110001",
			7490 => "0001011110010000000100",
			7491 => "0000000111010100110001",
			7492 => "0000000111010100110001",
			7493 => "0000110100001100001000",
			7494 => "0000011101011000000100",
			7495 => "0000000111010100110001",
			7496 => "0000000111010100110001",
			7497 => "0011101011100000000100",
			7498 => "0000000111010100110001",
			7499 => "0000000111010100110001",
			7500 => "0010110011011100001000",
			7501 => "0001101001100100000100",
			7502 => "1111111111011001010101",
			7503 => "0000000111011001010101",
			7504 => "0001000011000000110000",
			7505 => "0000110111110000010000",
			7506 => "0010011011111100001000",
			7507 => "0001111101111000000100",
			7508 => "1111111111011001010101",
			7509 => "0000000111011001010101",
			7510 => "0011011010001100000100",
			7511 => "0000000111011001010101",
			7512 => "0000000111011001010101",
			7513 => "0010101000100100011100",
			7514 => "0010110000011100010000",
			7515 => "0011010101110100001000",
			7516 => "0001111100101000000100",
			7517 => "0000000111011001010101",
			7518 => "0000001111011001010101",
			7519 => "0000111100000000000100",
			7520 => "1111111111011001010101",
			7521 => "0000000111011001010101",
			7522 => "0000010101011100000100",
			7523 => "1111111111011001010101",
			7524 => "0001101001100100000100",
			7525 => "0000001111011001010101",
			7526 => "0000000111011001010101",
			7527 => "0000001111011001010101",
			7528 => "0001101001100100111100",
			7529 => "0000010110101000011100",
			7530 => "0000111010011100010000",
			7531 => "0001001111100000001000",
			7532 => "0011101000000000000100",
			7533 => "1111111111011001010101",
			7534 => "0000000111011001010101",
			7535 => "0011000100000000000100",
			7536 => "0000001111011001010101",
			7537 => "1111111111011001010101",
			7538 => "0000101100000000001000",
			7539 => "0000000011010000000100",
			7540 => "0000000111011001010101",
			7541 => "0000001111011001010101",
			7542 => "1111111111011001010101",
			7543 => "0001000011110000010000",
			7544 => "0000000010111100001000",
			7545 => "0011010110100100000100",
			7546 => "1111111111011001010101",
			7547 => "0000000111011001010101",
			7548 => "0001111001110000000100",
			7549 => "0000000111011001010101",
			7550 => "0000001111011001010101",
			7551 => "0010110110000100001000",
			7552 => "0010011001011000000100",
			7553 => "1111111111011001010101",
			7554 => "0000000111011001010101",
			7555 => "0000001101010000000100",
			7556 => "0000000111011001010101",
			7557 => "1111111111011001010101",
			7558 => "0011001000111100001100",
			7559 => "0011000000101000001000",
			7560 => "0000010110101000000100",
			7561 => "0000001111011001010101",
			7562 => "1111111111011001010101",
			7563 => "0000001111011001010101",
			7564 => "0000001001110000010000",
			7565 => "0000011101011000001000",
			7566 => "0010010111101100000100",
			7567 => "0000000111011001010101",
			7568 => "0000000111011001010101",
			7569 => "0000000000111000000100",
			7570 => "1111111111011001010101",
			7571 => "0000000111011001010101",
			7572 => "1111111111011001010101",
			7573 => "0011101110101101100000",
			7574 => "0010111110001101000100",
			7575 => "0011011001001000101100",
			7576 => "0001010100011000011100",
			7577 => "0011011110110000001100",
			7578 => "0001000001101100000100",
			7579 => "1111111111100000101001",
			7580 => "0010111001110000000100",
			7581 => "0000000111100000101001",
			7582 => "0000000111100000101001",
			7583 => "0011111001010000001000",
			7584 => "0001111000111000000100",
			7585 => "0000000111100000101001",
			7586 => "0000000111100000101001",
			7587 => "0001111000111000000100",
			7588 => "0000000111100000101001",
			7589 => "0000000111100000101001",
			7590 => "0000100111011000001000",
			7591 => "0011000100000000000100",
			7592 => "0000000111100000101001",
			7593 => "1111111111100000101001",
			7594 => "0000101111010100000100",
			7595 => "0000000111100000101001",
			7596 => "0000000111100000101001",
			7597 => "0000000011010000001000",
			7598 => "0011111111010000000100",
			7599 => "0000000111100000101001",
			7600 => "0000001111100000101001",
			7601 => "0011100100000100001000",
			7602 => "0001111101100000000100",
			7603 => "0000001111100000101001",
			7604 => "0000000111100000101001",
			7605 => "0001111101100000000100",
			7606 => "1111111111100000101001",
			7607 => "0000000111100000101001",
			7608 => "0000010110101000001000",
			7609 => "0010100110011100000100",
			7610 => "1111111111100000101001",
			7611 => "0000000111100000101001",
			7612 => "0001011001001000001000",
			7613 => "0011110100101000000100",
			7614 => "0000000111100000101001",
			7615 => "0000001111100000101001",
			7616 => "0010010101011100000100",
			7617 => "0000000111100000101001",
			7618 => "0001001000001100000100",
			7619 => "0000000111100000101001",
			7620 => "1111111111100000101001",
			7621 => "0001001000001001001100",
			7622 => "0011001110001100010000",
			7623 => "0010110100001000001000",
			7624 => "0010100110011000000100",
			7625 => "0000000111100000101001",
			7626 => "0000000111100000101001",
			7627 => "0000011001011000000100",
			7628 => "1111111111100000101001",
			7629 => "0000000111100000101001",
			7630 => "0010000101000100100000",
			7631 => "0010100010101100010000",
			7632 => "0000100111011000001000",
			7633 => "0011001010111000000100",
			7634 => "0000000111100000101001",
			7635 => "0000000111100000101001",
			7636 => "0000010001000100000100",
			7637 => "0000000111100000101001",
			7638 => "0000001111100000101001",
			7639 => "0001001011101100001000",
			7640 => "0001010010110100000100",
			7641 => "0000000111100000101001",
			7642 => "1111111111100000101001",
			7643 => "0001000011000000000100",
			7644 => "0000000111100000101001",
			7645 => "0000000111100000101001",
			7646 => "0001110110110100001100",
			7647 => "0000011101011000001000",
			7648 => "0000000001110100000100",
			7649 => "0000000111100000101001",
			7650 => "0000000111100000101001",
			7651 => "0000000111100000101001",
			7652 => "0011110110001100001000",
			7653 => "0010010011101000000100",
			7654 => "0000000111100000101001",
			7655 => "0000000111100000101001",
			7656 => "0011101110100100000100",
			7657 => "0000000111100000101001",
			7658 => "0000000111100000101001",
			7659 => "0010001011010100101000",
			7660 => "0000001111000100011100",
			7661 => "0010010100101100001100",
			7662 => "0010100110011000001000",
			7663 => "0001000010111000000100",
			7664 => "0000000111100000101001",
			7665 => "0000001111100000101001",
			7666 => "0000000111100000101001",
			7667 => "0000001101010000001000",
			7668 => "0011001011000000000100",
			7669 => "0000000111100000101001",
			7670 => "0000000111100000101001",
			7671 => "0010010000001000000100",
			7672 => "0000000111100000101001",
			7673 => "0000000111100000101001",
			7674 => "0011101011110000000100",
			7675 => "1111111111100000101001",
			7676 => "0001110001011000000100",
			7677 => "0000000111100000101001",
			7678 => "0000000111100000101001",
			7679 => "0011000011011100000100",
			7680 => "0000000111100000101001",
			7681 => "0001110100001000000100",
			7682 => "0000001111100000101001",
			7683 => "0011100011010100001000",
			7684 => "0010100110011100000100",
			7685 => "0000000111100000101001",
			7686 => "0000000111100000101001",
			7687 => "0000001100001000000100",
			7688 => "0000001111100000101001",
			7689 => "0000000111100000101001",
			7690 => "0000111001110100100000",
			7691 => "0000010111100100011100",
			7692 => "0000101001100000000100",
			7693 => "1111111111100101111101",
			7694 => "0011000100000000001100",
			7695 => "0010001000110000000100",
			7696 => "1111111111100101111101",
			7697 => "0001010000001100000100",
			7698 => "1111111111100101111101",
			7699 => "0000001111100101111101",
			7700 => "0001111000111000001000",
			7701 => "0001111000111000000100",
			7702 => "1111111111100101111101",
			7703 => "0000000111100101111101",
			7704 => "1111111111100101111101",
			7705 => "0000001111100101111101",
			7706 => "0011001000011001100100",
			7707 => "0010000001110000110000",
			7708 => "0000001100000100010000",
			7709 => "0010010101010000001100",
			7710 => "0011010100010000001000",
			7711 => "0000011011101000000100",
			7712 => "1111111111100101111101",
			7713 => "0000010111100101111101",
			7714 => "1111111111100101111101",
			7715 => "0000001111100101111101",
			7716 => "0001010111100000010000",
			7717 => "0010110100000100001000",
			7718 => "0011100110111100000100",
			7719 => "0000000111100101111101",
			7720 => "0000001111100101111101",
			7721 => "0001111001001000000100",
			7722 => "0000000111100101111101",
			7723 => "0000001111100101111101",
			7724 => "0010011001111100001000",
			7725 => "0001010101110000000100",
			7726 => "1111111111100101111101",
			7727 => "0000001111100101111101",
			7728 => "0000001010101100000100",
			7729 => "1111111111100101111101",
			7730 => "0000000111100101111101",
			7731 => "0010010111101100100000",
			7732 => "0011001000111000010000",
			7733 => "0001010111001000001000",
			7734 => "0001000011110100000100",
			7735 => "1111111111100101111101",
			7736 => "0000000111100101111101",
			7737 => "0000010111100100000100",
			7738 => "0000001111100101111101",
			7739 => "0000001111100101111101",
			7740 => "0000111110010000001000",
			7741 => "0001110101101100000100",
			7742 => "0000000111100101111101",
			7743 => "1111111111100101111101",
			7744 => "0011000110000100000100",
			7745 => "0000001111100101111101",
			7746 => "0000000111100101111101",
			7747 => "0010111011110100001000",
			7748 => "0001001110111000000100",
			7749 => "0000001111100101111101",
			7750 => "0000000111100101111101",
			7751 => "0011101011110000000100",
			7752 => "1111111111100101111101",
			7753 => "0011001001110100000100",
			7754 => "1111111111100101111101",
			7755 => "0000001111100101111101",
			7756 => "0010011000010100100000",
			7757 => "0010001011010100011100",
			7758 => "0011011010000100010000",
			7759 => "0000010001111000001000",
			7760 => "0000010001111000000100",
			7761 => "0000000111100101111101",
			7762 => "0000011111100101111101",
			7763 => "0011010110111100000100",
			7764 => "1111111111100101111101",
			7765 => "0000000111100101111101",
			7766 => "0011101000011100000100",
			7767 => "0000010111100101111101",
			7768 => "0001110111110000000100",
			7769 => "1111111111100101111101",
			7770 => "0000010111100101111101",
			7771 => "1111111111100101111101",
			7772 => "0000000010111100000100",
			7773 => "0000000111100101111101",
			7774 => "0000001111100101111101",
			7775 => "0001101011001101001100",
			7776 => "0010011000010000100100",
			7777 => "0001101101011000011000",
			7778 => "0001101001011000001000",
			7779 => "0001010110100100000100",
			7780 => "1111111111101100111001",
			7781 => "0000001111101100111001",
			7782 => "0001000101110000001100",
			7783 => "0010101001111100000100",
			7784 => "1111111111101100111001",
			7785 => "0001011110101100000100",
			7786 => "0000010111101100111001",
			7787 => "0000000111101100111001",
			7788 => "1111111111101100111001",
			7789 => "0000111010001100000100",
			7790 => "1111111111101100111001",
			7791 => "0000100010000100000100",
			7792 => "0000010111101100111001",
			7793 => "1111111111101100111001",
			7794 => "0001111001001000001000",
			7795 => "0011100111111100000100",
			7796 => "0000001111101100111001",
			7797 => "1111111111101100111001",
			7798 => "0001110110100100010000",
			7799 => "0011100010000000000100",
			7800 => "1111111111101100111001",
			7801 => "0000010001000100000100",
			7802 => "0000000111101100111001",
			7803 => "0001110110100100000100",
			7804 => "0000010111101100111001",
			7805 => "0000001111101100111001",
			7806 => "0000001001101000001000",
			7807 => "0010110101100100000100",
			7808 => "0000001111101100111001",
			7809 => "1111111111101100111001",
			7810 => "0011001001110100000100",
			7811 => "0000010111101100111001",
			7812 => "1111111111101100111001",
			7813 => "0011001000011001101000",
			7814 => "0001101000010000111100",
			7815 => "0001111101100000011100",
			7816 => "0000010110101000010000",
			7817 => "0011110111111100001000",
			7818 => "0001010111001000000100",
			7819 => "0000000111101100111001",
			7820 => "0000001111101100111001",
			7821 => "0000000000111000000100",
			7822 => "1111111111101100111001",
			7823 => "0000000111101100111001",
			7824 => "0001101001100100000100",
			7825 => "0000000111101100111001",
			7826 => "0000010111100100000100",
			7827 => "0000001111101100111001",
			7828 => "0000001111101100111001",
			7829 => "0000111100010000010000",
			7830 => "0010111101111000001000",
			7831 => "0000010111100100000100",
			7832 => "1111111111101100111001",
			7833 => "0000001111101100111001",
			7834 => "0001101000010000000100",
			7835 => "1111111111101100111001",
			7836 => "0000000111101100111001",
			7837 => "0001010001000000001000",
			7838 => "0010100111110100000100",
			7839 => "0000000111101100111001",
			7840 => "0000001111101100111001",
			7841 => "0010011001111100000100",
			7842 => "0000001111101100111001",
			7843 => "1111111111101100111001",
			7844 => "0010111011110100011000",
			7845 => "0001000011010100001100",
			7846 => "0010101001000100000100",
			7847 => "0000000111101100111001",
			7848 => "0010011010011000000100",
			7849 => "0000001111101100111001",
			7850 => "0000001111101100111001",
			7851 => "0001110001111100000100",
			7852 => "0000001111101100111001",
			7853 => "0001101001111100000100",
			7854 => "1111111111101100111001",
			7855 => "0000000111101100111001",
			7856 => "0011110010110000001000",
			7857 => "0011001000011000000100",
			7858 => "1111111111101100111001",
			7859 => "0000000111101100111001",
			7860 => "0010100001010000000100",
			7861 => "1111111111101100111001",
			7862 => "0001001011100000000100",
			7863 => "0000001111101100111001",
			7864 => "0000001111101100111001",
			7865 => "0010011000010100100100",
			7866 => "0010101010110000100000",
			7867 => "0010011010100000010000",
			7868 => "0001110100010000001000",
			7869 => "0001101000010000000100",
			7870 => "0000001111101100111001",
			7871 => "1111111111101100111001",
			7872 => "0010100001010000000100",
			7873 => "0000011111101100111001",
			7874 => "0000001111101100111001",
			7875 => "0010110110100000001000",
			7876 => "0011001000011000000100",
			7877 => "0000000111101100111001",
			7878 => "1111111111101100111001",
			7879 => "0001000110001100000100",
			7880 => "0000011111101100111001",
			7881 => "1111111111101100111001",
			7882 => "1111111111101100111001",
			7883 => "0000000010111100000100",
			7884 => "1111111111101100111001",
			7885 => "0000001111101100111001",
			7886 => "0000010110101001001100",
			7887 => "0001000010111000010100",
			7888 => "0010010101011100010000",
			7889 => "0011111110000100000100",
			7890 => "0000000111110011111101",
			7891 => "0001111101100000001000",
			7892 => "0001111000111000000100",
			7893 => "0000000111110011111101",
			7894 => "1111111111110011111101",
			7895 => "0000000111110011111101",
			7896 => "0000000111110011111101",
			7897 => "0011000100000000100000",
			7898 => "0001011010111000010100",
			7899 => "0001101001100100001100",
			7900 => "0011000100010100000100",
			7901 => "0000000111110011111101",
			7902 => "0001000111011100000100",
			7903 => "0000000111110011111101",
			7904 => "0000000111110011111101",
			7905 => "0010110011011100000100",
			7906 => "0000000111110011111101",
			7907 => "0000000111110011111101",
			7908 => "0011010100011000000100",
			7909 => "0000000111110011111101",
			7910 => "0001111001110000000100",
			7911 => "0000001111110011111101",
			7912 => "0000000111110011111101",
			7913 => "0001000010010000010000",
			7914 => "0000010110101000001100",
			7915 => "0010011011101000000100",
			7916 => "0000000111110011111101",
			7917 => "0001111000111000000100",
			7918 => "0000000111110011111101",
			7919 => "1111111111110011111101",
			7920 => "0000000111110011111101",
			7921 => "0001101111000000000100",
			7922 => "0000000111110011111101",
			7923 => "0000000111110011111101",
			7924 => "0000100110111100110100",
			7925 => "0001101001100100100100",
			7926 => "0001001100001100100000",
			7927 => "0001110110100100010000",
			7928 => "0011001110001100001000",
			7929 => "0001111101100000000100",
			7930 => "0000000111110011111101",
			7931 => "0000000111110011111101",
			7932 => "0000010111101000000100",
			7933 => "0000000111110011111101",
			7934 => "0000000111110011111101",
			7935 => "0010001000100100001000",
			7936 => "0000010000111100000100",
			7937 => "0000000111110011111101",
			7938 => "0000000111110011111101",
			7939 => "0000011110010100000100",
			7940 => "0000000111110011111101",
			7941 => "0000000111110011111101",
			7942 => "0000000111110011111101",
			7943 => "0001001011110000001000",
			7944 => "0001001111101000000100",
			7945 => "0000000111110011111101",
			7946 => "0000000111110011111101",
			7947 => "0010100001010000000100",
			7948 => "0000000111110011111101",
			7949 => "0000001111110011111101",
			7950 => "0011111011110000110100",
			7951 => "0000100010010100100000",
			7952 => "0011110000010000010000",
			7953 => "0001101111000000001000",
			7954 => "0011001011000000000100",
			7955 => "1111111111110011111101",
			7956 => "0000000111110011111101",
			7957 => "0010111101111000000100",
			7958 => "0000000111110011111101",
			7959 => "0000000111110011111101",
			7960 => "0001110110100100001000",
			7961 => "0011011110000100000100",
			7962 => "0000000111110011111101",
			7963 => "0000000111110011111101",
			7964 => "0000010101011100000100",
			7965 => "0000000111110011111101",
			7966 => "0000000111110011111101",
			7967 => "0001100101010000001100",
			7968 => "0001101111000000000100",
			7969 => "0000000111110011111101",
			7970 => "0001001000110100000100",
			7971 => "0000000111110011111101",
			7972 => "1111111111110011111101",
			7973 => "0001110110100100000100",
			7974 => "0000000111110011111101",
			7975 => "0000000111110011111101",
			7976 => "0010111011110100010000",
			7977 => "0000010111101000000100",
			7978 => "0000000111110011111101",
			7979 => "0011110011001100001000",
			7980 => "0010010010101100000100",
			7981 => "0000001111110011111101",
			7982 => "0000000111110011111101",
			7983 => "0000000111110011111101",
			7984 => "0001101001111100010000",
			7985 => "0001110000011100001000",
			7986 => "0010010011101000000100",
			7987 => "0000000111110011111101",
			7988 => "0000000111110011111101",
			7989 => "0000011100011000000100",
			7990 => "0000000111110011111101",
			7991 => "0000000111110011111101",
			7992 => "0000110011011000001000",
			7993 => "0001110010001000000100",
			7994 => "0000000111110011111101",
			7995 => "0000000111110011111101",
			7996 => "0000100011111000000100",
			7997 => "0000000111110011111101",
			7998 => "0000000111110011111101",
			7999 => "0001101101011001000100",
			8000 => "0010010101010000100000",
			8001 => "0000010111100100001100",
			8002 => "0000111010001100000100",
			8003 => "1111111111111011001011",
			8004 => "0011100110100100000100",
			8005 => "0000000111111011001011",
			8006 => "1111111111111011001011",
			8007 => "0001110011100000010000",
			8008 => "0011001110001100000100",
			8009 => "1111111111111011001011",
			8010 => "0000000001110000000100",
			8011 => "1111111111111011001011",
			8012 => "0000001101010000000100",
			8013 => "0000001111111011001011",
			8014 => "0000000111111011001011",
			8015 => "1111111111111011001011",
			8016 => "0010101010100100001000",
			8017 => "0010010101010000000100",
			8018 => "0000000111111011001011",
			8019 => "0000010111111011001011",
			8020 => "0001111001001000000100",
			8021 => "1111111111111011001011",
			8022 => "0010000001010000010000",
			8023 => "0000011011111100001000",
			8024 => "0000010001000100000100",
			8025 => "0000000111111011001011",
			8026 => "1111111111111011001011",
			8027 => "0010000110011000000100",
			8028 => "0000000111111011001011",
			8029 => "0000010111111011001011",
			8030 => "0010100011101000000100",
			8031 => "1111111111111011001011",
			8032 => "0000000111111011001011",
			8033 => "0011001000011001110100",
			8034 => "0001101001100100111000",
			8035 => "0000101001100000011000",
			8036 => "0000110100000100001100",
			8037 => "0001001001001100000100",
			8038 => "1111111111111011001011",
			8039 => "0000111010111100000100",
			8040 => "1111111111111011001011",
			8041 => "0000001111111011001011",
			8042 => "0000000011111100001000",
			8043 => "0001101011001100000100",
			8044 => "0000000111111011001011",
			8045 => "0000001111111011001011",
			8046 => "0000001111111011001011",
			8047 => "0000111100010000010000",
			8048 => "0011111110010000001000",
			8049 => "0010001001101000000100",
			8050 => "1111110111111011001011",
			8051 => "0000000111111011001011",
			8052 => "0000101100010000000100",
			8053 => "0000000111111011001011",
			8054 => "1111111111111011001011",
			8055 => "0011111010000100001000",
			8056 => "0000010001111000000100",
			8057 => "0000010111111011001011",
			8058 => "1111111111111011001011",
			8059 => "0000001011010100000100",
			8060 => "1111111111111011001011",
			8061 => "0000000111111011001011",
			8062 => "0010000001110000100000",
			8063 => "0001111000011000010000",
			8064 => "0001001000000100001000",
			8065 => "0000000111000100000100",
			8066 => "1111111111111011001011",
			8067 => "0000001111111011001011",
			8068 => "0000111100111000000100",
			8069 => "1111111111111011001011",
			8070 => "0000001111111011001011",
			8071 => "0011010110010000001000",
			8072 => "0011010100101000000100",
			8073 => "0000000111111011001011",
			8074 => "1111111111111011001011",
			8075 => "0001110001011000000100",
			8076 => "0000001111111011001011",
			8077 => "0000000111111011001011",
			8078 => "0011100001011100010000",
			8079 => "0001111101100000001000",
			8080 => "0000010110101000000100",
			8081 => "0000001111111011001011",
			8082 => "0000001111111011001011",
			8083 => "0010001001101000000100",
			8084 => "0000001111111011001011",
			8085 => "0000000111111011001011",
			8086 => "0010000111000100001000",
			8087 => "0001101000010000000100",
			8088 => "0000010111111011001011",
			8089 => "0000001111111011001011",
			8090 => "0000000111111011001011",
			8091 => "0011010110111100010100",
			8092 => "0000010001111000010000",
			8093 => "0000010001111000001100",
			8094 => "0011011100000000000100",
			8095 => "1111111111111011001011",
			8096 => "0000001101010000000100",
			8097 => "0000001111111011001011",
			8098 => "0000000111111011001011",
			8099 => "0000010111111011001011",
			8100 => "1111111111111011001011",
			8101 => "0000000111000000001100",
			8102 => "0000111100001100001000",
			8103 => "0011000111010000000100",
			8104 => "0000000111111011001011",
			8105 => "0000001111111011001011",
			8106 => "0000100111111011001011",
			8107 => "0000001011000100001100",
			8108 => "0001001010110100000100",
			8109 => "1111111111111011001011",
			8110 => "0010100001010000000100",
			8111 => "0000001111111011001011",
			8112 => "0000000111111011001011",
			8113 => "1111111111111011001011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2750, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5367, initial_addr_3'length));
	end generate gen_rom_9;

	gen_rom_10: if SELECT_ROM = 10 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0001001111100100000100",
			21 => "0000000000000001100101",
			22 => "0000011100011000000100",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0001100100111100000100",
			26 => "0000000000000001111001",
			27 => "0001101001111100000100",
			28 => "0000000000000001111001",
			29 => "0000000000000001111001",
			30 => "0000010100110100001000",
			31 => "0010010111101100000100",
			32 => "0000000000000010001101",
			33 => "0000000000000010001101",
			34 => "0000000000000010001101",
			35 => "0000011100011000001000",
			36 => "0000000001110000000100",
			37 => "0000000000000010100001",
			38 => "0000000000000010100001",
			39 => "0000000000000010100001",
			40 => "0010011010100100001000",
			41 => "0011101011110000000100",
			42 => "0000000000000010110101",
			43 => "0000000000000010110101",
			44 => "0000000000000010110101",
			45 => "0000000010101000001100",
			46 => "0000000010101000000100",
			47 => "0000000000000011010001",
			48 => "0010000101000100000100",
			49 => "0000000000000011010001",
			50 => "0000000000000011010001",
			51 => "0000000000000011010001",
			52 => "0011101100001100001100",
			53 => "0000011100011000001000",
			54 => "0011101011111000000100",
			55 => "0000000000000011101101",
			56 => "0000000000000011101101",
			57 => "0000000000000011101101",
			58 => "0000000000000011101101",
			59 => "0001001000011100000100",
			60 => "0000000000000100001001",
			61 => "0001001011100000001000",
			62 => "0010010100101100000100",
			63 => "0000000000000100001001",
			64 => "0000000000000100001001",
			65 => "0000000000000100001001",
			66 => "0010011010100000000100",
			67 => "0000000000000100100101",
			68 => "0001010111011000001000",
			69 => "0010010011101000000100",
			70 => "0000000000000100100101",
			71 => "0000000000000100100101",
			72 => "0000000000000100100101",
			73 => "0000000010101000001100",
			74 => "0010011010100100000100",
			75 => "0000000000000101010001",
			76 => "0011110011000000000100",
			77 => "0000000000000101010001",
			78 => "0000000000000101010001",
			79 => "0011110101000000001000",
			80 => "0000001010101100000100",
			81 => "0000000000000101010001",
			82 => "0000000000000101010001",
			83 => "0000000000000101010001",
			84 => "0010111011011100000100",
			85 => "0000000000000101110101",
			86 => "0001101001111100001100",
			87 => "0001100100111100000100",
			88 => "0000000000000101110101",
			89 => "0010110110100000000100",
			90 => "0000000000000101110101",
			91 => "0000000000000101110101",
			92 => "0000000000000101110101",
			93 => "0001110110100100001000",
			94 => "0011001101010100000100",
			95 => "0000000000000110100001",
			96 => "0000000000000110100001",
			97 => "0000010111101000000100",
			98 => "0000000000000110100001",
			99 => "0010011010100100001000",
			100 => "0010010100101100000100",
			101 => "0000000000000110100001",
			102 => "0000000000000110100001",
			103 => "0000000000000110100001",
			104 => "0001110001101000010000",
			105 => "0000000010101000001100",
			106 => "0001111000000000000100",
			107 => "0000000000000111001101",
			108 => "0000000001010100000100",
			109 => "0000000000000111001101",
			110 => "0000000000000111001101",
			111 => "0000000000000111001101",
			112 => "0001110111010000000100",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0000001010101100001100",
			116 => "0010011010100100000100",
			117 => "0000000000001000001001",
			118 => "0000110001011100000100",
			119 => "0000000000001000001001",
			120 => "0000000000001000001001",
			121 => "0011101110000000001000",
			122 => "0000011100011000000100",
			123 => "0000000000001000001001",
			124 => "0000000000001000001001",
			125 => "0011011111100100001000",
			126 => "0001110111010000000100",
			127 => "0000000000001000001001",
			128 => "0000000000001000001001",
			129 => "0000000000001000001001",
			130 => "0001001011110000010100",
			131 => "0000111101101100010000",
			132 => "0011001000000000001100",
			133 => "0011001101010100000100",
			134 => "0000000000001000111101",
			135 => "0001000010000100000100",
			136 => "0000000000001000111101",
			137 => "0000000000001000111101",
			138 => "0000000000001000111101",
			139 => "0000000000001000111101",
			140 => "0000111000000100000100",
			141 => "0000000000001000111101",
			142 => "0000000000001000111101",
			143 => "0010111011011100000100",
			144 => "0000000000001001101001",
			145 => "0001101001111100010000",
			146 => "0001100100111100000100",
			147 => "0000000000001001101001",
			148 => "0001010111011000001000",
			149 => "0001011100100100000100",
			150 => "0000000000001001101001",
			151 => "0000000000001001101001",
			152 => "0000000000001001101001",
			153 => "0000000000001001101001",
			154 => "0010010111101100010000",
			155 => "0001110111010000001100",
			156 => "0011101000101000001000",
			157 => "0001100100110100000100",
			158 => "0000000000001010101101",
			159 => "0000000000001010101101",
			160 => "0000000000001010101101",
			161 => "0000000000001010101101",
			162 => "0010010011101000010000",
			163 => "0001101001111100001100",
			164 => "0010100011101000000100",
			165 => "0000000000001010101101",
			166 => "0011100110010000000100",
			167 => "0000000000001010101101",
			168 => "0000000000001010101101",
			169 => "0000000000001010101101",
			170 => "0000000000001010101101",
			171 => "0001110110100100010100",
			172 => "0011001101010100000100",
			173 => "0000000000001011110001",
			174 => "0010000001010100001100",
			175 => "0010001000010100000100",
			176 => "0000000000001011110001",
			177 => "0001110011100000000100",
			178 => "0000000000001011110001",
			179 => "0000000000001011110001",
			180 => "0000000000001011110001",
			181 => "0000010111101000000100",
			182 => "0000000000001011110001",
			183 => "0010011010100100001000",
			184 => "0010010100101100000100",
			185 => "0000000000001011110001",
			186 => "0000000000001011110001",
			187 => "0000000000001011110001",
			188 => "0001001011110000010100",
			189 => "0011101011101100010000",
			190 => "0010001010110000000100",
			191 => "0000000000001101000101",
			192 => "0011100110010000000100",
			193 => "0000000000001101000101",
			194 => "0000000010101000000100",
			195 => "0000000000001101000101",
			196 => "0000000000001101000101",
			197 => "0000000000001101000101",
			198 => "0011101110000000001100",
			199 => "0010011001111100000100",
			200 => "0000000000001101000101",
			201 => "0010010010101100000100",
			202 => "0000000000001101000101",
			203 => "0000000000001101000101",
			204 => "0001011111010100001000",
			205 => "0010111011110100000100",
			206 => "0000000000001101000101",
			207 => "0000000000001101000101",
			208 => "0000000000001101000101",
			209 => "0001001011110000011000",
			210 => "0011101011101100010100",
			211 => "0011011110101100000100",
			212 => "0000000000001110000001",
			213 => "0011011100010100001100",
			214 => "0010001000100100000100",
			215 => "0000000000001110000001",
			216 => "0000001010101100000100",
			217 => "0000000000001110000001",
			218 => "0000000000001110000001",
			219 => "0000000000001110000001",
			220 => "0000000000001110000001",
			221 => "0011100010010100000100",
			222 => "0000000000001110000001",
			223 => "0000000000001110000001",
			224 => "0011011111100100011000",
			225 => "0001101011001100000100",
			226 => "0000000000001110110101",
			227 => "0001101001111100010000",
			228 => "0011001101010100000100",
			229 => "0000000000001110110101",
			230 => "0000000000111000001000",
			231 => "0010100011101000000100",
			232 => "0000000000001110110101",
			233 => "0000000000001110110101",
			234 => "0000000000001110110101",
			235 => "0000000000001110110101",
			236 => "0000000000001110110101",
			237 => "0001011001010000000100",
			238 => "0000000000001111101001",
			239 => "0011011011111000010100",
			240 => "0010010010101100010000",
			241 => "0000000010101000000100",
			242 => "0000000000001111101001",
			243 => "0011101100111000000100",
			244 => "0000000000001111101001",
			245 => "0001000111011100000100",
			246 => "0000000000001111101001",
			247 => "0000000000001111101001",
			248 => "0000000000001111101001",
			249 => "0000000000001111101001",
			250 => "0011011110010000011000",
			251 => "0010010000001000000100",
			252 => "0000000000010000110101",
			253 => "0011101111101000010000",
			254 => "0001111000011000001100",
			255 => "0010101001000100001000",
			256 => "0010001010110000000100",
			257 => "0000000000010000110101",
			258 => "0000000000010000110101",
			259 => "0000000000010000110101",
			260 => "0000000000010000110101",
			261 => "0000000000010000110101",
			262 => "0000010111101000000100",
			263 => "0000000000010000110101",
			264 => "0000100011110100001000",
			265 => "0010010100101100000100",
			266 => "0000000000010000110101",
			267 => "0000000000010000110101",
			268 => "0000000000010000110101",
			269 => "0000000001110100010100",
			270 => "0000111111100100010000",
			271 => "0001100100110100000100",
			272 => "0000000000010010010001",
			273 => "0011011110010000001000",
			274 => "0011001101010100000100",
			275 => "0000000000010010010001",
			276 => "0000000000010010010001",
			277 => "0000000000010010010001",
			278 => "0000000000010010010001",
			279 => "0001111111011100001100",
			280 => "0010011010100100001000",
			281 => "0000011100011000000100",
			282 => "0000000000010010010001",
			283 => "0000000000010010010001",
			284 => "0000000000010010010001",
			285 => "0000010100110100001100",
			286 => "0011011111100100001000",
			287 => "0010011111000000000100",
			288 => "0000000000010010010001",
			289 => "0000000000010010010001",
			290 => "0000000000010010010001",
			291 => "0000000000010010010001",
			292 => "0010010111101100001100",
			293 => "0001101000010000001000",
			294 => "0011001000011000000100",
			295 => "0000000000010011011101",
			296 => "0000000000010011011101",
			297 => "0000000000010011011101",
			298 => "0011011110010000011000",
			299 => "0011101111101000010100",
			300 => "0001011100100100000100",
			301 => "0000000000010011011101",
			302 => "0000000111000100000100",
			303 => "0000000000010011011101",
			304 => "0011001001001000001000",
			305 => "0010000001110000000100",
			306 => "0000000000010011011101",
			307 => "0000000000010011011101",
			308 => "0000000000010011011101",
			309 => "0000000000010011011101",
			310 => "0000000000010011011101",
			311 => "0001100100111100001100",
			312 => "0001001011101100000100",
			313 => "0000000000010100101001",
			314 => "0000011010011000000100",
			315 => "0000000000010100101001",
			316 => "0000000000010100101001",
			317 => "0011000001011000011000",
			318 => "0000000010101000000100",
			319 => "0000000000010100101001",
			320 => "0000000010111100010000",
			321 => "0010110010001000000100",
			322 => "0000000000010100101001",
			323 => "0011000100011000000100",
			324 => "0000000000010100101001",
			325 => "0011010111010100000100",
			326 => "0000000000010100101001",
			327 => "0000000000010100101001",
			328 => "0000000000010100101001",
			329 => "0000000000010100101001",
			330 => "0000001010101100011100",
			331 => "0010110101110100011000",
			332 => "0010010000001000000100",
			333 => "0000000000010101101101",
			334 => "0001111000011000010000",
			335 => "0000101000101000001100",
			336 => "0001011100100100000100",
			337 => "0000000000010101101101",
			338 => "0000000111000100000100",
			339 => "0000000000010101101101",
			340 => "0000000000010101101101",
			341 => "0000000000010101101101",
			342 => "0000000000010101101101",
			343 => "0000000000010101101101",
			344 => "0001101000010000000100",
			345 => "0000000000010101101101",
			346 => "0000000000010101101101",
			347 => "0010010111101100010100",
			348 => "0001101000010000001000",
			349 => "0000000111000100000100",
			350 => "0000000000010111011001",
			351 => "0000000000010111011001",
			352 => "0001000000010100001000",
			353 => "0001010111111100000100",
			354 => "0000000000010111011001",
			355 => "0000000000010111011001",
			356 => "0000000000010111011001",
			357 => "0010110001000000100000",
			358 => "0000010100110100010000",
			359 => "0010100011101000000100",
			360 => "0000000000010111011001",
			361 => "0000001011010100000100",
			362 => "0000000000010111011001",
			363 => "0011100110010000000100",
			364 => "0000000000010111011001",
			365 => "0000000000010111011001",
			366 => "0000000111000000001000",
			367 => "0000000001110100000100",
			368 => "0000000000010111011001",
			369 => "0000000000010111011001",
			370 => "0000000010011000000100",
			371 => "0000000000010111011001",
			372 => "0000000000010111011001",
			373 => "0000000000010111011001",
			374 => "0001100100111100000100",
			375 => "0000000000011000010101",
			376 => "0011011111100100011000",
			377 => "0001101001111100010100",
			378 => "0011010111111100000100",
			379 => "0000000000011000010101",
			380 => "0010100110011100001100",
			381 => "0010110110110100000100",
			382 => "0000000000011000010101",
			383 => "0010101000010100000100",
			384 => "0000000000011000010101",
			385 => "0000000000011000010101",
			386 => "0000000000011000010101",
			387 => "0000000000011000010101",
			388 => "0000000000011000010101",
			389 => "0010111011011100001000",
			390 => "0001001011101100000100",
			391 => "0000000000011001110001",
			392 => "0000000000011001110001",
			393 => "0010110010110100011000",
			394 => "0001101001100100000100",
			395 => "0000000000011001110001",
			396 => "0010001011010100010000",
			397 => "0010010011101000001100",
			398 => "0011000100011000000100",
			399 => "0000000000011001110001",
			400 => "0001110001101000000100",
			401 => "0000000000011001110001",
			402 => "0000000000011001110001",
			403 => "0000000000011001110001",
			404 => "0000000000011001110001",
			405 => "0010001111001000001100",
			406 => "0011001111011100000100",
			407 => "0000000000011001110001",
			408 => "0001110010001000000100",
			409 => "0000000000011001110001",
			410 => "0000000000011001110001",
			411 => "0000000000011001110001",
			412 => "0000000010101000010100",
			413 => "0010010000001000000100",
			414 => "0000000000011011010101",
			415 => "0001111000011000001100",
			416 => "0000101000101000001000",
			417 => "0011100110010000000100",
			418 => "0000000000011011010101",
			419 => "0000000000011011010101",
			420 => "0000000000011011010101",
			421 => "0000000000011011010101",
			422 => "0001111111011100000100",
			423 => "0000000000011011010101",
			424 => "0001101000010000001000",
			425 => "0001110101100100000100",
			426 => "0000000000011011010101",
			427 => "0000000000011011010101",
			428 => "0011011011111000010000",
			429 => "0010010010101100001100",
			430 => "0001101001111100001000",
			431 => "0011101100111000000100",
			432 => "0000000000011011010101",
			433 => "0000000000011011010101",
			434 => "0000000000011011010101",
			435 => "0000000000011011010101",
			436 => "0000000000011011010101",
			437 => "0010010111101100011100",
			438 => "0011100001011100001100",
			439 => "0001001100010000000100",
			440 => "0000000000011101100001",
			441 => "0011001111011100000100",
			442 => "0000000000011101100001",
			443 => "0000000000011101100001",
			444 => "0001010010000100001100",
			445 => "0001110111010000000100",
			446 => "0000000000011101100001",
			447 => "0001000011010100000100",
			448 => "0000000000011101100001",
			449 => "0000000000011101100001",
			450 => "0000000000011101100001",
			451 => "0011101011101100010000",
			452 => "0001011100100100000100",
			453 => "0000000000011101100001",
			454 => "0000001010101100001000",
			455 => "0000000111000100000100",
			456 => "0000000000011101100001",
			457 => "0000000000011101100001",
			458 => "0000000000011101100001",
			459 => "0000000111000000001000",
			460 => "0010000001010100000100",
			461 => "0000000000011101100001",
			462 => "0000000000011101100001",
			463 => "0001010110111100010000",
			464 => "0001101000010000000100",
			465 => "0000000000011101100001",
			466 => "0001011001010000000100",
			467 => "0000000000011101100001",
			468 => "0001101001111100000100",
			469 => "0000000000011101100001",
			470 => "0000000000011101100001",
			471 => "0000000000011101100001",
			472 => "0001001000110100011100",
			473 => "0011011100010100011000",
			474 => "0001101000010000010100",
			475 => "0000000010101000010000",
			476 => "0001100100110100000100",
			477 => "0000000000011111010101",
			478 => "0000101000101000001000",
			479 => "0001110011100000000100",
			480 => "0000000000011111010101",
			481 => "0000000000011111010101",
			482 => "0000000000011111010101",
			483 => "0000000000011111010101",
			484 => "0000000000011111010101",
			485 => "0000000000011111010101",
			486 => "0001010111111100001000",
			487 => "0000001010101100000100",
			488 => "0000000000011111010101",
			489 => "0000000000011111010101",
			490 => "0001110100010000010000",
			491 => "0001001110111000001100",
			492 => "0010101000010100000100",
			493 => "0000000000011111010101",
			494 => "0010010010101100000100",
			495 => "0000000000011111010101",
			496 => "0000000000011111010101",
			497 => "0000000000011111010101",
			498 => "0011101110100100000100",
			499 => "0000000000011111010101",
			500 => "0000000000011111010101",
			501 => "0000001101010000101100",
			502 => "0011000100011000010000",
			503 => "0001001000100000001100",
			504 => "0010100011101000000100",
			505 => "0000000000100001011001",
			506 => "0011100110010000000100",
			507 => "0000000000100001011001",
			508 => "0000000000100001011001",
			509 => "0000000000100001011001",
			510 => "0001110101100100010100",
			511 => "0010010011101000010000",
			512 => "0011010101110000000100",
			513 => "0000000000100001011001",
			514 => "0010001100000100001000",
			515 => "0010101000100100000100",
			516 => "0000000000100001011001",
			517 => "0000000000100001011001",
			518 => "0000000000100001011001",
			519 => "0000000000100001011001",
			520 => "0010000001110000000100",
			521 => "0000000000100001011001",
			522 => "0000000000100001011001",
			523 => "0011101100001100000100",
			524 => "0000000000100001011001",
			525 => "0010011010100100010000",
			526 => "0011011011111000001100",
			527 => "0000110101000000000100",
			528 => "0000000000100001011001",
			529 => "0000001000111100000100",
			530 => "0000000000100001011001",
			531 => "0000000000100001011001",
			532 => "0000000000100001011001",
			533 => "0000000000100001011001",
			534 => "0001001000110100011100",
			535 => "0011011100010100011000",
			536 => "0001101000010000010100",
			537 => "0001100100110100000100",
			538 => "0000000000100011010101",
			539 => "0000101000101000001100",
			540 => "0010101000010100001000",
			541 => "0001110011100000000100",
			542 => "0000000000100011010101",
			543 => "0000000000100011010101",
			544 => "0000000000100011010101",
			545 => "0000000000100011010101",
			546 => "0000000000100011010101",
			547 => "0000000000100011010101",
			548 => "0011101000110100001100",
			549 => "0000011110010100000100",
			550 => "0000000000100011010101",
			551 => "0010011001111100000100",
			552 => "0000000000100011010101",
			553 => "0000000000100011010101",
			554 => "0011011111100100010100",
			555 => "0001110111010000000100",
			556 => "0000000000100011010101",
			557 => "0000010001000100000100",
			558 => "0000000000100011010101",
			559 => "0000011100011000001000",
			560 => "0011101000011100000100",
			561 => "0000000000100011010101",
			562 => "0000000000100011010101",
			563 => "0000000000100011010101",
			564 => "0000000000100011010101",
			565 => "0001111000011000100100",
			566 => "0011000100011000001100",
			567 => "0001001000100000000100",
			568 => "0000000000100101100001",
			569 => "0000011100011000000100",
			570 => "0000000000100101100001",
			571 => "0000000000100101100001",
			572 => "0011001000000000010100",
			573 => "0011011110010000010000",
			574 => "0010101001000100001100",
			575 => "0001110110100100000100",
			576 => "0000000000100101100001",
			577 => "0001100100110100000100",
			578 => "0000000000100101100001",
			579 => "0000000000100101100001",
			580 => "0000000000100101100001",
			581 => "0000000000100101100001",
			582 => "0000000000100101100001",
			583 => "0001111111011100000100",
			584 => "0000000000100101100001",
			585 => "0001010110111100011000",
			586 => "0000010100110100010000",
			587 => "0000010101011100000100",
			588 => "0000000000100101100001",
			589 => "0011001001110100000100",
			590 => "0000000000100101100001",
			591 => "0001010101110000000100",
			592 => "0000000000100101100001",
			593 => "0000000000100101100001",
			594 => "0001111111011100000100",
			595 => "0000000000100101100001",
			596 => "0000000000100101100001",
			597 => "0011000100000100000100",
			598 => "0000000000100101100001",
			599 => "0000000000100101100001",
			600 => "0010011010100000101000",
			601 => "0001111111011100001000",
			602 => "0001000110101100000100",
			603 => "0000000000101000001101",
			604 => "1111111000101000001101",
			605 => "0001110010001000010100",
			606 => "0001000011001100010000",
			607 => "0011110000010000000100",
			608 => "0000000000101000001101",
			609 => "0000000110001000000100",
			610 => "0000000000101000001101",
			611 => "0001011100010100000100",
			612 => "0000000000101000001101",
			613 => "0000000000101000001101",
			614 => "0000000000101000001101",
			615 => "0011111000001000001000",
			616 => "0011001111011100000100",
			617 => "0000000000101000001101",
			618 => "0000000000101000001101",
			619 => "0000000000101000001101",
			620 => "0011001001110100011100",
			621 => "0000001000101100011000",
			622 => "0001011100100100001000",
			623 => "0011001010111000000100",
			624 => "0000000000101000001101",
			625 => "0000000000101000001101",
			626 => "0011000100011000000100",
			627 => "0000000000101000001101",
			628 => "0000011101111100000100",
			629 => "0000000000101000001101",
			630 => "0010011010100000000100",
			631 => "0000000000101000001101",
			632 => "0000001000101000001101",
			633 => "0000000000101000001101",
			634 => "0000010100110100001100",
			635 => "0001101000010000000100",
			636 => "0000000000101000001101",
			637 => "0001010111111100000100",
			638 => "0000000000101000001101",
			639 => "0000000000101000001101",
			640 => "0001000110111000000100",
			641 => "0000000000101000001101",
			642 => "0000000000101000001101",
			643 => "0001001000000100100100",
			644 => "0010011010100100011000",
			645 => "0001101001100100010100",
			646 => "0001100100110100000100",
			647 => "0000000000101010110001",
			648 => "0000011101111100001100",
			649 => "0001010101110000001000",
			650 => "0001111000000000000100",
			651 => "0000000000101010110001",
			652 => "0000000000101010110001",
			653 => "0000000000101010110001",
			654 => "0000000000101010110001",
			655 => "0000000000101010110001",
			656 => "0001111111011100001000",
			657 => "0000101000101000000100",
			658 => "0000001000101010110001",
			659 => "0000000000101010110001",
			660 => "0000000000101010110001",
			661 => "0011101100001100011100",
			662 => "0001001010110100011000",
			663 => "0001010111111100001000",
			664 => "0000011100011000000100",
			665 => "0000000000101010110001",
			666 => "0000000000101010110001",
			667 => "0001000110001100000100",
			668 => "0000000000101010110001",
			669 => "0011010111011000001000",
			670 => "0000011100011000000100",
			671 => "0000000000101010110001",
			672 => "0000000000101010110001",
			673 => "0000000000101010110001",
			674 => "1111111000101010110001",
			675 => "0010110001000000010000",
			676 => "0010110000110100000100",
			677 => "0000000000101010110001",
			678 => "0010010010101100001000",
			679 => "0000011011111100000100",
			680 => "0000000000101010110001",
			681 => "0000001000101010110001",
			682 => "0000000000101010110001",
			683 => "0000000000101010110001",
			684 => "0000010101011100011000",
			685 => "0000000111000100010000",
			686 => "0010100011101000001100",
			687 => "0010011011111100001000",
			688 => "0001011111011100000100",
			689 => "1111111000101101010101",
			690 => "0000011000101101010101",
			691 => "1111111000101101010101",
			692 => "0000011000101101010101",
			693 => "0000011001011000000100",
			694 => "1111111000101101010101",
			695 => "1111111000101101010101",
			696 => "0010010010101100110100",
			697 => "0001011001010000011100",
			698 => "0010011010100000001100",
			699 => "0001001111100100001000",
			700 => "0001101011001100000100",
			701 => "1111111000101101010101",
			702 => "0000011000101101010101",
			703 => "1111111000101101010101",
			704 => "0000101111100100000100",
			705 => "0000010000101101010101",
			706 => "0000011100011000001000",
			707 => "0000011100011000000100",
			708 => "1111111000101101010101",
			709 => "0000000000101101010101",
			710 => "0000011000101101010101",
			711 => "0010000101000100001000",
			712 => "0010010101010000000100",
			713 => "0000000000101101010101",
			714 => "1111111000101101010101",
			715 => "0000100010010100000100",
			716 => "0000011000101101010101",
			717 => "0001010111011000001000",
			718 => "0001100100111100000100",
			719 => "1111111000101101010101",
			720 => "0000001000101101010101",
			721 => "1111111000101101010101",
			722 => "0001110001101000000100",
			723 => "0000000000101101010101",
			724 => "1111111000101101010101",
			725 => "0000000010111101000100",
			726 => "0011101000110100110100",
			727 => "0000001000101100101000",
			728 => "0010111011110100011000",
			729 => "0001011001010000001100",
			730 => "0000111111100100001000",
			731 => "0010010000001000000100",
			732 => "0000000000101111101001",
			733 => "0000000000101111101001",
			734 => "0000000000101111101001",
			735 => "0001111000011000000100",
			736 => "0000000000101111101001",
			737 => "0001001111101000000100",
			738 => "0000000000101111101001",
			739 => "0000001000101111101001",
			740 => "0000000111000000001000",
			741 => "0000111111101000000100",
			742 => "0000000000101111101001",
			743 => "0000000000101111101001",
			744 => "0011011110110100000100",
			745 => "0000000000101111101001",
			746 => "0000000000101111101001",
			747 => "0011101110000000001000",
			748 => "0010011010100100000100",
			749 => "0000000000101111101001",
			750 => "0000000000101111101001",
			751 => "0000000000101111101001",
			752 => "0001010111111100000100",
			753 => "0000000000101111101001",
			754 => "0010100110011000000100",
			755 => "0000000000101111101001",
			756 => "0000011010011000000100",
			757 => "0000001000101111101001",
			758 => "0000000000101111101001",
			759 => "0011100010110000000100",
			760 => "1111111000101111101001",
			761 => "0000000000101111101001",
			762 => "0011001101010100000100",
			763 => "1111111000110001101101",
			764 => "0000101000100000100000",
			765 => "0001101011001100001100",
			766 => "0000011011101000001000",
			767 => "0001111001001000000100",
			768 => "0000000000110001101101",
			769 => "0000001000110001101101",
			770 => "1111111000110001101101",
			771 => "0010000101000100010000",
			772 => "0011101011111000001100",
			773 => "0011100110010000000100",
			774 => "0000000000110001101101",
			775 => "0010100011101000000100",
			776 => "0000000000110001101101",
			777 => "0000001000110001101101",
			778 => "0000000000110001101101",
			779 => "0000000000110001101101",
			780 => "0010110010001000000100",
			781 => "1111111000110001101101",
			782 => "0011001000000000001100",
			783 => "0011001011000000000100",
			784 => "0000000000110001101101",
			785 => "0000010100110100000100",
			786 => "0000000000110001101101",
			787 => "0000001000110001101101",
			788 => "0010011010100100001100",
			789 => "0001111111011100000100",
			790 => "1111111000110001101101",
			791 => "0011011111100100000100",
			792 => "0000000000110001101101",
			793 => "1111111000110001101101",
			794 => "1111111000110001101101",
			795 => "0001011001010100000100",
			796 => "1111111000110011001001",
			797 => "0011011111100100101000",
			798 => "0010010010101100100000",
			799 => "0001100100110100000100",
			800 => "1111111000110011001001",
			801 => "0011101100001100010000",
			802 => "0000001101010000001000",
			803 => "0001101000010000000100",
			804 => "0000000000110011001001",
			805 => "0000001000110011001001",
			806 => "0011101000011100000100",
			807 => "1111111000110011001001",
			808 => "0000000000110011001001",
			809 => "0000000000110000001000",
			810 => "0001010011001000000100",
			811 => "0000000000110011001001",
			812 => "0000001000110011001001",
			813 => "0000000000110011001001",
			814 => "0001011110000100000100",
			815 => "0000000000110011001001",
			816 => "1111111000110011001001",
			817 => "1111111000110011001001",
			818 => "0001010110111100111100",
			819 => "0000110011110000110000",
			820 => "0010001100000100101000",
			821 => "0001101000010000011100",
			822 => "0011101011111000001100",
			823 => "0000110000010000000100",
			824 => "0000000000110101000101",
			825 => "0001101111000000000100",
			826 => "0000000000110101000101",
			827 => "0000000000110101000101",
			828 => "0001100100111100001000",
			829 => "0000010001000100000100",
			830 => "0000000000110101000101",
			831 => "0000000000110101000101",
			832 => "0011111000000100000100",
			833 => "0000000000110101000101",
			834 => "0000000000110101000101",
			835 => "0001111000011000000100",
			836 => "0000000000110101000101",
			837 => "0010010010101100000100",
			838 => "0000000000110101000101",
			839 => "0000000000110101000101",
			840 => "0011101000110100000100",
			841 => "0000000000110101000101",
			842 => "0000000000110101000101",
			843 => "0010010010101100001000",
			844 => "0001000001100100000100",
			845 => "0000000000110101000101",
			846 => "0000000000110101000101",
			847 => "0000000000110101000101",
			848 => "0000000000110101000101",
			849 => "0001110110100100001100",
			850 => "0010011010100100000100",
			851 => "1111111000110111001001",
			852 => "0000011100011000000100",
			853 => "0000001000110111001001",
			854 => "0000000000110111001001",
			855 => "0011011111100100110100",
			856 => "0010010010101100101100",
			857 => "0011011001011100010000",
			858 => "0011010110100000000100",
			859 => "0000001000110111001001",
			860 => "0010011010100000000100",
			861 => "1111111000110111001001",
			862 => "0001100100111100000100",
			863 => "0000001000110111001001",
			864 => "1111111000110111001001",
			865 => "0000101110000000010000",
			866 => "0010111010010100001000",
			867 => "0000000110001000000100",
			868 => "1111111000110111001001",
			869 => "0000010000110111001001",
			870 => "0000011011111100000100",
			871 => "0000001000110111001001",
			872 => "1111111000110111001001",
			873 => "0010111011110100000100",
			874 => "1111111000110111001001",
			875 => "0001101000010000000100",
			876 => "1111111000110111001001",
			877 => "0000001000110111001001",
			878 => "0010110110110100000100",
			879 => "0000001000110111001001",
			880 => "1111111000110111001001",
			881 => "1111111000110111001001",
			882 => "0010011010100001000000",
			883 => "0001111111011100011000",
			884 => "0000000110001000010100",
			885 => "0010110100000100010000",
			886 => "0001111000000000000100",
			887 => "0000000000111010100101",
			888 => "0011001101010100000100",
			889 => "0000000000111010100101",
			890 => "0001110110100100000100",
			891 => "0000001000111010100101",
			892 => "0000000000111010100101",
			893 => "0000000000111010100101",
			894 => "1111111000111010100101",
			895 => "0001011110110100011000",
			896 => "0000111110000000010000",
			897 => "0011111000110100001100",
			898 => "0001101001100100000100",
			899 => "0000000000111010100101",
			900 => "0001110101100100000100",
			901 => "0000000000111010100101",
			902 => "0000000000111010100101",
			903 => "0000000000111010100101",
			904 => "0000000000110000000100",
			905 => "0000001000111010100101",
			906 => "0000000000111010100101",
			907 => "0010100001010000000100",
			908 => "1111111000111010100101",
			909 => "0011011000001100001000",
			910 => "0011111111100000000100",
			911 => "0000000000111010100101",
			912 => "0000000000111010100101",
			913 => "0000000000111010100101",
			914 => "0000111101101100010000",
			915 => "0000001010101100001100",
			916 => "0010111011011100001000",
			917 => "0010110000011100000100",
			918 => "0000000000111010100101",
			919 => "0000000000111010100101",
			920 => "0000001000111010100101",
			921 => "0000000000111010100101",
			922 => "0000000010101000000100",
			923 => "0000000000111010100101",
			924 => "0000001101010000010100",
			925 => "0010010010101100001100",
			926 => "0011011010001000000100",
			927 => "0000000000111010100101",
			928 => "0001111011011100000100",
			929 => "0000001000111010100101",
			930 => "0000000000111010100101",
			931 => "0011001000000000000100",
			932 => "0000000000111010100101",
			933 => "0000000000111010100101",
			934 => "0011100011110000000100",
			935 => "0000000000111010100101",
			936 => "0000000000111010100101",
			937 => "0000000010101000101100",
			938 => "0010101000100100100000",
			939 => "0011101011111000011000",
			940 => "0001101011001100001000",
			941 => "0010010000001000000100",
			942 => "0000000000111101110001",
			943 => "0000000000111101110001",
			944 => "0010000101000100001100",
			945 => "0010001100011100000100",
			946 => "0000000000111101110001",
			947 => "0000110111011000000100",
			948 => "0000000000111101110001",
			949 => "0000001000111101110001",
			950 => "0000000000111101110001",
			951 => "0000000010101000000100",
			952 => "0000000000111101110001",
			953 => "0000000000111101110001",
			954 => "0001101000010000001000",
			955 => "0000110001011100000100",
			956 => "0000001000111101110001",
			957 => "0000000000111101110001",
			958 => "0000000000111101110001",
			959 => "0011100001011100000100",
			960 => "1111111000111101110001",
			961 => "0010110110100000100100",
			962 => "0011011100010100010100",
			963 => "0001101000010000001100",
			964 => "0011001011000000000100",
			965 => "0000000000111101110001",
			966 => "0010110100010000000100",
			967 => "0000000000111101110001",
			968 => "0000000000111101110001",
			969 => "0001111000011000000100",
			970 => "0000000000111101110001",
			971 => "0000000000111101110001",
			972 => "0010010010101100001100",
			973 => "0001101000010000000100",
			974 => "0000000000111101110001",
			975 => "0010000110001000000100",
			976 => "0000001000111101110001",
			977 => "0000000000111101110001",
			978 => "0000000000111101110001",
			979 => "0001101001111100001000",
			980 => "0011011111010100000100",
			981 => "0000000000111101110001",
			982 => "0000000000111101110001",
			983 => "0010011010100100001000",
			984 => "0010010100101100000100",
			985 => "0000000000111101110001",
			986 => "0000000000111101110001",
			987 => "0000000000111101110001",
			988 => "0000000010011001001000",
			989 => "0000111000110100110100",
			990 => "0000001000110000101100",
			991 => "0010111011110100011000",
			992 => "0001011001010000001100",
			993 => "0000111111100100001000",
			994 => "0010010000001000000100",
			995 => "0000000001000000001101",
			996 => "0000000001000000001101",
			997 => "0000000001000000001101",
			998 => "0001111000011000000100",
			999 => "0000000001000000001101",
			1000 => "0001001111101000000100",
			1001 => "0000000001000000001101",
			1002 => "0000001001000000001101",
			1003 => "0000000111000000001100",
			1004 => "0000111111101000000100",
			1005 => "0000000001000000001101",
			1006 => "0001001100001100000100",
			1007 => "0000000001000000001101",
			1008 => "0000000001000000001101",
			1009 => "0001010011001000000100",
			1010 => "0000000001000000001101",
			1011 => "0000000001000000001101",
			1012 => "0000111110000000000100",
			1013 => "1111111001000000001101",
			1014 => "0000000001000000001101",
			1015 => "0010100110011000000100",
			1016 => "0000000001000000001101",
			1017 => "0000011100011000001100",
			1018 => "0001000100001100001000",
			1019 => "0000000010011000000100",
			1020 => "0000001001000000001101",
			1021 => "0000000001000000001101",
			1022 => "0000000001000000001101",
			1023 => "0000000001000000001101",
			1024 => "0011100011110000000100",
			1025 => "1111111001000000001101",
			1026 => "0000000001000000001101",
			1027 => "0001001011110000101100",
			1028 => "0001101011001100001000",
			1029 => "0000011101111100000100",
			1030 => "0000000001000011011001",
			1031 => "0000000001000011011001",
			1032 => "0011101011101100011100",
			1033 => "0001011100100100010000",
			1034 => "0000100110111100001000",
			1035 => "0000110010000100000100",
			1036 => "0000000001000011011001",
			1037 => "0000000001000011011001",
			1038 => "0011000111001000000100",
			1039 => "0000000001000011011001",
			1040 => "0000000001000011011001",
			1041 => "0010100011101000000100",
			1042 => "0000000001000011011001",
			1043 => "0000000110001000000100",
			1044 => "0000000001000011011001",
			1045 => "0000001001000011011001",
			1046 => "0011001000000000000100",
			1047 => "0000000001000011011001",
			1048 => "0000000001000011011001",
			1049 => "0011100001011100001000",
			1050 => "0010010010101100000100",
			1051 => "1111111001000011011001",
			1052 => "0000000001000011011001",
			1053 => "0000000111000000001000",
			1054 => "0011101000101000000100",
			1055 => "0000000001000011011001",
			1056 => "0000000001000011011001",
			1057 => "0010110110100000010100",
			1058 => "0010111011110100001000",
			1059 => "0010101001000100000100",
			1060 => "0000000001000011011001",
			1061 => "0000000001000011011001",
			1062 => "0001001110111000001000",
			1063 => "0001101000010000000100",
			1064 => "0000000001000011011001",
			1065 => "0000001001000011011001",
			1066 => "0000000001000011011001",
			1067 => "0001101001111100001100",
			1068 => "0011011111010100000100",
			1069 => "0000000001000011011001",
			1070 => "0001001010110100000100",
			1071 => "0000000001000011011001",
			1072 => "0000000001000011011001",
			1073 => "0000010100110100001000",
			1074 => "0000011110010100000100",
			1075 => "0000000001000011011001",
			1076 => "0000000001000011011001",
			1077 => "0000000001000011011001",
			1078 => "0000010101011100011000",
			1079 => "0000000111000000010000",
			1080 => "0000111000100000001100",
			1081 => "0011001011000000000100",
			1082 => "1111111001000110011101",
			1083 => "0010011101011000000100",
			1084 => "0000011001000110011101",
			1085 => "1111111001000110011101",
			1086 => "0000011001000110011101",
			1087 => "0010011001100100000100",
			1088 => "1111111001000110011101",
			1089 => "1111110001000110011101",
			1090 => "0010010010101101000100",
			1091 => "0001011001010000100000",
			1092 => "0001000110111000011000",
			1093 => "0010011010100000001100",
			1094 => "0010010000001000000100",
			1095 => "1111111001000110011101",
			1096 => "0000010001111000000100",
			1097 => "0000100001000110011101",
			1098 => "0000000001000110011101",
			1099 => "0011101000001100000100",
			1100 => "0000011001000110011101",
			1101 => "0000111011101100000100",
			1102 => "0000001001000110011101",
			1103 => "1111111001000110011101",
			1104 => "0000011100011000000100",
			1105 => "1111111001000110011101",
			1106 => "0000000001000110011101",
			1107 => "0010000001010100010000",
			1108 => "0010010101010000001000",
			1109 => "0010111011110100000100",
			1110 => "0000000001000110011101",
			1111 => "0000001001000110011101",
			1112 => "0001110101110100000100",
			1113 => "1111111001000110011101",
			1114 => "1111110001000110011101",
			1115 => "0001010111011000010000",
			1116 => "0001000110001100001000",
			1117 => "0011001001110100000100",
			1118 => "0000011001000110011101",
			1119 => "0000001001000110011101",
			1120 => "0011101011110000000100",
			1121 => "0000000001000110011101",
			1122 => "0000001001000110011101",
			1123 => "1111111001000110011101",
			1124 => "0001001011110000000100",
			1125 => "0000001001000110011101",
			1126 => "1111111001000110011101",
			1127 => "0010111010011100000100",
			1128 => "1111111001001000000001",
			1129 => "0001011111010100101100",
			1130 => "0010010010101100100100",
			1131 => "0001100100110100000100",
			1132 => "1111111001001000000001",
			1133 => "0000001101010000010000",
			1134 => "0001101000010000001000",
			1135 => "0011111011110000000100",
			1136 => "0000000001001000000001",
			1137 => "1111111001001000000001",
			1138 => "0001111000011000000100",
			1139 => "0000000001001000000001",
			1140 => "0000001001001000000001",
			1141 => "0011101110100100001000",
			1142 => "0011101000011100000100",
			1143 => "1111111001001000000001",
			1144 => "0000000001001000000001",
			1145 => "0001010011001000000100",
			1146 => "1111111001001000000001",
			1147 => "0000001001001000000001",
			1148 => "0010110110110100000100",
			1149 => "0000000001001000000001",
			1150 => "1111111001001000000001",
			1151 => "1111111001001000000001",
			1152 => "0010010111101100110000",
			1153 => "0011001000000000001000",
			1154 => "0011111000000100000100",
			1155 => "1111111001001011100101",
			1156 => "0000000001001011100101",
			1157 => "0011011010000100100000",
			1158 => "0000010101011100010000",
			1159 => "0011000110100100001000",
			1160 => "0000011101011100000100",
			1161 => "0000000001001011100101",
			1162 => "0000000001001011100101",
			1163 => "0011100010010100000100",
			1164 => "0000000001001011100101",
			1165 => "0000000001001011100101",
			1166 => "0000000010101000000100",
			1167 => "0000000001001011100101",
			1168 => "0001000011010100001000",
			1169 => "0010101010110000000100",
			1170 => "0000001001001011100101",
			1171 => "0000000001001011100101",
			1172 => "0000000001001011100101",
			1173 => "0011100101000000000100",
			1174 => "0000000001001011100101",
			1175 => "0000000001001011100101",
			1176 => "0000111000100000011100",
			1177 => "0001011100100100010100",
			1178 => "0001001011101100001100",
			1179 => "0010010000001000000100",
			1180 => "0000000001001011100101",
			1181 => "0011101110110100000100",
			1182 => "0000000001001011100101",
			1183 => "0000000001001011100101",
			1184 => "0011001010111000000100",
			1185 => "0000000001001011100101",
			1186 => "0000000001001011100101",
			1187 => "0000000111000100000100",
			1188 => "0000000001001011100101",
			1189 => "0000001001001011100101",
			1190 => "0010000001010100000100",
			1191 => "0000000001001011100101",
			1192 => "0010000001110000010000",
			1193 => "0010010010101100001100",
			1194 => "0001010001000000000100",
			1195 => "0000000001001011100101",
			1196 => "0001010111111100000100",
			1197 => "0000001001001011100101",
			1198 => "0000000001001011100101",
			1199 => "0000000001001011100101",
			1200 => "0011011100010100000100",
			1201 => "1111111001001011100101",
			1202 => "0001001110111000001000",
			1203 => "0011001000011000000100",
			1204 => "0000001001001011100101",
			1205 => "0000000001001011100101",
			1206 => "0011100011110000000100",
			1207 => "0000000001001011100101",
			1208 => "0000000001001011100101",
			1209 => "0000011101111101000000",
			1210 => "0011000100011000001000",
			1211 => "0000110010010100000100",
			1212 => "1111111001001111011001",
			1213 => "0000000001001111011001",
			1214 => "0001000101000000010100",
			1215 => "0001101001100100001100",
			1216 => "0000101010001000001000",
			1217 => "0001000010000000000100",
			1218 => "0000000001001111011001",
			1219 => "0000000001001111011001",
			1220 => "1111111001001111011001",
			1221 => "0010110110110100000100",
			1222 => "0000000001001111011001",
			1223 => "0000001001001111011001",
			1224 => "0011101000011100010000",
			1225 => "0010011001111100001100",
			1226 => "0010011000010000000100",
			1227 => "0000000001001111011001",
			1228 => "0000001000101100000100",
			1229 => "0000000001001111011001",
			1230 => "0000000001001111011001",
			1231 => "1111111001001111011001",
			1232 => "0010110111100000001100",
			1233 => "0000111110100100000100",
			1234 => "0000000001001111011001",
			1235 => "0000001100001000000100",
			1236 => "0000001001001111011001",
			1237 => "0000000001001111011001",
			1238 => "0011011111100100000100",
			1239 => "0000000001001111011001",
			1240 => "0000000001001111011001",
			1241 => "0011001000011000110000",
			1242 => "0011010111111100010100",
			1243 => "0001100100111100010000",
			1244 => "0001001111101000001000",
			1245 => "0010011010100000000100",
			1246 => "0000000001001111011001",
			1247 => "0000001001001111011001",
			1248 => "0011001011000000000100",
			1249 => "0000000001001111011001",
			1250 => "0000000001001111011001",
			1251 => "1111111001001111011001",
			1252 => "0000000010101000001000",
			1253 => "0010110010001000000100",
			1254 => "0000000001001111011001",
			1255 => "0000000001001111011001",
			1256 => "0011101111101000001000",
			1257 => "0000001000101100000100",
			1258 => "0000001001001111011001",
			1259 => "0000000001001111011001",
			1260 => "0001001100001100000100",
			1261 => "1111111001001111011001",
			1262 => "0011010011001000000100",
			1263 => "0000000001001111011001",
			1264 => "0000001001001111011001",
			1265 => "0000010100110100000100",
			1266 => "0000000001001111011001",
			1267 => "0011100010111000000100",
			1268 => "1111111001001111011001",
			1269 => "0000000001001111011001",
			1270 => "0000011101111101000100",
			1271 => "0011000100011000001000",
			1272 => "0000110010010100000100",
			1273 => "1111111001010011010101",
			1274 => "0000000001010011010101",
			1275 => "0001000101000000011000",
			1276 => "0000111011111000001000",
			1277 => "0011111010001000000100",
			1278 => "0000000001010011010101",
			1279 => "0000000001010011010101",
			1280 => "0001010111111100001100",
			1281 => "0000000110001000000100",
			1282 => "0000000001010011010101",
			1283 => "0000010001111000000100",
			1284 => "0000001001010011010101",
			1285 => "0000000001010011010101",
			1286 => "0000000001010011010101",
			1287 => "0011101000011100010000",
			1288 => "0010011001111100001100",
			1289 => "0010011000010000000100",
			1290 => "0000000001010011010101",
			1291 => "0001011100010100000100",
			1292 => "0000000001010011010101",
			1293 => "0000000001010011010101",
			1294 => "1111111001010011010101",
			1295 => "0010110111100000001100",
			1296 => "0000111110100100000100",
			1297 => "0000000001010011010101",
			1298 => "0000001100001000000100",
			1299 => "0000001001010011010101",
			1300 => "0000000001010011010101",
			1301 => "0011011111100100000100",
			1302 => "0000000001010011010101",
			1303 => "0000000001010011010101",
			1304 => "0011001000011000110000",
			1305 => "0011010100101000010100",
			1306 => "0010100111110100001000",
			1307 => "0010011010100000000100",
			1308 => "0000000001010011010101",
			1309 => "0000001001010011010101",
			1310 => "0010011010100100001000",
			1311 => "0000011101111100000100",
			1312 => "0000000001010011010101",
			1313 => "1111111001010011010101",
			1314 => "0000000001010011010101",
			1315 => "0011110011000000001000",
			1316 => "0010011010100100000100",
			1317 => "0000000001010011010101",
			1318 => "0000001001010011010101",
			1319 => "0000000111000000001000",
			1320 => "0000011010011000000100",
			1321 => "1111111001010011010101",
			1322 => "0000000001010011010101",
			1323 => "0001011001010000000100",
			1324 => "0000000001010011010101",
			1325 => "0010001001101000000100",
			1326 => "0000001001010011010101",
			1327 => "0000000001010011010101",
			1328 => "0000010100110100000100",
			1329 => "0000000001010011010101",
			1330 => "0011100010111000000100",
			1331 => "1111111001010011010101",
			1332 => "0000000001010011010101",
			1333 => "0011001010111000001000",
			1334 => "0000011100011000000100",
			1335 => "1111111001010110100001",
			1336 => "0000000001010110100001",
			1337 => "0001000011001101000000",
			1338 => "0010101000010100100100",
			1339 => "0001011110101100001100",
			1340 => "0001000110101100001000",
			1341 => "0000000001010100000100",
			1342 => "0000000001010110100001",
			1343 => "0000001001010110100001",
			1344 => "0000000001010110100001",
			1345 => "0000001111001000001000",
			1346 => "0010110100000100000100",
			1347 => "0000000001010110100001",
			1348 => "1111111001010110100001",
			1349 => "0000101100111000001000",
			1350 => "0011010101110000000100",
			1351 => "0000000001010110100001",
			1352 => "0000001001010110100001",
			1353 => "0000000010101000000100",
			1354 => "0000000001010110100001",
			1355 => "0000000001010110100001",
			1356 => "0011010010000100010100",
			1357 => "0001111000011000001000",
			1358 => "0001110110100100000100",
			1359 => "0000000001010110100001",
			1360 => "0000000001010110100001",
			1361 => "0010100001010000001000",
			1362 => "0011011001011100000100",
			1363 => "0000000001010110100001",
			1364 => "0000001001010110100001",
			1365 => "0000000001010110100001",
			1366 => "0010001100000100000100",
			1367 => "0000000001010110100001",
			1368 => "0000000001010110100001",
			1369 => "0011101000110100001000",
			1370 => "0001000011001100000100",
			1371 => "0000000001010110100001",
			1372 => "1111111001010110100001",
			1373 => "0001011100010000010000",
			1374 => "0010011010100100001100",
			1375 => "0001011110010000000100",
			1376 => "0000000001010110100001",
			1377 => "0000100011110100000100",
			1378 => "0000001001010110100001",
			1379 => "0000000001010110100001",
			1380 => "0000000001010110100001",
			1381 => "0001101001111100000100",
			1382 => "1111111001010110100001",
			1383 => "0000000001010110100001",
			1384 => "0000010101011100011100",
			1385 => "0000000111000000011000",
			1386 => "0000000001010100000100",
			1387 => "1111111001011001100101",
			1388 => "0000000001010100000100",
			1389 => "0000000001011001100101",
			1390 => "0000000111000000001100",
			1391 => "0000000110001000000100",
			1392 => "1111111001011001100101",
			1393 => "0000001111001000000100",
			1394 => "0000010001011001100101",
			1395 => "1111111001011001100101",
			1396 => "0000000001011001100101",
			1397 => "1111111001011001100101",
			1398 => "0000011100011001000000",
			1399 => "0001011001010000100000",
			1400 => "0001001011110000011100",
			1401 => "0000011101111100010000",
			1402 => "0010000110011100001000",
			1403 => "0000101100000000000100",
			1404 => "0000000001011001100101",
			1405 => "1111111001011001100101",
			1406 => "0001011100100100000100",
			1407 => "1111111001011001100101",
			1408 => "0000101001011001100101",
			1409 => "0010000110011100000100",
			1410 => "0000100001011001100101",
			1411 => "0000010100110100000100",
			1412 => "1111111001011001100101",
			1413 => "0000001001011001100101",
			1414 => "1111111001011001100101",
			1415 => "0001100100111100001100",
			1416 => "0010110101110100000100",
			1417 => "0000010001011001100101",
			1418 => "0000000111000000000100",
			1419 => "1111111001011001100101",
			1420 => "1111110001011001100101",
			1421 => "0000101110000000001000",
			1422 => "0001001000011100000100",
			1423 => "0000000001011001100101",
			1424 => "0000011001011001100101",
			1425 => "0010111100100100001000",
			1426 => "0011100010010100000100",
			1427 => "1111111001011001100101",
			1428 => "0000001001011001100101",
			1429 => "0000000001011001100101",
			1430 => "0000110001011100000100",
			1431 => "0000010001011001100101",
			1432 => "1111111001011001100101",
			1433 => "0011001101010100000100",
			1434 => "1111111001011100010001",
			1435 => "0010011010100101000000",
			1436 => "0010110111010000010000",
			1437 => "0000000110001000001100",
			1438 => "0001100100110100000100",
			1439 => "0000000001011100010001",
			1440 => "0001110011100000000100",
			1441 => "0000000001011100010001",
			1442 => "0000001001011100010001",
			1443 => "0000000001011100010001",
			1444 => "0010110110110100011000",
			1445 => "0010110100000100001100",
			1446 => "0000100110111100001000",
			1447 => "0000101100010000000100",
			1448 => "0000000001011100010001",
			1449 => "0000000001011100010001",
			1450 => "0000000001011100010001",
			1451 => "0001011100100100000100",
			1452 => "1111111001011100010001",
			1453 => "0001010111100000000100",
			1454 => "0000000001011100010001",
			1455 => "0000000001011100010001",
			1456 => "0000111100111000001100",
			1457 => "0001101001100100000100",
			1458 => "0000000001011100010001",
			1459 => "0000000010101000000100",
			1460 => "0000001001011100010001",
			1461 => "0000000001011100010001",
			1462 => "0001111111011100000100",
			1463 => "1111111001011100010001",
			1464 => "0011010111010100000100",
			1465 => "0000000001011100010001",
			1466 => "0000000001011100010001",
			1467 => "0011001000000000010000",
			1468 => "0011001011000000001000",
			1469 => "0010110101100100000100",
			1470 => "0000000001011100010001",
			1471 => "0000000001011100010001",
			1472 => "0000001101010000000100",
			1473 => "0000001001011100010001",
			1474 => "0000000001011100010001",
			1475 => "1111111001011100010001",
			1476 => "0011001101010100000100",
			1477 => "1111111001011111011101",
			1478 => "0010011010100000101100",
			1479 => "0001111111011100001100",
			1480 => "0000101110010000001000",
			1481 => "0001100100110100000100",
			1482 => "0000000001011111011101",
			1483 => "0000000001011111011101",
			1484 => "1111111001011111011101",
			1485 => "0011010111010100011000",
			1486 => "0011100110111000010000",
			1487 => "0001111011011100001000",
			1488 => "0000001000110000000100",
			1489 => "0000000001011111011101",
			1490 => "0000000001011111011101",
			1491 => "0001100101010000000100",
			1492 => "1111111001011111011101",
			1493 => "0000000001011111011101",
			1494 => "0000000011010000000100",
			1495 => "0000001001011111011101",
			1496 => "0000000001011111011101",
			1497 => "0000010111101000000100",
			1498 => "1111111001011111011101",
			1499 => "0000000001011111011101",
			1500 => "0011001000000000010100",
			1501 => "0010011010100100001000",
			1502 => "0001101111000000000100",
			1503 => "0000000001011111011101",
			1504 => "1111111001011111011101",
			1505 => "0000001000101100001000",
			1506 => "0010111011011100000100",
			1507 => "0000000001011111011101",
			1508 => "0000001001011111011101",
			1509 => "0000000001011111011101",
			1510 => "0010000001110000001100",
			1511 => "0010011010100100001000",
			1512 => "0010011010100100000100",
			1513 => "0000000001011111011101",
			1514 => "0000000001011111011101",
			1515 => "1111111001011111011101",
			1516 => "0011011110110100001100",
			1517 => "0010001100000100001000",
			1518 => "0000010100110100000100",
			1519 => "0000000001011111011101",
			1520 => "0000000001011111011101",
			1521 => "0000000001011111011101",
			1522 => "0011101110000000000100",
			1523 => "0000000001011111011101",
			1524 => "0000011100011000000100",
			1525 => "0000001001011111011101",
			1526 => "0000000001011111011101",
			1527 => "0001110011100000000100",
			1528 => "1111111001100010010001",
			1529 => "0010111010001100010000",
			1530 => "0010100111110100001100",
			1531 => "0001001111100100001000",
			1532 => "0011111001011100000100",
			1533 => "0000000001100010010001",
			1534 => "0000001001100010010001",
			1535 => "0000000001100010010001",
			1536 => "0000000001100010010001",
			1537 => "0000011100011000110000",
			1538 => "0011100010010100011100",
			1539 => "0000101000100000010000",
			1540 => "0001000001011100001000",
			1541 => "0010110100000100000100",
			1542 => "0000000001100010010001",
			1543 => "1111111001100010010001",
			1544 => "0001011100100100000100",
			1545 => "0000000001100010010001",
			1546 => "0000001001100010010001",
			1547 => "0011001001001000000100",
			1548 => "1111111001100010010001",
			1549 => "0001111111011100000100",
			1550 => "0000000001100010010001",
			1551 => "1111111001100010010001",
			1552 => "0010110001000000001100",
			1553 => "0001101000010000000100",
			1554 => "1111111001100010010001",
			1555 => "0010111011110100000100",
			1556 => "0000000001100010010001",
			1557 => "0000001001100010010001",
			1558 => "0001011111010100000100",
			1559 => "0000000001100010010001",
			1560 => "1111111001100010010001",
			1561 => "0001110000011100010100",
			1562 => "0010110010001000001000",
			1563 => "0001101000010000000100",
			1564 => "0000000001100010010001",
			1565 => "0000000001100010010001",
			1566 => "0010001001101000001000",
			1567 => "0010010010101100000100",
			1568 => "0000001001100010010001",
			1569 => "0000000001100010010001",
			1570 => "0000000001100010010001",
			1571 => "1111111001100010010001",
			1572 => "0011001010111000001000",
			1573 => "0010010010101100000100",
			1574 => "1111111001100100111101",
			1575 => "0000000001100100111101",
			1576 => "0011011111100101001100",
			1577 => "0011100101000000111100",
			1578 => "0000101110000000100000",
			1579 => "0000000111000000010000",
			1580 => "0011101101101100001000",
			1581 => "0001001111101000000100",
			1582 => "0000000001100100111101",
			1583 => "0000001001100100111101",
			1584 => "0000011101111100000100",
			1585 => "0000000001100100111101",
			1586 => "1111111001100100111101",
			1587 => "0010011010100100001000",
			1588 => "0001110111010000000100",
			1589 => "1111111001100100111101",
			1590 => "0000000001100100111101",
			1591 => "0011000001101000000100",
			1592 => "0000001001100100111101",
			1593 => "0000000001100100111101",
			1594 => "0011101011110000010000",
			1595 => "0000101000110100001000",
			1596 => "0000010111101000000100",
			1597 => "0000000001100100111101",
			1598 => "0000000001100100111101",
			1599 => "0010101001000100000100",
			1600 => "0000000001100100111101",
			1601 => "1111111001100100111101",
			1602 => "0010001100000100000100",
			1603 => "1111111001100100111101",
			1604 => "0010001001101000000100",
			1605 => "0000001001100100111101",
			1606 => "1111111001100100111101",
			1607 => "0000011100011000001100",
			1608 => "0000001011000100001000",
			1609 => "0001110111010000000100",
			1610 => "0000000001100100111101",
			1611 => "0000001001100100111101",
			1612 => "0000000001100100111101",
			1613 => "0000000001100100111101",
			1614 => "1111111001100100111101",
			1615 => "0000011101011100000100",
			1616 => "1111111001100111010011",
			1617 => "0010010010101101000000",
			1618 => "0001101011001100000100",
			1619 => "1111111001100111010011",
			1620 => "0001001011110000011100",
			1621 => "0001011100100100010000",
			1622 => "0001001111100100001000",
			1623 => "0010010111101100000100",
			1624 => "0000000001100111010011",
			1625 => "0000001001100111010011",
			1626 => "0010011010100100000100",
			1627 => "1111111001100111010011",
			1628 => "0000000001100111010011",
			1629 => "0000111101101100001000",
			1630 => "0000000110001000000100",
			1631 => "0000000001100111010011",
			1632 => "0000010001100111010011",
			1633 => "0000000001100111010011",
			1634 => "0000000111000000010000",
			1635 => "0000110001011100001000",
			1636 => "0001100100111100000100",
			1637 => "1111111001100111010011",
			1638 => "0000001001100111010011",
			1639 => "0000000111000000000100",
			1640 => "1111111001100111010011",
			1641 => "0000000001100111010011",
			1642 => "0000001000101100001000",
			1643 => "0010101000010100000100",
			1644 => "1111111001100111010011",
			1645 => "0000001001100111010011",
			1646 => "0001010111111100000100",
			1647 => "1111111001100111010011",
			1648 => "0000000001100111010011",
			1649 => "0011010100101000000100",
			1650 => "0000000001100111010011",
			1651 => "1111111001100111010011",
			1652 => "0000000001100111010101",
			1653 => "0000000001100111011001",
			1654 => "0000000001100111011101",
			1655 => "0000000001100111100001",
			1656 => "0000000001100111100101",
			1657 => "0000000001100111101001",
			1658 => "0000000001100111101101",
			1659 => "0000000001100111110001",
			1660 => "0000000001100111110101",
			1661 => "0000000001100111111001",
			1662 => "0000000001100111111101",
			1663 => "0000000001101000000001",
			1664 => "0000000001101000000101",
			1665 => "0000000001101000001001",
			1666 => "0000000001101000001101",
			1667 => "0000000001101000010001",
			1668 => "0000000001101000010101",
			1669 => "0000000001101000011001",
			1670 => "0000000001101000011101",
			1671 => "0000000001101000100001",
			1672 => "0001100100111100000100",
			1673 => "0000000001101000110101",
			1674 => "0001101001111100000100",
			1675 => "0000000001101000110101",
			1676 => "0000000001101000110101",
			1677 => "0011101100001100001000",
			1678 => "0000111011101100000100",
			1679 => "0000000001101001001001",
			1680 => "0000000001101001001001",
			1681 => "0000000001101001001001",
			1682 => "0001100100111100000100",
			1683 => "0000000001101001011101",
			1684 => "0001101001111100000100",
			1685 => "0000000001101001011101",
			1686 => "0000000001101001011101",
			1687 => "0010001011010100001000",
			1688 => "0010001010110000000100",
			1689 => "0000000001101001110001",
			1690 => "0000000001101001110001",
			1691 => "0000000001101001110001",
			1692 => "0001111111011100001000",
			1693 => "0001110001101000000100",
			1694 => "0000000001101010001101",
			1695 => "0000000001101010001101",
			1696 => "0001110100010000000100",
			1697 => "0000000001101010001101",
			1698 => "0000000001101010001101",
			1699 => "0000000010101000001100",
			1700 => "0000000010101000000100",
			1701 => "0000000001101010101001",
			1702 => "0010000101000100000100",
			1703 => "0000000001101010101001",
			1704 => "0000000001101010101001",
			1705 => "0000000001101010101001",
			1706 => "0011011111100100001100",
			1707 => "0010111011110100000100",
			1708 => "0000000001101011000101",
			1709 => "0011010011001000000100",
			1710 => "0000000001101011000101",
			1711 => "0000000001101011000101",
			1712 => "0000000001101011000101",
			1713 => "0000011100011000001100",
			1714 => "0001111000011000000100",
			1715 => "0000000001101011100001",
			1716 => "0000000011111100000100",
			1717 => "0000000001101011100001",
			1718 => "0000000001101011100001",
			1719 => "0000000001101011100001",
			1720 => "0010011010100000000100",
			1721 => "0000000001101011111101",
			1722 => "0001010111011000001000",
			1723 => "0010010011101000000100",
			1724 => "0000000001101011111101",
			1725 => "0000000001101011111101",
			1726 => "0000000001101011111101",
			1727 => "0000001101010000010000",
			1728 => "0010011010100000000100",
			1729 => "0000000001101100100001",
			1730 => "0011001001110100001000",
			1731 => "0010101001000100000100",
			1732 => "0000000001101100100001",
			1733 => "0000000001101100100001",
			1734 => "0000000001101100100001",
			1735 => "0000000001101100100001",
			1736 => "0000110011110000010000",
			1737 => "0001001011110000000100",
			1738 => "0000000001101101000101",
			1739 => "0000011100011000001000",
			1740 => "0000010111101000000100",
			1741 => "0000000001101101000101",
			1742 => "0000000001101101000101",
			1743 => "0000000001101101000101",
			1744 => "0000000001101101000101",
			1745 => "0001001000011100010000",
			1746 => "0010010000001000000100",
			1747 => "0000000001101101110001",
			1748 => "0000110010010100001000",
			1749 => "0010100011101000000100",
			1750 => "0000000001101101110001",
			1751 => "0000000001101101110001",
			1752 => "0000000001101101110001",
			1753 => "0010010100101100000100",
			1754 => "0000000001101101110001",
			1755 => "0000000001101101110001",
			1756 => "0000000010101000010000",
			1757 => "0011110011000000001100",
			1758 => "0010001010110000000100",
			1759 => "0000000001101110011101",
			1760 => "0011111100010000000100",
			1761 => "0000000001101110011101",
			1762 => "0000000001101110011101",
			1763 => "0000000001101110011101",
			1764 => "0000100011110100000100",
			1765 => "0000000001101110011101",
			1766 => "0000000001101110011101",
			1767 => "0000001010101100001100",
			1768 => "0010011010100100000100",
			1769 => "0000000001101111011001",
			1770 => "0000100001011100000100",
			1771 => "0000000001101111011001",
			1772 => "0000000001101111011001",
			1773 => "0011101110000000001000",
			1774 => "0000011100011000000100",
			1775 => "0000000001101111011001",
			1776 => "0000000001101111011001",
			1777 => "0011011111100100001000",
			1778 => "0001110111010000000100",
			1779 => "0000000001101111011001",
			1780 => "0000000001101111011001",
			1781 => "0000000001101111011001",
			1782 => "0001110001101000010100",
			1783 => "0000000010101000010000",
			1784 => "0000111100111000001100",
			1785 => "0001111000000000000100",
			1786 => "0000000001110000001101",
			1787 => "0000000001010100000100",
			1788 => "0000000001110000001101",
			1789 => "0000000001110000001101",
			1790 => "0000000001110000001101",
			1791 => "0000000001110000001101",
			1792 => "0001110111010000000100",
			1793 => "0000000001110000001101",
			1794 => "0000000001110000001101",
			1795 => "0010011010100000000100",
			1796 => "0000000001110000111001",
			1797 => "0011001000011000010000",
			1798 => "0001101001111100001100",
			1799 => "0010010011101000001000",
			1800 => "0010011010100000000100",
			1801 => "0000000001110000111001",
			1802 => "0000000001110000111001",
			1803 => "0000000001110000111001",
			1804 => "0000000001110000111001",
			1805 => "0000000001110000111001",
			1806 => "0010000001010100010100",
			1807 => "0001011100100100000100",
			1808 => "0000000001110001111101",
			1809 => "0000001111001000000100",
			1810 => "0000000001110001111101",
			1811 => "0010110101110100001000",
			1812 => "0000101000101000000100",
			1813 => "0000000001110001111101",
			1814 => "0000000001110001111101",
			1815 => "0000000001110001111101",
			1816 => "0011101110000000001100",
			1817 => "0000011100011000001000",
			1818 => "0001001000110100000100",
			1819 => "0000000001110001111101",
			1820 => "0000000001110001111101",
			1821 => "0000000001110001111101",
			1822 => "0000000001110001111101",
			1823 => "0010000001010100011000",
			1824 => "0001011100100100001000",
			1825 => "0000000001110000000100",
			1826 => "0000000001110011010001",
			1827 => "0000000001110011010001",
			1828 => "0000001111001000000100",
			1829 => "0000000001110011010001",
			1830 => "0000110010010100001000",
			1831 => "0001110000011100000100",
			1832 => "0000000001110011010001",
			1833 => "0000000001110011010001",
			1834 => "0000000001110011010001",
			1835 => "0001010111111100001000",
			1836 => "0001000110111000000100",
			1837 => "0000000001110011010001",
			1838 => "0000000001110011010001",
			1839 => "0001001110111000001000",
			1840 => "0001000110001100000100",
			1841 => "0000000001110011010001",
			1842 => "0000000001110011010001",
			1843 => "0000000001110011010001",
			1844 => "0001001011110000011000",
			1845 => "0011101011101100010100",
			1846 => "0001111000000000000100",
			1847 => "0000000001110100001101",
			1848 => "0010001000100100000100",
			1849 => "0000000001110100001101",
			1850 => "0011011100010100001000",
			1851 => "0010101000010100000100",
			1852 => "0000000001110100001101",
			1853 => "0000000001110100001101",
			1854 => "0000000001110100001101",
			1855 => "0000000001110100001101",
			1856 => "0011100010010100000100",
			1857 => "0000000001110100001101",
			1858 => "0000000001110100001101",
			1859 => "0010001100000100011000",
			1860 => "0001101011001100000100",
			1861 => "0000000001110101001001",
			1862 => "0011011110110100010000",
			1863 => "0000101000011100001100",
			1864 => "0001011100100100000100",
			1865 => "0000000001110101001001",
			1866 => "0010001100011100000100",
			1867 => "0000000001110101001001",
			1868 => "0000000001110101001001",
			1869 => "0000000001110101001001",
			1870 => "0000000001110101001001",
			1871 => "0000100011110100000100",
			1872 => "0000000001110101001001",
			1873 => "0000000001110101001001",
			1874 => "0011011111100100011000",
			1875 => "0000010101011100000100",
			1876 => "0000000001110101111101",
			1877 => "0001111111011100000100",
			1878 => "0000000001110101111101",
			1879 => "0000010100110100001100",
			1880 => "0011010011001000000100",
			1881 => "0000000001110101111101",
			1882 => "0001101000010000000100",
			1883 => "0000000001110101111101",
			1884 => "0000000001110101111101",
			1885 => "0000000001110101111101",
			1886 => "0000000001110101111101",
			1887 => "0001011001010000000100",
			1888 => "0000000001110110110001",
			1889 => "0011011011111000010100",
			1890 => "0010010010101100010000",
			1891 => "0011011110010000000100",
			1892 => "0000000001110110110001",
			1893 => "0001101001100100000100",
			1894 => "0000000001110110110001",
			1895 => "0010100110011100000100",
			1896 => "0000000001110110110001",
			1897 => "0000000001110110110001",
			1898 => "0000000001110110110001",
			1899 => "0000000001110110110001",
			1900 => "0000001010101100011000",
			1901 => "0010110101110100010100",
			1902 => "0011001001110100010000",
			1903 => "0001100100110100000100",
			1904 => "0000000001110111111101",
			1905 => "0011001010111000000100",
			1906 => "0000000001110111111101",
			1907 => "0000101000101000000100",
			1908 => "0000000001110111111101",
			1909 => "0000000001110111111101",
			1910 => "0000000001110111111101",
			1911 => "0000000001110111111101",
			1912 => "0001101000010000000100",
			1913 => "0000000001110111111101",
			1914 => "0010101010110000001000",
			1915 => "0010101001000100000100",
			1916 => "0000000001110111111101",
			1917 => "0000000001110111111101",
			1918 => "0000000001110111111101",
			1919 => "0001111000011000100000",
			1920 => "0011000100011000001100",
			1921 => "0001001000100000000100",
			1922 => "0000000001111001011001",
			1923 => "0000011100011000000100",
			1924 => "0000000001111001011001",
			1925 => "0000000001111001011001",
			1926 => "0011001000000000010000",
			1927 => "0000001000101100001100",
			1928 => "0001110110100100000100",
			1929 => "0000000001111001011001",
			1930 => "0001100100110100000100",
			1931 => "0000000001111001011001",
			1932 => "0000000001111001011001",
			1933 => "0000000001111001011001",
			1934 => "0000000001111001011001",
			1935 => "0000100011110100001100",
			1936 => "0000010111101000000100",
			1937 => "0000000001111001011001",
			1938 => "0001101001111100000100",
			1939 => "0000000001111001011001",
			1940 => "0000000001111001011001",
			1941 => "0000000001111001011001",
			1942 => "0001001110111000100000",
			1943 => "0010111011011100001000",
			1944 => "0001001011101100000100",
			1945 => "0000000001111010100101",
			1946 => "0000000001111010100101",
			1947 => "0001110100010000010100",
			1948 => "0001101001100100000100",
			1949 => "0000000001111010100101",
			1950 => "0010010011101000001100",
			1951 => "0011000100011000000100",
			1952 => "0000000001111010100101",
			1953 => "0010001011010100000100",
			1954 => "0000000001111010100101",
			1955 => "0000000001111010100101",
			1956 => "0000000001111010100101",
			1957 => "0000000001111010100101",
			1958 => "0010101100011100000100",
			1959 => "0000000001111010100101",
			1960 => "0000000001111010100101",
			1961 => "0011001011000000001000",
			1962 => "0011101000101000000100",
			1963 => "0000000001111011101001",
			1964 => "0000000001111011101001",
			1965 => "0011011111100100011000",
			1966 => "0010110010001000000100",
			1967 => "0000000001111011101001",
			1968 => "0001001011110000000100",
			1969 => "0000000001111011101001",
			1970 => "0010110010110100001100",
			1971 => "0001001001001100001000",
			1972 => "0011011010001000000100",
			1973 => "0000000001111011101001",
			1974 => "0000000001111011101001",
			1975 => "0000000001111011101001",
			1976 => "0000000001111011101001",
			1977 => "0000000001111011101001",
			1978 => "0000000010101000010100",
			1979 => "0010010000001000000100",
			1980 => "0000000001111101001101",
			1981 => "0001111000011000001100",
			1982 => "0000101000101000001000",
			1983 => "0011100110010000000100",
			1984 => "0000000001111101001101",
			1985 => "0000000001111101001101",
			1986 => "0000000001111101001101",
			1987 => "0000000001111101001101",
			1988 => "0001111111011100000100",
			1989 => "0000000001111101001101",
			1990 => "0001110101100100001100",
			1991 => "0010001011010100001000",
			1992 => "0010010010101100000100",
			1993 => "0000000001111101001101",
			1994 => "0000000001111101001101",
			1995 => "0000000001111101001101",
			1996 => "0001100101010000001000",
			1997 => "0001000110001100000100",
			1998 => "0000000001111101001101",
			1999 => "0000000001111101001101",
			2000 => "0001101001111100000100",
			2001 => "0000000001111101001101",
			2002 => "0000000001111101001101",
			2003 => "0010000110011100010100",
			2004 => "0010100011101000000100",
			2005 => "0000000001111111000001",
			2006 => "0010100111110100001100",
			2007 => "0001101111000000001000",
			2008 => "0001101011001100000100",
			2009 => "0000000001111111000001",
			2010 => "0000000001111111000001",
			2011 => "0000000001111111000001",
			2012 => "0000000001111111000001",
			2013 => "0001101000010000001100",
			2014 => "0010011010100100001000",
			2015 => "0000010001000100000100",
			2016 => "0000000001111111000001",
			2017 => "0000000001111111000001",
			2018 => "0000000001111111000001",
			2019 => "0001001001001100010000",
			2020 => "0001111000011000000100",
			2021 => "0000000001111111000001",
			2022 => "0010001001101000001000",
			2023 => "0010101000010100000100",
			2024 => "0000000001111111000001",
			2025 => "0000000001111111000001",
			2026 => "0000000001111111000001",
			2027 => "0010101010110000001000",
			2028 => "0001001110111000000100",
			2029 => "0000000001111111000001",
			2030 => "0000000001111111000001",
			2031 => "0000000001111111000001",
			2032 => "0001111000011000100000",
			2033 => "0010000001110000011000",
			2034 => "0011001000000000010100",
			2035 => "0011000100011000000100",
			2036 => "0000000010000000110101",
			2037 => "0001101000010000001100",
			2038 => "0001110110100100000100",
			2039 => "0000000010000000110101",
			2040 => "0001100100110100000100",
			2041 => "0000000010000000110101",
			2042 => "0000000010000000110101",
			2043 => "0000000010000000110101",
			2044 => "0000000010000000110101",
			2045 => "0010110101110100000100",
			2046 => "0000000010000000110101",
			2047 => "0000000010000000110101",
			2048 => "0011101111101000001100",
			2049 => "0000011100011000001000",
			2050 => "0001110111010000000100",
			2051 => "0000000010000000110101",
			2052 => "0000000010000000110101",
			2053 => "0000000010000000110101",
			2054 => "0010110001000000001100",
			2055 => "0001111111011100000100",
			2056 => "0000000010000000110101",
			2057 => "0001011001010000000100",
			2058 => "0000000010000000110101",
			2059 => "0000000010000000110101",
			2060 => "0000000010000000110101",
			2061 => "0010010111101100001100",
			2062 => "0011001000000000001000",
			2063 => "0011101000101000000100",
			2064 => "0000000010000010100001",
			2065 => "0000000010000010100001",
			2066 => "0000000010000010100001",
			2067 => "0011000100011000010000",
			2068 => "0010000001010100001100",
			2069 => "0010010000001000000100",
			2070 => "0000000010000010100001",
			2071 => "0011100110010000000100",
			2072 => "0000000010000010100001",
			2073 => "0000000010000010100001",
			2074 => "0000000010000010100001",
			2075 => "0001101000010000001000",
			2076 => "0000111000100000000100",
			2077 => "0000000010000010100001",
			2078 => "0000000010000010100001",
			2079 => "0010110001000000010000",
			2080 => "0001010010011100000100",
			2081 => "0000000010000010100001",
			2082 => "0011100011000000000100",
			2083 => "0000000010000010100001",
			2084 => "0010100110011100000100",
			2085 => "0000000010000010100001",
			2086 => "0000000010000010100001",
			2087 => "0000000010000010100001",
			2088 => "0010000001110000011100",
			2089 => "0011011100010100010100",
			2090 => "0011000100011000000100",
			2091 => "0000000010000100010101",
			2092 => "0011010101110000000100",
			2093 => "0000000010000100010101",
			2094 => "0000000111000100000100",
			2095 => "0000000010000100010101",
			2096 => "0001101000010000000100",
			2097 => "0000000010000100010101",
			2098 => "0000000010000100010101",
			2099 => "0001100100111100000100",
			2100 => "0000000010000100010101",
			2101 => "0000000010000100010101",
			2102 => "0001111111011100000100",
			2103 => "0000000010000100010101",
			2104 => "0000010100110100010100",
			2105 => "0000011110010100001000",
			2106 => "0001011110110100000100",
			2107 => "0000000010000100010101",
			2108 => "0000000010000100010101",
			2109 => "0011100011000000000100",
			2110 => "0000000010000100010101",
			2111 => "0001010101110000000100",
			2112 => "0000000010000100010101",
			2113 => "0000000010000100010101",
			2114 => "0011111000110100000100",
			2115 => "0000000010000100010101",
			2116 => "0000000010000100010101",
			2117 => "0010000110011100010100",
			2118 => "0010100011101000000100",
			2119 => "0000000010000110010001",
			2120 => "0010100111110100001100",
			2121 => "0001101111000000001000",
			2122 => "0001101011001100000100",
			2123 => "0000000010000110010001",
			2124 => "0000000010000110010001",
			2125 => "0000000010000110010001",
			2126 => "0000000010000110010001",
			2127 => "0001101000010000001100",
			2128 => "0010011010100100001000",
			2129 => "0010010101010000000100",
			2130 => "0000000010000110010001",
			2131 => "0000000010000110010001",
			2132 => "0000000010000110010001",
			2133 => "0000001101010000010100",
			2134 => "0001111000011000000100",
			2135 => "0000000010000110010001",
			2136 => "0000000111000000000100",
			2137 => "0000000010000110010001",
			2138 => "0001011001010000000100",
			2139 => "0000000010000110010001",
			2140 => "0010000001110000000100",
			2141 => "0000000010000110010001",
			2142 => "0000000010000110010001",
			2143 => "0000000011111100001000",
			2144 => "0010101100011100000100",
			2145 => "0000000010000110010001",
			2146 => "0000000010000110010001",
			2147 => "0000000010000110010001",
			2148 => "0010000001110000101000",
			2149 => "0001110001101000010100",
			2150 => "0010010000001000000100",
			2151 => "0000000010001000011101",
			2152 => "0000001010101100001100",
			2153 => "0000111100111000001000",
			2154 => "0011100110010000000100",
			2155 => "0000000010001000011101",
			2156 => "0000000010001000011101",
			2157 => "0000000010001000011101",
			2158 => "0000000010001000011101",
			2159 => "0000000111000000001100",
			2160 => "0001110111010000001000",
			2161 => "0010110000011100000100",
			2162 => "0000000010001000011101",
			2163 => "0000000010001000011101",
			2164 => "0000000010001000011101",
			2165 => "0011100110111000000100",
			2166 => "0000000010001000011101",
			2167 => "0000000010001000011101",
			2168 => "0001111111011100000100",
			2169 => "0000000010001000011101",
			2170 => "0000010100110100010100",
			2171 => "0000011110010100001000",
			2172 => "0001011110110100000100",
			2173 => "0000000010001000011101",
			2174 => "0000000010001000011101",
			2175 => "0011100011000000000100",
			2176 => "0000000010001000011101",
			2177 => "0001010101110000000100",
			2178 => "0000000010001000011101",
			2179 => "0000000010001000011101",
			2180 => "0011111000110100000100",
			2181 => "0000000010001000011101",
			2182 => "0000000010001000011101",
			2183 => "0000010001111000010000",
			2184 => "0011100001011100001100",
			2185 => "0001001100010000000100",
			2186 => "0000000010001010100001",
			2187 => "0011001111011100000100",
			2188 => "0000000010001010100001",
			2189 => "0000000010001010100001",
			2190 => "0000000010001010100001",
			2191 => "0011101011101100010000",
			2192 => "0001110110100100000100",
			2193 => "0000000010001010100001",
			2194 => "0000000111000100000100",
			2195 => "0000000010001010100001",
			2196 => "0000000010101000000100",
			2197 => "0000000010001010100001",
			2198 => "0000000010001010100001",
			2199 => "0000000111000000001000",
			2200 => "0010000001010100000100",
			2201 => "0000000010001010100001",
			2202 => "0000000010001010100001",
			2203 => "0001110101100100010000",
			2204 => "0001001110111000001100",
			2205 => "0011011010001000000100",
			2206 => "0000000010001010100001",
			2207 => "0001111000011000000100",
			2208 => "0000000010001010100001",
			2209 => "0000000010001010100001",
			2210 => "0000000010001010100001",
			2211 => "0001001110111000001000",
			2212 => "0001111011011100000100",
			2213 => "0000000010001010100001",
			2214 => "0000000010001010100001",
			2215 => "0000000010001010100001",
			2216 => "0001001011110000010000",
			2217 => "0011101011101100001100",
			2218 => "0010110110110100001000",
			2219 => "0010011010100000000100",
			2220 => "0000000010001100001101",
			2221 => "0000000010001100001101",
			2222 => "0000000010001100001101",
			2223 => "0000000010001100001101",
			2224 => "0001011001010000000100",
			2225 => "1111111010001100001101",
			2226 => "0010110001000000100000",
			2227 => "0000000111000000001100",
			2228 => "0011101000101000000100",
			2229 => "0000000010001100001101",
			2230 => "0000000111000000000100",
			2231 => "0000000010001100001101",
			2232 => "0000000010001100001101",
			2233 => "0011101000101000000100",
			2234 => "0000000010001100001101",
			2235 => "0000000010011000001000",
			2236 => "0010010010101100000100",
			2237 => "0000000010001100001101",
			2238 => "0000000010001100001101",
			2239 => "0011100011110000000100",
			2240 => "0000000010001100001101",
			2241 => "0000000010001100001101",
			2242 => "0000000010001100001101",
			2243 => "0001110001101000010100",
			2244 => "0001001000100000001100",
			2245 => "0010101010100000000100",
			2246 => "0000000010001110111001",
			2247 => "0011001101010100000100",
			2248 => "0000000010001110111001",
			2249 => "0000000010001110111001",
			2250 => "0010010010101100000100",
			2251 => "1111111010001110111001",
			2252 => "0000000010001110111001",
			2253 => "0011001001110100011000",
			2254 => "0010110110110100001000",
			2255 => "0000111011111000000100",
			2256 => "0000000010001110111001",
			2257 => "0000000010001110111001",
			2258 => "0010001100000100001000",
			2259 => "0001001111101000000100",
			2260 => "0000000010001110111001",
			2261 => "0000001010001110111001",
			2262 => "0011001001110100000100",
			2263 => "0000000010001110111001",
			2264 => "0000000010001110111001",
			2265 => "0011101000011100011000",
			2266 => "0010010100101100001100",
			2267 => "0001001101001000001000",
			2268 => "0001001000110100000100",
			2269 => "0000000010001110111001",
			2270 => "0000000010001110111001",
			2271 => "0000000010001110111001",
			2272 => "0001010010011100000100",
			2273 => "0000000010001110111001",
			2274 => "0011101110000000000100",
			2275 => "0000000010001110111001",
			2276 => "0000000010001110111001",
			2277 => "0010110111100000010000",
			2278 => "0010000110001000001100",
			2279 => "0010010010101100001000",
			2280 => "0001000010111000000100",
			2281 => "0000000010001110111001",
			2282 => "0000001010001110111001",
			2283 => "0000000010001110111001",
			2284 => "0000000010001110111001",
			2285 => "0000000010001110111001",
			2286 => "0010011010100000011000",
			2287 => "0011101011110000001000",
			2288 => "0000001000101100000100",
			2289 => "0000000010010000111101",
			2290 => "0000000010010000111101",
			2291 => "0001000011110100001100",
			2292 => "0000001000110000000100",
			2293 => "0000000010010000111101",
			2294 => "0001011110010000000100",
			2295 => "0000000010010000111101",
			2296 => "0000000010010000111101",
			2297 => "0000000010010000111101",
			2298 => "0011001011011100101000",
			2299 => "0010111011011100001000",
			2300 => "0001000011000000000100",
			2301 => "0000000010010000111101",
			2302 => "0000000010010000111101",
			2303 => "0000000111000100000100",
			2304 => "0000000010010000111101",
			2305 => "0011101111101000001100",
			2306 => "0001111111011100001000",
			2307 => "0011000100011000000100",
			2308 => "0000000010010000111101",
			2309 => "0000001010010000111101",
			2310 => "0000000010010000111101",
			2311 => "0011100110001100001000",
			2312 => "0010011010100100000100",
			2313 => "0000000010010000111101",
			2314 => "0000000010010000111101",
			2315 => "0010010010101100000100",
			2316 => "0000000010010000111101",
			2317 => "0000000010010000111101",
			2318 => "0000000010010000111101",
			2319 => "0010011010100000101100",
			2320 => "0001111111011100001000",
			2321 => "0001000110101100000100",
			2322 => "0000000010010011110001",
			2323 => "1111111010010011110001",
			2324 => "0010110010110100010100",
			2325 => "0001000011001100010000",
			2326 => "0011110000010000000100",
			2327 => "0000000010010011110001",
			2328 => "0010001100011100000100",
			2329 => "0000000010010011110001",
			2330 => "0001011100010100000100",
			2331 => "0000000010010011110001",
			2332 => "0000000010010011110001",
			2333 => "0000000010010011110001",
			2334 => "0011001111011100000100",
			2335 => "0000000010010011110001",
			2336 => "0010001011010100001000",
			2337 => "0001110010001000000100",
			2338 => "0000000010010011110001",
			2339 => "0000000010010011110001",
			2340 => "0000000010010011110001",
			2341 => "0011001001110100011100",
			2342 => "0000001000101100011000",
			2343 => "0001011100100100001000",
			2344 => "0011001010111000000100",
			2345 => "0000000010010011110001",
			2346 => "0000000010010011110001",
			2347 => "0011000100011000000100",
			2348 => "0000000010010011110001",
			2349 => "0000011101111100000100",
			2350 => "0000000010010011110001",
			2351 => "0010011010100000000100",
			2352 => "0000000010010011110001",
			2353 => "0000001010010011110001",
			2354 => "0000000010010011110001",
			2355 => "0000010100110100001100",
			2356 => "0001101000010000000100",
			2357 => "0000000010010011110001",
			2358 => "0001010111111100000100",
			2359 => "0000000010010011110001",
			2360 => "0000000010010011110001",
			2361 => "0010110101110100000100",
			2362 => "0000000010010011110001",
			2363 => "0000000010010011110001",
			2364 => "0011101110110100010000",
			2365 => "0001110110100100000100",
			2366 => "1111111010010101110101",
			2367 => "0001110110100100001000",
			2368 => "0011010001000000000100",
			2369 => "0000000010010101110101",
			2370 => "0000000010010101110101",
			2371 => "0000000010010101110101",
			2372 => "0011011111100100110000",
			2373 => "0011100110001100011100",
			2374 => "0010001001101000010100",
			2375 => "0010100011101000000100",
			2376 => "1111111010010101110101",
			2377 => "0000101000100000001000",
			2378 => "0001101001100100000100",
			2379 => "0000001010010101110101",
			2380 => "0000000010010101110101",
			2381 => "0000000111000000000100",
			2382 => "0000000010010101110101",
			2383 => "0000000010010101110101",
			2384 => "0011101100001100000100",
			2385 => "1111111010010101110101",
			2386 => "0000000010010101110101",
			2387 => "0010000111000100010000",
			2388 => "0001001001001100000100",
			2389 => "0000000010010101110101",
			2390 => "0000011010011000001000",
			2391 => "0011011100000000000100",
			2392 => "0000010010010101110101",
			2393 => "0000001010010101110101",
			2394 => "0000000010010101110101",
			2395 => "0000000010010101110101",
			2396 => "1111111010010101110101",
			2397 => "0000000010101000011000",
			2398 => "0000010001111000000100",
			2399 => "0000000010011000001001",
			2400 => "0001111000011000010000",
			2401 => "0000101000101000001100",
			2402 => "0010100011101000000100",
			2403 => "0000000010011000001001",
			2404 => "0011100110010000000100",
			2405 => "0000000010011000001001",
			2406 => "0000000010011000001001",
			2407 => "0000000010011000001001",
			2408 => "0000000010011000001001",
			2409 => "0001111111011100000100",
			2410 => "0000000010011000001001",
			2411 => "0001110101100100010000",
			2412 => "0010001011010100001100",
			2413 => "0010000001010100000100",
			2414 => "0000000010011000001001",
			2415 => "0000011100011000000100",
			2416 => "0000000010011000001001",
			2417 => "0000000010011000001001",
			2418 => "0000000010011000001001",
			2419 => "0011101000011100010000",
			2420 => "0001000110001100000100",
			2421 => "0000000010011000001001",
			2422 => "0001100101010000001000",
			2423 => "0011000001011000000100",
			2424 => "0000000010011000001001",
			2425 => "0000000010011000001001",
			2426 => "0000000010011000001001",
			2427 => "0011011011111000001100",
			2428 => "0001101001111100001000",
			2429 => "0001101000010000000100",
			2430 => "0000000010011000001001",
			2431 => "0000000010011000001001",
			2432 => "0000000010011000001001",
			2433 => "0000000010011000001001",
			2434 => "0001001011110000011100",
			2435 => "0011101011101100011000",
			2436 => "0001100100110100000100",
			2437 => "0000000010011010001101",
			2438 => "0010110110110100010000",
			2439 => "0010011010100000001100",
			2440 => "0000100110111100001000",
			2441 => "0000000110001000000100",
			2442 => "0000000010011010001101",
			2443 => "0000000010011010001101",
			2444 => "0000000010011010001101",
			2445 => "0000001010011010001101",
			2446 => "0000000010011010001101",
			2447 => "0000000010011010001101",
			2448 => "0001100100111100000100",
			2449 => "1111111010011010001101",
			2450 => "0010110001000000100000",
			2451 => "0001010111111100010000",
			2452 => "0001000110001100001100",
			2453 => "0010010010101100001000",
			2454 => "0011011110010000000100",
			2455 => "0000000010011010001101",
			2456 => "0000000010011010001101",
			2457 => "0000000010011010001101",
			2458 => "0000000010011010001101",
			2459 => "0001101001111100001100",
			2460 => "0010010010101100001000",
			2461 => "0000010101011100000100",
			2462 => "0000000010011010001101",
			2463 => "0000000010011010001101",
			2464 => "0000000010011010001101",
			2465 => "0000000010011010001101",
			2466 => "0000000010011010001101",
			2467 => "0011001000000000100000",
			2468 => "0000010001111000001000",
			2469 => "0011101111101000000100",
			2470 => "0000000010011100100001",
			2471 => "0000000010011100100001",
			2472 => "0010110110110100001000",
			2473 => "0010110100000100000100",
			2474 => "0000000010011100100001",
			2475 => "0000000010011100100001",
			2476 => "0010110100010000001100",
			2477 => "0000011100011000001000",
			2478 => "0001010111100000000100",
			2479 => "0000000010011100100001",
			2480 => "0000000010011100100001",
			2481 => "0000000010011100100001",
			2482 => "0000000010011100100001",
			2483 => "0001010110111100101000",
			2484 => "0000011010011000100100",
			2485 => "0000001111001000000100",
			2486 => "0000000010011100100001",
			2487 => "0001110101100100010000",
			2488 => "0001101000010000001000",
			2489 => "0001000011001100000100",
			2490 => "0000000010011100100001",
			2491 => "0000000010011100100001",
			2492 => "0010111010010100000100",
			2493 => "0000000010011100100001",
			2494 => "0000000010011100100001",
			2495 => "0011101000011100001000",
			2496 => "0001101000010000000100",
			2497 => "0000000010011100100001",
			2498 => "0000000010011100100001",
			2499 => "0001101001111100000100",
			2500 => "0000000010011100100001",
			2501 => "0000000010011100100001",
			2502 => "0000000010011100100001",
			2503 => "0000000010011100100001",
			2504 => "0010011010100000101100",
			2505 => "0011001011000000001000",
			2506 => "0001000110101100000100",
			2507 => "0000000010011111001101",
			2508 => "0000000010011111001101",
			2509 => "0000100010010100001100",
			2510 => "0010001000100100000100",
			2511 => "0000000010011111001101",
			2512 => "0001001000011100000100",
			2513 => "0000000010011111001101",
			2514 => "0000000010011111001101",
			2515 => "0011101011110000001000",
			2516 => "0011111000110100000100",
			2517 => "0000000010011111001101",
			2518 => "0000000010011111001101",
			2519 => "0000110100001100001100",
			2520 => "0011101000000100000100",
			2521 => "0000000010011111001101",
			2522 => "0011111111100000000100",
			2523 => "0000000010011111001101",
			2524 => "0000000010011111001101",
			2525 => "0000000010011111001101",
			2526 => "0011001011011100101000",
			2527 => "0010111011011100001000",
			2528 => "0001000011000000000100",
			2529 => "0000000010011111001101",
			2530 => "0000000010011111001101",
			2531 => "0001000110111000000100",
			2532 => "0000000010011111001101",
			2533 => "0011101111101000001100",
			2534 => "0001111111011100001000",
			2535 => "0011000100011000000100",
			2536 => "0000000010011111001101",
			2537 => "0000001010011111001101",
			2538 => "0000000010011111001101",
			2539 => "0011100110001100001000",
			2540 => "0000011100011000000100",
			2541 => "0000000010011111001101",
			2542 => "0000000010011111001101",
			2543 => "0000011100011000000100",
			2544 => "0000000010011111001101",
			2545 => "0000000010011111001101",
			2546 => "0000000010011111001101",
			2547 => "0011001101010100000100",
			2548 => "1111111010100001010001",
			2549 => "0011000001011000110100",
			2550 => "0000110011110000101000",
			2551 => "0001110001101000010000",
			2552 => "0000000010101000001100",
			2553 => "0010010000001000000100",
			2554 => "0000000010100001010001",
			2555 => "0000111100111000000100",
			2556 => "0000001010100001010001",
			2557 => "0000000010100001010001",
			2558 => "0000000010100001010001",
			2559 => "0001001010110100010000",
			2560 => "0001110111010000001000",
			2561 => "0010011010100100000100",
			2562 => "1111111010100001010001",
			2563 => "0000000010100001010001",
			2564 => "0010011010100100000100",
			2565 => "0000000010100001010001",
			2566 => "0000000010100001010001",
			2567 => "0011101000011100000100",
			2568 => "1111111010100001010001",
			2569 => "0000000010100001010001",
			2570 => "0010010010101100001000",
			2571 => "0000001011000100000100",
			2572 => "0000001010100001010001",
			2573 => "0000000010100001010001",
			2574 => "0000000010100001010001",
			2575 => "0001110100010000000100",
			2576 => "0000000010100001010001",
			2577 => "0010101010110000000100",
			2578 => "1111111010100001010001",
			2579 => "0000000010100001010001",
			2580 => "0010011010100000111100",
			2581 => "0001111111011100011000",
			2582 => "0001001111100100010100",
			2583 => "0010110100000100010000",
			2584 => "0001010001001000000100",
			2585 => "0000000010100100101101",
			2586 => "0000000001010100000100",
			2587 => "0000000010100100101101",
			2588 => "0001111000000000000100",
			2589 => "0000000010100100101101",
			2590 => "0000001010100100101101",
			2591 => "0000000010100100101101",
			2592 => "1111111010100100101101",
			2593 => "0011010111010100011100",
			2594 => "0001101000010000001100",
			2595 => "0001110101100100001000",
			2596 => "0001101001100100000100",
			2597 => "0000000010100100101101",
			2598 => "0000000010100100101101",
			2599 => "0000000010100100101101",
			2600 => "0001000011101100001000",
			2601 => "0001010111111100000100",
			2602 => "0000000010100100101101",
			2603 => "0000001010100100101101",
			2604 => "0010111101000100000100",
			2605 => "0000000010100100101101",
			2606 => "0000000010100100101101",
			2607 => "0001101001111100000100",
			2608 => "1111111010100100101101",
			2609 => "0000000010100100101101",
			2610 => "0000111101101100010000",
			2611 => "0000001010101100001100",
			2612 => "0010111011011100001000",
			2613 => "0010110000011100000100",
			2614 => "0000000010100100101101",
			2615 => "0000000010100100101101",
			2616 => "0000001010100100101101",
			2617 => "0000000010100100101101",
			2618 => "0000000010101000000100",
			2619 => "0000000010100100101101",
			2620 => "0000001101010000010100",
			2621 => "0010010010101100001100",
			2622 => "0011011010001000000100",
			2623 => "0000000010100100101101",
			2624 => "0001110101100100000100",
			2625 => "0000001010100100101101",
			2626 => "0000000010100100101101",
			2627 => "0011001000000000000100",
			2628 => "0000000010100100101101",
			2629 => "0000000010100100101101",
			2630 => "0000110011110000001000",
			2631 => "0000001101010000000100",
			2632 => "0000000010100100101101",
			2633 => "0000000010100100101101",
			2634 => "0000000010100100101101",
			2635 => "0010011010100000111100",
			2636 => "0001111111011100011000",
			2637 => "0001001111100100010100",
			2638 => "0010110100000100010000",
			2639 => "0001010001001000000100",
			2640 => "0000000010101000001001",
			2641 => "0000000001010100000100",
			2642 => "0000000010101000001001",
			2643 => "0001111000000000000100",
			2644 => "0000000010101000001001",
			2645 => "0000001010101000001001",
			2646 => "0000000010101000001001",
			2647 => "1111111010101000001001",
			2648 => "0011010111010100011100",
			2649 => "0001101000010000001100",
			2650 => "0001110101100100001000",
			2651 => "0001101001100100000100",
			2652 => "0000000010101000001001",
			2653 => "0000000010101000001001",
			2654 => "0000000010101000001001",
			2655 => "0001000011101100001000",
			2656 => "0001010111111100000100",
			2657 => "0000000010101000001001",
			2658 => "0000001010101000001001",
			2659 => "0010111101000100000100",
			2660 => "0000000010101000001001",
			2661 => "0000000010101000001001",
			2662 => "0001101001111100000100",
			2663 => "1111111010101000001001",
			2664 => "0000000010101000001001",
			2665 => "0001001011110000010000",
			2666 => "0000101101101100001100",
			2667 => "0001011100100100001000",
			2668 => "0001011101000100000100",
			2669 => "0000000010101000001001",
			2670 => "0000000010101000001001",
			2671 => "0000001010101000001001",
			2672 => "0000000010101000001001",
			2673 => "0010110010001000000100",
			2674 => "0000000010101000001001",
			2675 => "0000001101010000011000",
			2676 => "0000000010101000001000",
			2677 => "0001001011110000000100",
			2678 => "0000000010101000001001",
			2679 => "0000000010101000001001",
			2680 => "0011010010000100001000",
			2681 => "0000001101010000000100",
			2682 => "0000001010101000001001",
			2683 => "0000000010101000001001",
			2684 => "0011000001101000000100",
			2685 => "0000000010101000001001",
			2686 => "0000000010101000001001",
			2687 => "0000100011001100000100",
			2688 => "0000000010101000001001",
			2689 => "0000000010101000001001",
			2690 => "0000010101011100010100",
			2691 => "0000000111000000010000",
			2692 => "0000111000100000001100",
			2693 => "0011001011000000000100",
			2694 => "1111111010101010110101",
			2695 => "0011100111111100000100",
			2696 => "0000010010101010110101",
			2697 => "1111111010101010110101",
			2698 => "0000010010101010110101",
			2699 => "1111111010101010110101",
			2700 => "0010010010101100111100",
			2701 => "0001011001010000100000",
			2702 => "0001001011110000011100",
			2703 => "0010011010100000001100",
			2704 => "0000101100000000001000",
			2705 => "0000101100010000000100",
			2706 => "1111111010101010110101",
			2707 => "0000001010101010110101",
			2708 => "1111111010101010110101",
			2709 => "0000101111100100001000",
			2710 => "0001101001100100000100",
			2711 => "0000010010101010110101",
			2712 => "0000001010101010110101",
			2713 => "0010110010001000000100",
			2714 => "1111111010101010110101",
			2715 => "0000010010101010110101",
			2716 => "1111111010101010110101",
			2717 => "0010000101000100001000",
			2718 => "0010010101010000000100",
			2719 => "0000000010101010110101",
			2720 => "1111111010101010110101",
			2721 => "0000100110111000001000",
			2722 => "0000111111101000000100",
			2723 => "0000011010101010110101",
			2724 => "0000001010101010110101",
			2725 => "0011101000101000000100",
			2726 => "1111111010101010110101",
			2727 => "0010111110101000000100",
			2728 => "0000001010101010110101",
			2729 => "0000000010101010110101",
			2730 => "0000011100011000000100",
			2731 => "0000000010101010110101",
			2732 => "1111111010101010110101",
			2733 => "0010111010001100000100",
			2734 => "1111111010101100100001",
			2735 => "0011011111100100110000",
			2736 => "0011100110001100100000",
			2737 => "0000000010011000011100",
			2738 => "0010100011101000001100",
			2739 => "0010110100000100001000",
			2740 => "0001110110100100000100",
			2741 => "0000000010101100100001",
			2742 => "0000000010101100100001",
			2743 => "1111111010101100100001",
			2744 => "0001101001100100001000",
			2745 => "0000101000100000000100",
			2746 => "0000001010101100100001",
			2747 => "0000000010101100100001",
			2748 => "0011000100011000000100",
			2749 => "1111111010101100100001",
			2750 => "0000000010101100100001",
			2751 => "1111111010101100100001",
			2752 => "0010000111000100001100",
			2753 => "0001001001001100000100",
			2754 => "0000000010101100100001",
			2755 => "0000011010011000000100",
			2756 => "0000001010101100100001",
			2757 => "0000000010101100100001",
			2758 => "0000000010101100100001",
			2759 => "1111111010101100100001",
			2760 => "0000000001110100101100",
			2761 => "0011101011111000101000",
			2762 => "0010100011101000011000",
			2763 => "0010110111010000010000",
			2764 => "0010111010011100000100",
			2765 => "0000000010101111110101",
			2766 => "0001001000001100001000",
			2767 => "0001000010000100000100",
			2768 => "0000000010101111110101",
			2769 => "0000000010101111110101",
			2770 => "0000000010101111110101",
			2771 => "0010110100000100000100",
			2772 => "0000000010101111110101",
			2773 => "0000000010101111110101",
			2774 => "0011101110110100000100",
			2775 => "0000000010101111110101",
			2776 => "0011011100100100000100",
			2777 => "0000000010101111110101",
			2778 => "0001000010010100000100",
			2779 => "0000001010101111110101",
			2780 => "0000000010101111110101",
			2781 => "0000000010101111110101",
			2782 => "0011101000101000010000",
			2783 => "0010010010101100001000",
			2784 => "0000011010011000000100",
			2785 => "1111111010101111110101",
			2786 => "0000000010101111110101",
			2787 => "0000011010011000000100",
			2788 => "0000000010101111110101",
			2789 => "0000000010101111110101",
			2790 => "0000000111000000001000",
			2791 => "0000101110000000000100",
			2792 => "1111111010101111110101",
			2793 => "0000000010101111110101",
			2794 => "0000101110000000001100",
			2795 => "0011011010001000000100",
			2796 => "0000000010101111110101",
			2797 => "0011011001100000000100",
			2798 => "0000001010101111110101",
			2799 => "0000000010101111110101",
			2800 => "0010110010110100010000",
			2801 => "0011001000011000001000",
			2802 => "0011010010000100000100",
			2803 => "0000000010101111110101",
			2804 => "0000000010101111110101",
			2805 => "0001101000010000000100",
			2806 => "0000000010101111110101",
			2807 => "0000000010101111110101",
			2808 => "0011001111011100000100",
			2809 => "0000000010101111110101",
			2810 => "0011111001001100000100",
			2811 => "0000000010101111110101",
			2812 => "0000000010101111110101",
			2813 => "0000010101011100010100",
			2814 => "0000000111000100010000",
			2815 => "0000111000100000001100",
			2816 => "0000011101101000001000",
			2817 => "0001110100001000000100",
			2818 => "1111111010110010011001",
			2819 => "0000010010110010011001",
			2820 => "1111111010110010011001",
			2821 => "0000010010110010011001",
			2822 => "1111111010110010011001",
			2823 => "0000011010011000111100",
			2824 => "0001011001010000011100",
			2825 => "0001001011110000011000",
			2826 => "0000011101111100001100",
			2827 => "0000101100000000001000",
			2828 => "0000101100010000000100",
			2829 => "1111111010110010011001",
			2830 => "0000001010110010011001",
			2831 => "1111111010110010011001",
			2832 => "0000111100111000001000",
			2833 => "0000001010101100000100",
			2834 => "0000001010110010011001",
			2835 => "1111111010110010011001",
			2836 => "1111111010110010011001",
			2837 => "1111111010110010011001",
			2838 => "0010000101000100001000",
			2839 => "0000010001000100000100",
			2840 => "0000000010110010011001",
			2841 => "1111111010110010011001",
			2842 => "0011010111010100001100",
			2843 => "0000101111101000000100",
			2844 => "0000011010110010011001",
			2845 => "0010101000010100000100",
			2846 => "1111111010110010011001",
			2847 => "0000001010110010011001",
			2848 => "0001101001111100000100",
			2849 => "1111110010110010011001",
			2850 => "0010001011010100000100",
			2851 => "0000000010110010011001",
			2852 => "0000001010110010011001",
			2853 => "1111111010110010011001",
			2854 => "0010011000010000011100",
			2855 => "0000000111000000011000",
			2856 => "0000000001010100000100",
			2857 => "1111111010110101010101",
			2858 => "0000000001010100000100",
			2859 => "0000000010110101010101",
			2860 => "0000000111000000001100",
			2861 => "0000000110001000000100",
			2862 => "1111111010110101010101",
			2863 => "0000001111001000000100",
			2864 => "0000011010110101010101",
			2865 => "1111111010110101010101",
			2866 => "0000000010110101010101",
			2867 => "1111111010110101010101",
			2868 => "0010010010101100111100",
			2869 => "0011011110010000011100",
			2870 => "0010011010100100010100",
			2871 => "0000101100000000001000",
			2872 => "0010100011101000000100",
			2873 => "1111111010110101010101",
			2874 => "0001100010110101010101",
			2875 => "0001000010010100001000",
			2876 => "0000000111000100000100",
			2877 => "1111111010110101010101",
			2878 => "0000011010110101010101",
			2879 => "1111111010110101010101",
			2880 => "0010101000010100000100",
			2881 => "0000010010110101010101",
			2882 => "1111111010110101010101",
			2883 => "0001100100111100001100",
			2884 => "0001010010011100000100",
			2885 => "0000010010110101010101",
			2886 => "0000000111000000000100",
			2887 => "1111111010110101010101",
			2888 => "1111110010110101010101",
			2889 => "0000101110000000000100",
			2890 => "0000110010110101010101",
			2891 => "0010011010100000001000",
			2892 => "0011010111010100000100",
			2893 => "0000001010110101010101",
			2894 => "0000000010110101010101",
			2895 => "0001001110111000000100",
			2896 => "0000011010110101010101",
			2897 => "0000001010110101010101",
			2898 => "0000110001011100000100",
			2899 => "0000010010110101010101",
			2900 => "1111111010110101010101",
			2901 => "0011001010111000001000",
			2902 => "0000011100011000000100",
			2903 => "1111111010111000010001",
			2904 => "0000000010111000010001",
			2905 => "0001000011001100111100",
			2906 => "0010000101000100100000",
			2907 => "0001011110101100001100",
			2908 => "0001000110101100001000",
			2909 => "0000101010001000000100",
			2910 => "0000000010111000010001",
			2911 => "0000001010111000010001",
			2912 => "0000000010111000010001",
			2913 => "0011010011001000001100",
			2914 => "0010011010100100001000",
			2915 => "0010110100000100000100",
			2916 => "0000000010111000010001",
			2917 => "1111111010111000010001",
			2918 => "0000000010111000010001",
			2919 => "0010111011110100000100",
			2920 => "0000000010111000010001",
			2921 => "0000000010111000010001",
			2922 => "0011010110010000010000",
			2923 => "0010111011011100000100",
			2924 => "0000000010111000010001",
			2925 => "0010001100000100001000",
			2926 => "0011000100011000000100",
			2927 => "0000000010111000010001",
			2928 => "0000001010111000010001",
			2929 => "0000000010111000010001",
			2930 => "0001101000010000000100",
			2931 => "0000000010111000010001",
			2932 => "0000011100011000000100",
			2933 => "0000000010111000010001",
			2934 => "0000000010111000010001",
			2935 => "0011101000000100000100",
			2936 => "1111111010111000010001",
			2937 => "0001011100010000010000",
			2938 => "0011011001100000000100",
			2939 => "0000000010111000010001",
			2940 => "0000011100011000001000",
			2941 => "0000011011111100000100",
			2942 => "0000000010111000010001",
			2943 => "0000001010111000010001",
			2944 => "0000000010111000010001",
			2945 => "0001101001111100000100",
			2946 => "1111111010111000010001",
			2947 => "0000000010111000010001",
			2948 => "0011001101010100000100",
			2949 => "1111111010111010100101",
			2950 => "0011000001011000111100",
			2951 => "0001110001101000010100",
			2952 => "0000000010101000010000",
			2953 => "0010010000001000000100",
			2954 => "0000000010111010100101",
			2955 => "0011001000000000001000",
			2956 => "0001001011110000000100",
			2957 => "0000001010111010100101",
			2958 => "0000000010111010100101",
			2959 => "0000000010111010100101",
			2960 => "0000000010111010100101",
			2961 => "0011101000110100011000",
			2962 => "0001000011001100010000",
			2963 => "0000000111000000001000",
			2964 => "0000011001011000000100",
			2965 => "0000000010111010100101",
			2966 => "0000000010111010100101",
			2967 => "0010111011110100000100",
			2968 => "0000000010111010100101",
			2969 => "0000000010111010100101",
			2970 => "0011101000000100000100",
			2971 => "1111111010111010100101",
			2972 => "0000000010111010100101",
			2973 => "0010110000110100000100",
			2974 => "0000000010111010100101",
			2975 => "0010010010101100001000",
			2976 => "0000000100000000000100",
			2977 => "0000001010111010100101",
			2978 => "0000000010111010100101",
			2979 => "0000000010111010100101",
			2980 => "0001110100010000000100",
			2981 => "0000000010111010100101",
			2982 => "0001101001111100000100",
			2983 => "1111111010111010100101",
			2984 => "0000000010111010100101",
			2985 => "0000011101011100000100",
			2986 => "1111111010111100100001",
			2987 => "0010010010101100110100",
			2988 => "0000001011010100000100",
			2989 => "1111111010111100100001",
			2990 => "0001001011110000011000",
			2991 => "0001011100100100001100",
			2992 => "0001001111100100000100",
			2993 => "0000001010111100100001",
			2994 => "0000010100110100000100",
			2995 => "1111111010111100100001",
			2996 => "0000000010111100100001",
			2997 => "0011101011101100001000",
			2998 => "0000000110001000000100",
			2999 => "0000000010111100100001",
			3000 => "0000010010111100100001",
			3001 => "0000000010111100100001",
			3002 => "0011101100001100001100",
			3003 => "0001001001001100001000",
			3004 => "0010110010001000000100",
			3005 => "1111111010111100100001",
			3006 => "0000000010111100100001",
			3007 => "1111111010111100100001",
			3008 => "0010001001101000000100",
			3009 => "0000000010111100100001",
			3010 => "0010011010100000000100",
			3011 => "0000001010111100100001",
			3012 => "0000010010111100100001",
			3013 => "0001001011110000000100",
			3014 => "0000000010111100100001",
			3015 => "1111111010111100100001",
			3016 => "0011001101010100000100",
			3017 => "1111111010111111101101",
			3018 => "0010011010100000101100",
			3019 => "0011101000011100011000",
			3020 => "0010010101010000010000",
			3021 => "0001000011110000001100",
			3022 => "0001100100110100000100",
			3023 => "0000000010111111101101",
			3024 => "0011000100011000000100",
			3025 => "0000000010111111101101",
			3026 => "0000000010111111101101",
			3027 => "0000000010111111101101",
			3028 => "0011101011110000000100",
			3029 => "1111111010111111101101",
			3030 => "0000000010111111101101",
			3031 => "0000111110111000001100",
			3032 => "0000111110100100000100",
			3033 => "0000000010111111101101",
			3034 => "0000001011000100000100",
			3035 => "0000001010111111101101",
			3036 => "0000000010111111101101",
			3037 => "0001011100000000000100",
			3038 => "0000000010111111101101",
			3039 => "0000000010111111101101",
			3040 => "0011001000000000010100",
			3041 => "0010011010100100001000",
			3042 => "0001101111000000000100",
			3043 => "0000000010111111101101",
			3044 => "0000000010111111101101",
			3045 => "0000001000101100001000",
			3046 => "0010111011011100000100",
			3047 => "0000000010111111101101",
			3048 => "0000001010111111101101",
			3049 => "0000000010111111101101",
			3050 => "0010000001110000001100",
			3051 => "0010011010100100001000",
			3052 => "0010011010100100000100",
			3053 => "0000000010111111101101",
			3054 => "0000000010111111101101",
			3055 => "1111111010111111101101",
			3056 => "0001010011001000001100",
			3057 => "0010001100000100001000",
			3058 => "0010011010100100000100",
			3059 => "0000000010111111101101",
			3060 => "0000000010111111101101",
			3061 => "0000000010111111101101",
			3062 => "0011101110000000000100",
			3063 => "0000000010111111101101",
			3064 => "0010010010101100000100",
			3065 => "0000001010111111101101",
			3066 => "0000000010111111101101",
			3067 => "0001010001001000000100",
			3068 => "1111111011000010000001",
			3069 => "0000111100111000100000",
			3070 => "0010100011101000001000",
			3071 => "0000011111001100000100",
			3072 => "0000001011000010000001",
			3073 => "1111111011000010000001",
			3074 => "0000000010101000010100",
			3075 => "0001011100100100001100",
			3076 => "0001001111100100000100",
			3077 => "0000001011000010000001",
			3078 => "0010011010100100000100",
			3079 => "1111111011000010000001",
			3080 => "0000000011000010000001",
			3081 => "0001000001011100000100",
			3082 => "0000000011000010000001",
			3083 => "0000001011000010000001",
			3084 => "0000000011000010000001",
			3085 => "0000000010101000000100",
			3086 => "1111111011000010000001",
			3087 => "0010110010001000000100",
			3088 => "1111111011000010000001",
			3089 => "0011001000011000010000",
			3090 => "0000011100011000001000",
			3091 => "0001011001010000000100",
			3092 => "1111111011000010000001",
			3093 => "0000000011000010000001",
			3094 => "0010001001101000000100",
			3095 => "0000001011000010000001",
			3096 => "0000000011000010000001",
			3097 => "0010101001000100001000",
			3098 => "0001110000011100000100",
			3099 => "0000000011000010000001",
			3100 => "1111111011000010000001",
			3101 => "0011011111100100000100",
			3102 => "0000000011000010000001",
			3103 => "1111111011000010000001",
			3104 => "0000011101111101001000",
			3105 => "0011000100011000001000",
			3106 => "0000110010010100000100",
			3107 => "1111111011000110001101",
			3108 => "0000000011000110001101",
			3109 => "0000000111000000011100",
			3110 => "0001101001100100001100",
			3111 => "0000101010001000001000",
			3112 => "0011010001000000000100",
			3113 => "0000000011000110001101",
			3114 => "0000000011000110001101",
			3115 => "0000000011000110001101",
			3116 => "0010110110110100000100",
			3117 => "0000000011000110001101",
			3118 => "0001010111111100001000",
			3119 => "0000010001111000000100",
			3120 => "0000001011000110001101",
			3121 => "0000000011000110001101",
			3122 => "0000000011000110001101",
			3123 => "0011101000011100010000",
			3124 => "0010011001111100001100",
			3125 => "0010011000010000000100",
			3126 => "1111111011000110001101",
			3127 => "0010010101010000000100",
			3128 => "0000000011000110001101",
			3129 => "0000000011000110001101",
			3130 => "1111111011000110001101",
			3131 => "0010110111100000001100",
			3132 => "0000111110100100000100",
			3133 => "0000000011000110001101",
			3134 => "0000001100001000000100",
			3135 => "0000001011000110001101",
			3136 => "0000000011000110001101",
			3137 => "0011011111100100000100",
			3138 => "0000000011000110001101",
			3139 => "0000000011000110001101",
			3140 => "0011001000011000110100",
			3141 => "0011010111111100010000",
			3142 => "0000111111100100001100",
			3143 => "0010011010100000000100",
			3144 => "0000000011000110001101",
			3145 => "0000000001110100000100",
			3146 => "0000001011000110001101",
			3147 => "0000000011000110001101",
			3148 => "1111111011000110001101",
			3149 => "0001011110000100001000",
			3150 => "0010011010100100000100",
			3151 => "0000000011000110001101",
			3152 => "0000001011000110001101",
			3153 => "0000000111000000001100",
			3154 => "0000110001011100001000",
			3155 => "0010101000100100000100",
			3156 => "0000000011000110001101",
			3157 => "0000001011000110001101",
			3158 => "1111111011000110001101",
			3159 => "0010001001101000001000",
			3160 => "0001011001010000000100",
			3161 => "0000000011000110001101",
			3162 => "0000001011000110001101",
			3163 => "0000100011001100000100",
			3164 => "0000000011000110001101",
			3165 => "0000000011000110001101",
			3166 => "0000010100110100000100",
			3167 => "0000000011000110001101",
			3168 => "0011100010111000000100",
			3169 => "1111111011000110001101",
			3170 => "0000000011000110001101",
			3171 => "0011001101010100000100",
			3172 => "1111111011001001001001",
			3173 => "0010011010100101001000",
			3174 => "0010110111010000010100",
			3175 => "0000000110001000010000",
			3176 => "0001100100110100000100",
			3177 => "0000000011001001001001",
			3178 => "0001001111100100001000",
			3179 => "0001110011100000000100",
			3180 => "0000000011001001001001",
			3181 => "0000001011001001001001",
			3182 => "0000000011001001001001",
			3183 => "0000000011001001001001",
			3184 => "0010110110110100011000",
			3185 => "0010110100000100001100",
			3186 => "0001001111100100001000",
			3187 => "0010010111101100000100",
			3188 => "0000000011001001001001",
			3189 => "0000000011001001001001",
			3190 => "0000000011001001001001",
			3191 => "0001011100100100000100",
			3192 => "1111111011001001001001",
			3193 => "0001010111100000000100",
			3194 => "0000000011001001001001",
			3195 => "0000000011001001001001",
			3196 => "0000001000101100001100",
			3197 => "0001101001100100000100",
			3198 => "0000000011001001001001",
			3199 => "0000010001111000000100",
			3200 => "0000001011001001001001",
			3201 => "0000000011001001001001",
			3202 => "0011101011110000001000",
			3203 => "0000001000110000000100",
			3204 => "0000000011001001001001",
			3205 => "1111111011001001001001",
			3206 => "0011011111100100000100",
			3207 => "0000000011001001001001",
			3208 => "1111111011001001001001",
			3209 => "0011001000000000010000",
			3210 => "0011001011000000001000",
			3211 => "0010110101100100000100",
			3212 => "0000000011001001001001",
			3213 => "0000000011001001001001",
			3214 => "0000001101010000000100",
			3215 => "0000001011001001001001",
			3216 => "0000000011001001001001",
			3217 => "1111111011001001001001",
			3218 => "0011001010111000001000",
			3219 => "0000011100011000000100",
			3220 => "1111111011001011110101",
			3221 => "0000000011001011110101",
			3222 => "0011011111100101001100",
			3223 => "0011100101000000111100",
			3224 => "0000101110000000100000",
			3225 => "0000000111000000010000",
			3226 => "0011101101101100001000",
			3227 => "0001001111101000000100",
			3228 => "0000000011001011110101",
			3229 => "0000001011001011110101",
			3230 => "0000011101111100000100",
			3231 => "0000000011001011110101",
			3232 => "1111111011001011110101",
			3233 => "0010011010100100001000",
			3234 => "0001110111010000000100",
			3235 => "1111111011001011110101",
			3236 => "0000000011001011110101",
			3237 => "0011000001101000000100",
			3238 => "0000001011001011110101",
			3239 => "0000000011001011110101",
			3240 => "0011101011110000010000",
			3241 => "0000101000110100001000",
			3242 => "0000010111101000000100",
			3243 => "0000000011001011110101",
			3244 => "0000000011001011110101",
			3245 => "0010101001000100000100",
			3246 => "0000000011001011110101",
			3247 => "1111111011001011110101",
			3248 => "0010001100000100000100",
			3249 => "1111111011001011110101",
			3250 => "0010001001101000000100",
			3251 => "0000001011001011110101",
			3252 => "1111111011001011110101",
			3253 => "0000011100011000001100",
			3254 => "0000001011000100001000",
			3255 => "0001010011001000000100",
			3256 => "0000000011001011110101",
			3257 => "0000001011001011110101",
			3258 => "0000000011001011110101",
			3259 => "0000000011001011110101",
			3260 => "1111111011001011110101",
			3261 => "0011101110110100000100",
			3262 => "1111111011001110010011",
			3263 => "0011011111100101001000",
			3264 => "0011101100001100110100",
			3265 => "0001110101100100011100",
			3266 => "0010001100000100001100",
			3267 => "0001101011001100000100",
			3268 => "1111111011001110010011",
			3269 => "0001101111000000000100",
			3270 => "0000001011001110010011",
			3271 => "0000001011001110010011",
			3272 => "0011011001100000001000",
			3273 => "0010111010010100000100",
			3274 => "1111111011001110010011",
			3275 => "0000000011001110010011",
			3276 => "0001001010110100000100",
			3277 => "0000001011001110010011",
			3278 => "0000000011001110010011",
			3279 => "0011101000011100001100",
			3280 => "0001001101001000001000",
			3281 => "0010000001110000000100",
			3282 => "1111111011001110010011",
			3283 => "0000000011001110010011",
			3284 => "1111111011001110010011",
			3285 => "0000001000110000000100",
			3286 => "0000000011001110010011",
			3287 => "0000000010011000000100",
			3288 => "0000001011001110010011",
			3289 => "0000000011001110010011",
			3290 => "0010000111000100010000",
			3291 => "0001010011001000000100",
			3292 => "0000000011001110010011",
			3293 => "0001110101100100000100",
			3294 => "0000011011001110010011",
			3295 => "0010001100000100000100",
			3296 => "0000000011001110010011",
			3297 => "0000001011001110010011",
			3298 => "0000000011001110010011",
			3299 => "1111111011001110010011",
			3300 => "0000000011001110010101",
			3301 => "0000000011001110011001",
			3302 => "0000000011001110011101",
			3303 => "0000000011001110100001",
			3304 => "0000000011001110100101",
			3305 => "0000000011001110101001",
			3306 => "0000000011001110101101",
			3307 => "0000000011001110110001",
			3308 => "0000000011001110110101",
			3309 => "0000000011001110111001",
			3310 => "0000000011001110111101",
			3311 => "0000000011001111000001",
			3312 => "0000000011001111000101",
			3313 => "0000000011001111001001",
			3314 => "0000000011001111001101",
			3315 => "0000000011001111010001",
			3316 => "0000000011001111010101",
			3317 => "0000000011001111011001",
			3318 => "0000000011001111011101",
			3319 => "0010011010100100000100",
			3320 => "0000000011001111101001",
			3321 => "0000000011001111101001",
			3322 => "0001100100111100000100",
			3323 => "0000000011001111111101",
			3324 => "0001101001111100000100",
			3325 => "0000000011001111111101",
			3326 => "0000000011001111111101",
			3327 => "0000010100110100001000",
			3328 => "0000010111101000000100",
			3329 => "0000000011010000010001",
			3330 => "0000000011010000010001",
			3331 => "0000000011010000010001",
			3332 => "0000011100011000001000",
			3333 => "0000000001110000000100",
			3334 => "0000000011010000100101",
			3335 => "0000000011010000100101",
			3336 => "0000000011010000100101",
			3337 => "0010011010100100001000",
			3338 => "0001101001111100000100",
			3339 => "0000000011010000111001",
			3340 => "0000000011010000111001",
			3341 => "0000000011010000111001",
			3342 => "0001111111011100001000",
			3343 => "0001110001101000000100",
			3344 => "0000000011010001010101",
			3345 => "0000000011010001010101",
			3346 => "0001110100010000000100",
			3347 => "0000000011010001010101",
			3348 => "0000000011010001010101",
			3349 => "0000000010101000001100",
			3350 => "0010001010110000000100",
			3351 => "0000000011010001110001",
			3352 => "0010000001010100000100",
			3353 => "0000000011010001110001",
			3354 => "0000000011010001110001",
			3355 => "0000000011010001110001",
			3356 => "0001001000011100000100",
			3357 => "0000000011010010001101",
			3358 => "0000100011110100001000",
			3359 => "0000010111101000000100",
			3360 => "0000000011010010001101",
			3361 => "0000000011010010001101",
			3362 => "0000000011010010001101",
			3363 => "0010011010100000000100",
			3364 => "0000000011010010101001",
			3365 => "0001010111011000001000",
			3366 => "0010010011101000000100",
			3367 => "0000000011010010101001",
			3368 => "0000000011010010101001",
			3369 => "0000000011010010101001",
			3370 => "0000000010101000001100",
			3371 => "0010011010100100000100",
			3372 => "0000000011010011010101",
			3373 => "0011110011000000000100",
			3374 => "0000000011010011010101",
			3375 => "0000000011010011010101",
			3376 => "0000111000110100001000",
			3377 => "0000001010101100000100",
			3378 => "0000000011010011010101",
			3379 => "0000000011010011010101",
			3380 => "0000000011010011010101",
			3381 => "0010111011011100000100",
			3382 => "0000000011010011111001",
			3383 => "0001101001111100001100",
			3384 => "0001100100111100000100",
			3385 => "0000000011010011111001",
			3386 => "0010110110100000000100",
			3387 => "0000000011010011111001",
			3388 => "0000000011010011111001",
			3389 => "0000000011010011111001",
			3390 => "0010011010100000000100",
			3391 => "0000000011010100011101",
			3392 => "0010110010110100001100",
			3393 => "0010010011101000001000",
			3394 => "0010011010100000000100",
			3395 => "0000000011010100011101",
			3396 => "0000000011010100011101",
			3397 => "0000000011010100011101",
			3398 => "0000000011010100011101",
			3399 => "0000001000101100010000",
			3400 => "0010100011101000000100",
			3401 => "0000000011010101001001",
			3402 => "0001010011001000001000",
			3403 => "0001011100100100000100",
			3404 => "0000000011010101001001",
			3405 => "0000000011010101001001",
			3406 => "0000000011010101001001",
			3407 => "0000100011110100000100",
			3408 => "0000000011010101001001",
			3409 => "0000000011010101001001",
			3410 => "0010010111101100000100",
			3411 => "0000000011010101110101",
			3412 => "0000010100110100001000",
			3413 => "0010001010110000000100",
			3414 => "0000000011010101110101",
			3415 => "0000000011010101110101",
			3416 => "0000111011101100000100",
			3417 => "0000000011010101110101",
			3418 => "0000110011110000000100",
			3419 => "0000000011010101110101",
			3420 => "0000000011010101110101",
			3421 => "0010011010100100010100",
			3422 => "0001110111010000001000",
			3423 => "0001001111100100000100",
			3424 => "0000000011010110110001",
			3425 => "0000000011010110110001",
			3426 => "0001110100010000001000",
			3427 => "0010111011110100000100",
			3428 => "0000000011010110110001",
			3429 => "0000000011010110110001",
			3430 => "0000000011010110110001",
			3431 => "0001111111011100001000",
			3432 => "0010010011101000000100",
			3433 => "0000000011010110110001",
			3434 => "0000000011010110110001",
			3435 => "0000000011010110110001",
			3436 => "0000001101010000010100",
			3437 => "0010100011101000000100",
			3438 => "0000000011010111011101",
			3439 => "0010011010100100001100",
			3440 => "0010011010011000000100",
			3441 => "0000000011010111011101",
			3442 => "0000001011010100000100",
			3443 => "0000000011010111011101",
			3444 => "0000000011010111011101",
			3445 => "0000000011010111011101",
			3446 => "0000000011010111011101",
			3447 => "0010000001010100001100",
			3448 => "0010011010100100000100",
			3449 => "0000000011011000100001",
			3450 => "0000100001011100000100",
			3451 => "0000000011011000100001",
			3452 => "0000000011011000100001",
			3453 => "0011101110000000001100",
			3454 => "0000011100011000001000",
			3455 => "0001000110111000000100",
			3456 => "0000000011011000100001",
			3457 => "0000000011011000100001",
			3458 => "0000000011011000100001",
			3459 => "0011011111100100001000",
			3460 => "0001110111010000000100",
			3461 => "0000000011011000100001",
			3462 => "0000000011011000100001",
			3463 => "0000000011011000100001",
			3464 => "0010000001010100010000",
			3465 => "0001011100100100000100",
			3466 => "0000000011011001100101",
			3467 => "0000001111001000000100",
			3468 => "0000000011011001100101",
			3469 => "0001010010011100000100",
			3470 => "0000000011011001100101",
			3471 => "0000000011011001100101",
			3472 => "0011101110000000010000",
			3473 => "0000011100011000001100",
			3474 => "0001001000110100000100",
			3475 => "0000000011011001100101",
			3476 => "0010011001111100000100",
			3477 => "0000000011011001100101",
			3478 => "0000000011011001100101",
			3479 => "0000000011011001100101",
			3480 => "0000000011011001100101",
			3481 => "0010010111101100010000",
			3482 => "0001110111010000001100",
			3483 => "0011101000101000001000",
			3484 => "0001100100110100000100",
			3485 => "0000000011011010111001",
			3486 => "0000000011011010111001",
			3487 => "0000000011011010111001",
			3488 => "0000000011011010111001",
			3489 => "0000010100110100001100",
			3490 => "0010100011101000000100",
			3491 => "0000000011011010111001",
			3492 => "0011100110010000000100",
			3493 => "0000000011011010111001",
			3494 => "0000000011011010111001",
			3495 => "0000111011101100000100",
			3496 => "0000000011011010111001",
			3497 => "0000110011110000001000",
			3498 => "0011001000000000000100",
			3499 => "0000000011011010111001",
			3500 => "0000000011011010111001",
			3501 => "0000000011011010111001",
			3502 => "0001001011110000011000",
			3503 => "0011101011101100010100",
			3504 => "0011011110101100000100",
			3505 => "0000000011011011110101",
			3506 => "0010001000100100000100",
			3507 => "0000000011011011110101",
			3508 => "0011011100010100001000",
			3509 => "0000001010101100000100",
			3510 => "0000000011011011110101",
			3511 => "0000000011011011110101",
			3512 => "0000000011011011110101",
			3513 => "0000000011011011110101",
			3514 => "0011100010010100000100",
			3515 => "0000000011011011110101",
			3516 => "0000000011011011110101",
			3517 => "0010110101110100011000",
			3518 => "0010000001110000010100",
			3519 => "0010111011011100000100",
			3520 => "0000000011011101000001",
			3521 => "0011111111100100000100",
			3522 => "0000000011011101000001",
			3523 => "0011000100011000000100",
			3524 => "0000000011011101000001",
			3525 => "0001001000101000000100",
			3526 => "0000000011011101000001",
			3527 => "0000000011011101000001",
			3528 => "0000000011011101000001",
			3529 => "0010000001110000001000",
			3530 => "0011100110111100000100",
			3531 => "0000000011011101000001",
			3532 => "0000000011011101000001",
			3533 => "0010001011010100000100",
			3534 => "0000000011011101000001",
			3535 => "0000000011011101000001",
			3536 => "0001011001010000000100",
			3537 => "0000000011011101110101",
			3538 => "0011011011111000010100",
			3539 => "0010010010101100010000",
			3540 => "0000000010101000000100",
			3541 => "0000000011011101110101",
			3542 => "0011101100111000000100",
			3543 => "0000000011011101110101",
			3544 => "0010000111000100000100",
			3545 => "0000000011011101110101",
			3546 => "0000000011011101110101",
			3547 => "0000000011011101110101",
			3548 => "0000000011011101110101",
			3549 => "0010011010100000000100",
			3550 => "0000000011011110101001",
			3551 => "0001110101100100010100",
			3552 => "0001001001001100010000",
			3553 => "0010011010100000000100",
			3554 => "0000000011011110101001",
			3555 => "0010010011101000001000",
			3556 => "0001011100010100000100",
			3557 => "0000000011011110101001",
			3558 => "0000000011011110101001",
			3559 => "0000000011011110101001",
			3560 => "0000000011011110101001",
			3561 => "0000000011011110101001",
			3562 => "0001001011110000011000",
			3563 => "0000111101101100010100",
			3564 => "0010001010110000000100",
			3565 => "0000000011011111110101",
			3566 => "0010000001010100001100",
			3567 => "0010111011011100000100",
			3568 => "0000000011011111110101",
			3569 => "0000111000001100000100",
			3570 => "0000000011011111110101",
			3571 => "0000000011011111110101",
			3572 => "0000000011011111110101",
			3573 => "0000000011011111110101",
			3574 => "0000111000000100000100",
			3575 => "0000000011011111110101",
			3576 => "0010111001010000001000",
			3577 => "0010111011110100000100",
			3578 => "0000000011011111110101",
			3579 => "0000000011011111110101",
			3580 => "0000000011011111110101",
			3581 => "0010000110011100010100",
			3582 => "0010100011101000000100",
			3583 => "0000000011100001011001",
			3584 => "0010100111110100001100",
			3585 => "0001101111000000001000",
			3586 => "0001101011001100000100",
			3587 => "0000000011100001011001",
			3588 => "0000000011100001011001",
			3589 => "0000000011100001011001",
			3590 => "0000000011100001011001",
			3591 => "0001101000010000001000",
			3592 => "0000011100011000000100",
			3593 => "0000000011100001011001",
			3594 => "0000000011100001011001",
			3595 => "0000001101010000001100",
			3596 => "0000100110111000000100",
			3597 => "0000000011100001011001",
			3598 => "0010000001110000000100",
			3599 => "0000000011100001011001",
			3600 => "0000000011100001011001",
			3601 => "0000000011111100001000",
			3602 => "0010101100011100000100",
			3603 => "0000000011100001011001",
			3604 => "0000000011100001011001",
			3605 => "0000000011100001011001",
			3606 => "0001100100111100001100",
			3607 => "0001001011101100000100",
			3608 => "0000000011100010100101",
			3609 => "0010010010101100000100",
			3610 => "0000000011100010100101",
			3611 => "0000000011100010100101",
			3612 => "0011000001011000011000",
			3613 => "0000000010101000000100",
			3614 => "0000000011100010100101",
			3615 => "0000000010111100010000",
			3616 => "0010110010001000000100",
			3617 => "0000000011100010100101",
			3618 => "0010010010101100001000",
			3619 => "0011010111111100000100",
			3620 => "0000000011100010100101",
			3621 => "0000000011100010100101",
			3622 => "0000000011100010100101",
			3623 => "0000000011100010100101",
			3624 => "0000000011100010100101",
			3625 => "0011001011000000001000",
			3626 => "0011110110111000000100",
			3627 => "0000000011100011101001",
			3628 => "0000000011100011101001",
			3629 => "0011011111100100011000",
			3630 => "0010110010001000000100",
			3631 => "0000000011100011101001",
			3632 => "0001001011110000000100",
			3633 => "0000000011100011101001",
			3634 => "0001110100010000001100",
			3635 => "0001001001001100001000",
			3636 => "0011011010001000000100",
			3637 => "0000000011100011101001",
			3638 => "0000000011100011101001",
			3639 => "0000000011100011101001",
			3640 => "0000000011100011101001",
			3641 => "0000000011100011101001",
			3642 => "0010011010100100010100",
			3643 => "0011001000000000001000",
			3644 => "0000000001110100000100",
			3645 => "0000000011100101000101",
			3646 => "0000000011100101000101",
			3647 => "0011000010001000001000",
			3648 => "0001001001000000000100",
			3649 => "0000000011100101000101",
			3650 => "0000000011100101000101",
			3651 => "0000000011100101000101",
			3652 => "0011001000011000011000",
			3653 => "0010010011101000010100",
			3654 => "0000000010101000000100",
			3655 => "0000000011100101000101",
			3656 => "0011000100011000000100",
			3657 => "0000000011100101000101",
			3658 => "0010001001101000001000",
			3659 => "0010000101000100000100",
			3660 => "0000000011100101000101",
			3661 => "0000000011100101000101",
			3662 => "0000000011100101000101",
			3663 => "0000000011100101000101",
			3664 => "0000000011100101000101",
			3665 => "0011101011111000011000",
			3666 => "0000000001110100010100",
			3667 => "0001100100110100000100",
			3668 => "0000000011100110110001",
			3669 => "0001010101110000001100",
			3670 => "0011001101010100000100",
			3671 => "0000000011100110110001",
			3672 => "0010001000100100000100",
			3673 => "0000000011100110110001",
			3674 => "0000000011100110110001",
			3675 => "0000000011100110110001",
			3676 => "0000000011100110110001",
			3677 => "0011000001101000001100",
			3678 => "0000100110111000001000",
			3679 => "0000011100011000000100",
			3680 => "0000000011100110110001",
			3681 => "0000000011100110110001",
			3682 => "0000000011100110110001",
			3683 => "0011011111100100010000",
			3684 => "0011101100001100000100",
			3685 => "0000000011100110110001",
			3686 => "0010010010101100001000",
			3687 => "0000000100000000000100",
			3688 => "0000000011100110110001",
			3689 => "0000000011100110110001",
			3690 => "0000000011100110110001",
			3691 => "0000000011100110110001",
			3692 => "0011001011000000001000",
			3693 => "0011101000101000000100",
			3694 => "0000000011101000001101",
			3695 => "0000000011101000001101",
			3696 => "0001110100010000011000",
			3697 => "0010110010001000000100",
			3698 => "0000000011101000001101",
			3699 => "0001001110111000010000",
			3700 => "0001001011110000000100",
			3701 => "0000000011101000001101",
			3702 => "0011011010001000000100",
			3703 => "0000000011101000001101",
			3704 => "0011011100000000000100",
			3705 => "0000000011101000001101",
			3706 => "0000000011101000001101",
			3707 => "0000000011101000001101",
			3708 => "0001001011100000001100",
			3709 => "0011001111011100000100",
			3710 => "0000000011101000001101",
			3711 => "0010110010110100000100",
			3712 => "0000000011101000001101",
			3713 => "0000000011101000001101",
			3714 => "0000000011101000001101",
			3715 => "0010010111101100010100",
			3716 => "0011100001011100001100",
			3717 => "0001001100010000000100",
			3718 => "0000000011101010001001",
			3719 => "0011001111011100000100",
			3720 => "0000000011101010001001",
			3721 => "0000000011101010001001",
			3722 => "0001010010000100000100",
			3723 => "0000000011101010001001",
			3724 => "0000000011101010001001",
			3725 => "0011101011101100010000",
			3726 => "0001011100100100000100",
			3727 => "0000000011101010001001",
			3728 => "0000000111000100000100",
			3729 => "0000000011101010001001",
			3730 => "0000001010101100000100",
			3731 => "0000000011101010001001",
			3732 => "0000000011101010001001",
			3733 => "0000000111000000001000",
			3734 => "0010000001010100000100",
			3735 => "0000000011101010001001",
			3736 => "0000000011101010001001",
			3737 => "0001010110111100010000",
			3738 => "0001101000010000000100",
			3739 => "0000000011101010001001",
			3740 => "0001011001010000000100",
			3741 => "0000000011101010001001",
			3742 => "0001101001111100000100",
			3743 => "0000000011101010001001",
			3744 => "0000000011101010001001",
			3745 => "0000000011101010001001",
			3746 => "0011001000000000010100",
			3747 => "0010010000001000001000",
			3748 => "0011100010010100000100",
			3749 => "0000000011101011111101",
			3750 => "0000000011101011111101",
			3751 => "0001010111100000001000",
			3752 => "0001010010110100000100",
			3753 => "0000000011101011111101",
			3754 => "0000000011101011111101",
			3755 => "0000000011101011111101",
			3756 => "0001010110111100100100",
			3757 => "0000110011110000011000",
			3758 => "0011111000110100010000",
			3759 => "0001100101010000001100",
			3760 => "0000001111001000000100",
			3761 => "0000000011101011111101",
			3762 => "0010010010101100000100",
			3763 => "0000000011101011111101",
			3764 => "0000000011101011111101",
			3765 => "0000000011101011111101",
			3766 => "0000111110000000000100",
			3767 => "0000000011101011111101",
			3768 => "0000000011101011111101",
			3769 => "0010010010101100001000",
			3770 => "0000000111111000000100",
			3771 => "0000000011101011111101",
			3772 => "0000000011101011111101",
			3773 => "0000000011101011111101",
			3774 => "0000000011101011111101",
			3775 => "0011101011111000011000",
			3776 => "0000000001110100010100",
			3777 => "0001100100110100000100",
			3778 => "0000000011101101111001",
			3779 => "0010111011110100001100",
			3780 => "0011001101010100000100",
			3781 => "0000000011101101111001",
			3782 => "0010001000100100000100",
			3783 => "0000000011101101111001",
			3784 => "0000000011101101111001",
			3785 => "0000000011101101111001",
			3786 => "0000000011101101111001",
			3787 => "0011000001101000010000",
			3788 => "0001000110001100001100",
			3789 => "0001110110100100000100",
			3790 => "0000000011101101111001",
			3791 => "0001100101010000000100",
			3792 => "0000000011101101111001",
			3793 => "0000000011101101111001",
			3794 => "0000000011101101111001",
			3795 => "0011011111100100010100",
			3796 => "0011101100001100001000",
			3797 => "0001001101001000000100",
			3798 => "0000000011101101111001",
			3799 => "0000000011101101111001",
			3800 => "0010010010101100001000",
			3801 => "0000000100000000000100",
			3802 => "0000000011101101111001",
			3803 => "0000000011101101111001",
			3804 => "0000000011101101111001",
			3805 => "0000000011101101111001",
			3806 => "0010010111101100011000",
			3807 => "0011001000000000001000",
			3808 => "0011101000101000000100",
			3809 => "0000000011110000000101",
			3810 => "0000000011110000000101",
			3811 => "0001011110110100001000",
			3812 => "0011010011001000000100",
			3813 => "0000000011110000000101",
			3814 => "0000000011110000000101",
			3815 => "0011011111010100000100",
			3816 => "0000000011110000000101",
			3817 => "0000000011110000000101",
			3818 => "0011000100011000010000",
			3819 => "0010000001010100001100",
			3820 => "0010010000001000000100",
			3821 => "0000000011110000000101",
			3822 => "0011100110010000000100",
			3823 => "0000000011110000000101",
			3824 => "0000000011110000000101",
			3825 => "0000000011110000000101",
			3826 => "0001101000010000001000",
			3827 => "0000100110101100000100",
			3828 => "0000000011110000000101",
			3829 => "0000000011110000000101",
			3830 => "0010110001000000010100",
			3831 => "0010110101110100001000",
			3832 => "0011110011000000000100",
			3833 => "0000000011110000000101",
			3834 => "0000000011110000000101",
			3835 => "0000000111000000000100",
			3836 => "0000000011110000000101",
			3837 => "0010000111000100000100",
			3838 => "0000000011110000000101",
			3839 => "0000000011110000000101",
			3840 => "0000000011110000000101",
			3841 => "0001001000110100011100",
			3842 => "0011011100010100011000",
			3843 => "0001101000010000010100",
			3844 => "0000000010101000010000",
			3845 => "0001100100110100000100",
			3846 => "0000000011110001111001",
			3847 => "0000101000101000001000",
			3848 => "0001110011100000000100",
			3849 => "0000000011110001111001",
			3850 => "0000000011110001111001",
			3851 => "0000000011110001111001",
			3852 => "0000000011110001111001",
			3853 => "0000000011110001111001",
			3854 => "0000000011110001111001",
			3855 => "0011101000110100001000",
			3856 => "0000011110010100000100",
			3857 => "0000000011110001111001",
			3858 => "0000000011110001111001",
			3859 => "0011011111100100010100",
			3860 => "0001110111010000000100",
			3861 => "0000000011110001111001",
			3862 => "0000010001000100000100",
			3863 => "0000000011110001111001",
			3864 => "0000011100011000001000",
			3865 => "0011101000011100000100",
			3866 => "0000000011110001111001",
			3867 => "0000000011110001111001",
			3868 => "0000000011110001111001",
			3869 => "0000000011110001111001",
			3870 => "0011101110110100010000",
			3871 => "0001110110100100000100",
			3872 => "1111111011110011101101",
			3873 => "0001110110100100001000",
			3874 => "0011010001000000000100",
			3875 => "0000000011110011101101",
			3876 => "0000000011110011101101",
			3877 => "0000000011110011101101",
			3878 => "0011011111100100101000",
			3879 => "0011100110001100011000",
			3880 => "0000000010011000010100",
			3881 => "0010100011101000000100",
			3882 => "1111111011110011101101",
			3883 => "0000101000100000001000",
			3884 => "0000011101111100000100",
			3885 => "0000001011110011101101",
			3886 => "0000000011110011101101",
			3887 => "0000000111000000000100",
			3888 => "0000000011110011101101",
			3889 => "0000000011110011101101",
			3890 => "1111111011110011101101",
			3891 => "0010000111000100001100",
			3892 => "0001110101100100000100",
			3893 => "0000010011110011101101",
			3894 => "0000011100011000000100",
			3895 => "0000001011110011101101",
			3896 => "0000000011110011101101",
			3897 => "0000000011110011101101",
			3898 => "1111111011110011101101",
			3899 => "0000001101010000101100",
			3900 => "0001101011001100000100",
			3901 => "0000000011110101010001",
			3902 => "0000111101101100010100",
			3903 => "0001011100100100000100",
			3904 => "0000000011110101010001",
			3905 => "0001101001100100000100",
			3906 => "0000000011110101010001",
			3907 => "0000001010101100001000",
			3908 => "0000000110001000000100",
			3909 => "0000000011110101010001",
			3910 => "0000000011110101010001",
			3911 => "0000000011110101010001",
			3912 => "0011110110111000000100",
			3913 => "0000000011110101010001",
			3914 => "0001101000010000000100",
			3915 => "0000000011110101010001",
			3916 => "0000110010010100000100",
			3917 => "0000000011110101010001",
			3918 => "0010101000010100000100",
			3919 => "0000000011110101010001",
			3920 => "0000000011110101010001",
			3921 => "0000100011110100000100",
			3922 => "0000000011110101010001",
			3923 => "0000000011110101010001",
			3924 => "0010011010100000101000",
			3925 => "0011001011000000001000",
			3926 => "0001000110101100000100",
			3927 => "0000000011110111100101",
			3928 => "0000000011110111100101",
			3929 => "0000100010010100010000",
			3930 => "0001100100110100000100",
			3931 => "0000000011110111100101",
			3932 => "0001001000011100001000",
			3933 => "0010001000100100000100",
			3934 => "0000000011110111100101",
			3935 => "0000000011110111100101",
			3936 => "0000000011110111100101",
			3937 => "0011101011110000000100",
			3938 => "0000000011110111100101",
			3939 => "0000111110111000001000",
			3940 => "0011101000000100000100",
			3941 => "0000000011110111100101",
			3942 => "0000000011110111100101",
			3943 => "0000000011110111100101",
			3944 => "0011001011011100100000",
			3945 => "0010111011011100001000",
			3946 => "0001000011000000000100",
			3947 => "0000000011110111100101",
			3948 => "0000000011110111100101",
			3949 => "0000000111000100000100",
			3950 => "0000000011110111100101",
			3951 => "0000011010011000010000",
			3952 => "0011101111101000001000",
			3953 => "0011010110010000000100",
			3954 => "0000001011110111100101",
			3955 => "0000000011110111100101",
			3956 => "0011100110001100000100",
			3957 => "0000000011110111100101",
			3958 => "0000000011110111100101",
			3959 => "0000000011110111100101",
			3960 => "0000000011110111100101",
			3961 => "0010011010100000101100",
			3962 => "0001111111011100001000",
			3963 => "0001000110101100000100",
			3964 => "0000000011111010011001",
			3965 => "1111111011111010011001",
			3966 => "0010110010110100010100",
			3967 => "0001000011001100010000",
			3968 => "0011110000010000000100",
			3969 => "0000000011111010011001",
			3970 => "0010100011101000000100",
			3971 => "0000000011111010011001",
			3972 => "0001011100010100000100",
			3973 => "0000000011111010011001",
			3974 => "0000000011111010011001",
			3975 => "0000000011111010011001",
			3976 => "0000111000001000001100",
			3977 => "0011001111011100000100",
			3978 => "0000000011111010011001",
			3979 => "0011000001011000000100",
			3980 => "0000000011111010011001",
			3981 => "0000000011111010011001",
			3982 => "0000000011111010011001",
			3983 => "0011001001110100011100",
			3984 => "0000001000101100011000",
			3985 => "0001011100100100001000",
			3986 => "0011001010111000000100",
			3987 => "0000000011111010011001",
			3988 => "0000000011111010011001",
			3989 => "0011000100011000000100",
			3990 => "0000000011111010011001",
			3991 => "0000011101111100000100",
			3992 => "0000000011111010011001",
			3993 => "0010011010100000000100",
			3994 => "0000000011111010011001",
			3995 => "0000001011111010011001",
			3996 => "0000000011111010011001",
			3997 => "0000010100110100001100",
			3998 => "0011100011000000000100",
			3999 => "0000000011111010011001",
			4000 => "0001010111111100000100",
			4001 => "0000000011111010011001",
			4002 => "0000000011111010011001",
			4003 => "0010110101110100000100",
			4004 => "0000000011111010011001",
			4005 => "0000000011111010011001",
			4006 => "0001110110100100001100",
			4007 => "0000011101111100000100",
			4008 => "1111111011111100010101",
			4009 => "0011011110000100000100",
			4010 => "0000001011111100010101",
			4011 => "1111111011111100010101",
			4012 => "0011011111100100110000",
			4013 => "0000011010011000101000",
			4014 => "0001011111010000010000",
			4015 => "0011010110100000000100",
			4016 => "0000010011111100010101",
			4017 => "0000011101111100000100",
			4018 => "1111111011111100010101",
			4019 => "0011101011101100000100",
			4020 => "0000001011111100010101",
			4021 => "1111111011111100010101",
			4022 => "0001000011101100001100",
			4023 => "0000011001011000000100",
			4024 => "0000011011111100010101",
			4025 => "0001100100111100000100",
			4026 => "1111111011111100010101",
			4027 => "0000001011111100010101",
			4028 => "0011101001001100000100",
			4029 => "1111111011111100010101",
			4030 => "0001111010010100000100",
			4031 => "0000000011111100010101",
			4032 => "0000010011111100010101",
			4033 => "0011001000000000000100",
			4034 => "0000001011111100010101",
			4035 => "1111111011111100010101",
			4036 => "1111111011111100010101",
			4037 => "0001110110100100001100",
			4038 => "0000011101111100000100",
			4039 => "1111111011111110011001",
			4040 => "0011011110000100000100",
			4041 => "0000001011111110011001",
			4042 => "1111111011111110011001",
			4043 => "0011011111100100110100",
			4044 => "0011100110001100100000",
			4045 => "0000001111000100011000",
			4046 => "0000011010011000010000",
			4047 => "0001101000010000001000",
			4048 => "0000011101011100000100",
			4049 => "0000001011111110011001",
			4050 => "0000000011111110011001",
			4051 => "0011011001011100000100",
			4052 => "1111111011111110011001",
			4053 => "0000001011111110011001",
			4054 => "0011011110010000000100",
			4055 => "0000001011111110011001",
			4056 => "1111111011111110011001",
			4057 => "0011101100001100000100",
			4058 => "1111111011111110011001",
			4059 => "0000000011111110011001",
			4060 => "0001110000011100000100",
			4061 => "0000100011111110011001",
			4062 => "0010000111000100001100",
			4063 => "0000011100011000001000",
			4064 => "0001000011101100000100",
			4065 => "0000001011111110011001",
			4066 => "0000001011111110011001",
			4067 => "0000000011111110011001",
			4068 => "0000000011111110011001",
			4069 => "1111111011111110011001",
			4070 => "0000000010101000100100",
			4071 => "0010011010100100011000",
			4072 => "0001101001100100010100",
			4073 => "0011010101110000010000",
			4074 => "0001100100110100000100",
			4075 => "0000000100000000111101",
			4076 => "0001110001101000001000",
			4077 => "0001111000000000000100",
			4078 => "0000000100000000111101",
			4079 => "0000000100000000111101",
			4080 => "0000000100000000111101",
			4081 => "0000000100000000111101",
			4082 => "0000000100000000111101",
			4083 => "0001111111011100001000",
			4084 => "0000110001011100000100",
			4085 => "0000001100000000111101",
			4086 => "0000000100000000111101",
			4087 => "0000000100000000111101",
			4088 => "0011100001011100000100",
			4089 => "1111111100000000111101",
			4090 => "0011101100001100011000",
			4091 => "0001001010110100010100",
			4092 => "0010011010100100001100",
			4093 => "0001110100010000001000",
			4094 => "0001010101110000000100",
			4095 => "0000000100000000111101",
			4096 => "0000000100000000111101",
			4097 => "0000000100000000111101",
			4098 => "0011100011000000000100",
			4099 => "0000000100000000111101",
			4100 => "0000000100000000111101",
			4101 => "0000000100000000111101",
			4102 => "0010110001000000010000",
			4103 => "0010110000110100000100",
			4104 => "0000000100000000111101",
			4105 => "0010010010101100001000",
			4106 => "0000001100001000000100",
			4107 => "0000001100000000111101",
			4108 => "0000000100000000111101",
			4109 => "0000000100000000111101",
			4110 => "0000000100000000111101",
			4111 => "0011001010111000001000",
			4112 => "0010010010101100000100",
			4113 => "1111111100000010111001",
			4114 => "0000000100000010111001",
			4115 => "0011011111100100110100",
			4116 => "0011100101000000100100",
			4117 => "0001001010110100011100",
			4118 => "0011101111101000010000",
			4119 => "0010011010100100001000",
			4120 => "0001101111000000000100",
			4121 => "0000000100000010111001",
			4122 => "0000000100000010111001",
			4123 => "0011001000000000000100",
			4124 => "0000001100000010111001",
			4125 => "0000000100000010111001",
			4126 => "0010010010101100001000",
			4127 => "0001110111010000000100",
			4128 => "0000000100000010111001",
			4129 => "0000001100000010111001",
			4130 => "1111111100000010111001",
			4131 => "0011101000110100000100",
			4132 => "1111111100000010111001",
			4133 => "0000000100000010111001",
			4134 => "0000011100011000001100",
			4135 => "0000001011000100001000",
			4136 => "0000110101000000000100",
			4137 => "0000000100000010111001",
			4138 => "0000001100000010111001",
			4139 => "0000000100000010111001",
			4140 => "0000000100000010111001",
			4141 => "1111111100000010111001",
			4142 => "0001000010010100101000",
			4143 => "0011101011111000100100",
			4144 => "0001101011001100010000",
			4145 => "0001001100010000001100",
			4146 => "0001000010000100000100",
			4147 => "0000000100000101111101",
			4148 => "0010011011001100000100",
			4149 => "0000000100000101111101",
			4150 => "0000000100000101111101",
			4151 => "0000000100000101111101",
			4152 => "0010101000100100010000",
			4153 => "0010100011101000000100",
			4154 => "0000000100000101111101",
			4155 => "0011100110010000000100",
			4156 => "0000000100000101111101",
			4157 => "0001011110101100000100",
			4158 => "0000000100000101111101",
			4159 => "0000001100000101111101",
			4160 => "0000000100000101111101",
			4161 => "0000000100000101111101",
			4162 => "0011101000101000010000",
			4163 => "0010010010101100001000",
			4164 => "0000011010011000000100",
			4165 => "1111111100000101111101",
			4166 => "0000000100000101111101",
			4167 => "0000011010011000000100",
			4168 => "0000000100000101111101",
			4169 => "0000000100000101111101",
			4170 => "0011100011000000010000",
			4171 => "0001101000010000001100",
			4172 => "0000100010010100000100",
			4173 => "0000000100000101111101",
			4174 => "0001100100111100000100",
			4175 => "0000000100000101111101",
			4176 => "0000000100000101111101",
			4177 => "0000000100000101111101",
			4178 => "0000011100011000011000",
			4179 => "0011000100000100001100",
			4180 => "0001101000010000000100",
			4181 => "0000000100000101111101",
			4182 => "0011001001110100000100",
			4183 => "0000000100000101111101",
			4184 => "0000000100000101111101",
			4185 => "0001101001111100001000",
			4186 => "0010011001111100000100",
			4187 => "0000000100000101111101",
			4188 => "0000000100000101111101",
			4189 => "0000000100000101111101",
			4190 => "1111111100000101111101",
			4191 => "0010110001000001000000",
			4192 => "0011101100001100110000",
			4193 => "0000001101010000101000",
			4194 => "0011111111101000010000",
			4195 => "0011011100010100001100",
			4196 => "0010011010100000000100",
			4197 => "0000000100001000000001",
			4198 => "0010011010100100000100",
			4199 => "0000000100001000000001",
			4200 => "0000000100001000000001",
			4201 => "0000000100001000000001",
			4202 => "0010111011110100001000",
			4203 => "0001111111011100000100",
			4204 => "0000000100001000000001",
			4205 => "0000000100001000000001",
			4206 => "0000000111000000001000",
			4207 => "0000110010010100000100",
			4208 => "0000000100001000000001",
			4209 => "0000000100001000000001",
			4210 => "0011100011000000000100",
			4211 => "0000000100001000000001",
			4212 => "0000000100001000000001",
			4213 => "0000001111000100000100",
			4214 => "0000000100001000000001",
			4215 => "0000000100001000000001",
			4216 => "0011000110100100000100",
			4217 => "0000000100001000000001",
			4218 => "0010010010101100001000",
			4219 => "0000000100000000000100",
			4220 => "0000001100001000000001",
			4221 => "0000000100001000000001",
			4222 => "0000000100001000000001",
			4223 => "0000000100001000000001",
			4224 => "0001000010010100101000",
			4225 => "0011101011111000100100",
			4226 => "0010000101000100100000",
			4227 => "0010100011101000010100",
			4228 => "0010110111010000001100",
			4229 => "0010111010011100000100",
			4230 => "0000000100001011001101",
			4231 => "0001001000001100000100",
			4232 => "0000000100001011001101",
			4233 => "0000000100001011001101",
			4234 => "0010110100000100000100",
			4235 => "0000000100001011001101",
			4236 => "0000000100001011001101",
			4237 => "0011011100100100000100",
			4238 => "0000000100001011001101",
			4239 => "0011101110110100000100",
			4240 => "0000000100001011001101",
			4241 => "0000001100001011001101",
			4242 => "0000000100001011001101",
			4243 => "0000000100001011001101",
			4244 => "0011101000101000010100",
			4245 => "0010010010101100001100",
			4246 => "0001001011110000000100",
			4247 => "0000000100001011001101",
			4248 => "0000011010011000000100",
			4249 => "1111111100001011001101",
			4250 => "0000000100001011001101",
			4251 => "0000011010011000000100",
			4252 => "0000000100001011001101",
			4253 => "0000000100001011001101",
			4254 => "0000011100011000100000",
			4255 => "0010110010110100010000",
			4256 => "0011010011001000000100",
			4257 => "0000000100001011001101",
			4258 => "0001001110111000001000",
			4259 => "0001001000011100000100",
			4260 => "0000000100001011001101",
			4261 => "0000001100001011001101",
			4262 => "0000000100001011001101",
			4263 => "0011101110100100000100",
			4264 => "0000000100001011001101",
			4265 => "0011010000010000001000",
			4266 => "0010110111100000000100",
			4267 => "0000000100001011001101",
			4268 => "0000000100001011001101",
			4269 => "0000000100001011001101",
			4270 => "0011100011000000001000",
			4271 => "0011001001110100000100",
			4272 => "0000000100001011001101",
			4273 => "0000000100001011001101",
			4274 => "1111111100001011001101",
			4275 => "0000101110100101000100",
			4276 => "0000101110000000101100",
			4277 => "0011100110010000001100",
			4278 => "0011001011000000000100",
			4279 => "1100000100001110101001",
			4280 => "0011001011000000000100",
			4281 => "1100001100001110101001",
			4282 => "1100000100001110101001",
			4283 => "0011011001100000011100",
			4284 => "0000011100011000010000",
			4285 => "0001110111010000001000",
			4286 => "0010011010100000000100",
			4287 => "1100000100001110101001",
			4288 => "1100001100001110101001",
			4289 => "0000000001110100000100",
			4290 => "1100010100001110101001",
			4291 => "1110011100001110101001",
			4292 => "0000101100111000000100",
			4293 => "1111100100001110101001",
			4294 => "0000011100011000000100",
			4295 => "1100101100001110101001",
			4296 => "1100001100001110101001",
			4297 => "1100000100001110101001",
			4298 => "0010010111101100001000",
			4299 => "0000000010011000000100",
			4300 => "0000101100001110101001",
			4301 => "1100000100001110101001",
			4302 => "0010011010100100001100",
			4303 => "0001010101110000000100",
			4304 => "1100000100001110101001",
			4305 => "0001110000011100000100",
			4306 => "1110111100001110101001",
			4307 => "1100011100001110101001",
			4308 => "1100000100001110101001",
			4309 => "0010001111001000100100",
			4310 => "0010010000001000001000",
			4311 => "0000111000000100000100",
			4312 => "1100000100001110101001",
			4313 => "0001000100001110101001",
			4314 => "0011100010111000010100",
			4315 => "0010011010100100001000",
			4316 => "0001010111111100000100",
			4317 => "1100000100001110101001",
			4318 => "1110110100001110101001",
			4319 => "0010010010101100001000",
			4320 => "0000100110001100000100",
			4321 => "1100000100001110101001",
			4322 => "1100011100001110101001",
			4323 => "1100000100001110101001",
			4324 => "0000011010011000000100",
			4325 => "1111011100001110101001",
			4326 => "1100000100001110101001",
			4327 => "0010000111000100000100",
			4328 => "1100011100001110101001",
			4329 => "1100000100001110101001",
			4330 => "0010010111101100101100",
			4331 => "0011001000000000001000",
			4332 => "0011111000000100000100",
			4333 => "1111111100010010001101",
			4334 => "0000000100010010001101",
			4335 => "0011011010000100011100",
			4336 => "0000010101011100001100",
			4337 => "0000011101011100001000",
			4338 => "0011111011110000000100",
			4339 => "0000000100010010001101",
			4340 => "0000000100010010001101",
			4341 => "0000000100010010001101",
			4342 => "0000000010101000000100",
			4343 => "0000000100010010001101",
			4344 => "0001000011010100001000",
			4345 => "0010101010110000000100",
			4346 => "0000001100010010001101",
			4347 => "0000000100010010001101",
			4348 => "0000000100010010001101",
			4349 => "0011100101000000000100",
			4350 => "0000000100010010001101",
			4351 => "0000000100010010001101",
			4352 => "0001001011110000011100",
			4353 => "0010110010001000010100",
			4354 => "0010010000001000000100",
			4355 => "0000000100010010001101",
			4356 => "0000000010101000001100",
			4357 => "0011011100100100000100",
			4358 => "0000000100010010001101",
			4359 => "0010100011101000000100",
			4360 => "0000000100010010001101",
			4361 => "0000001100010010001101",
			4362 => "0000000100010010001101",
			4363 => "0000111011101100000100",
			4364 => "0000000100010010001101",
			4365 => "0000000100010010001101",
			4366 => "0001111111011100001100",
			4367 => "0000011010011000000100",
			4368 => "1111111100010010001101",
			4369 => "0000001000110000000100",
			4370 => "0000000100010010001101",
			4371 => "0000000100010010001101",
			4372 => "0001110101100100010000",
			4373 => "0010001001101000001100",
			4374 => "0000000111000000000100",
			4375 => "0000000100010010001101",
			4376 => "0010010010101100000100",
			4377 => "0000001100010010001101",
			4378 => "0000000100010010001101",
			4379 => "0000000100010010001101",
			4380 => "0000010100110100001100",
			4381 => "0010100110011000000100",
			4382 => "0000000100010010001101",
			4383 => "0011000001011000000100",
			4384 => "0000000100010010001101",
			4385 => "0000000100010010001101",
			4386 => "0000000100010010001101",
			4387 => "0011001101010100000100",
			4388 => "1111111100010100110001",
			4389 => "0001110101100100111000",
			4390 => "0010011010100100100100",
			4391 => "0001101001100100010100",
			4392 => "0010010000001000001000",
			4393 => "0000011001011000000100",
			4394 => "0000000100010100110001",
			4395 => "0000000100010100110001",
			4396 => "0011000100011000001000",
			4397 => "0011011100100100000100",
			4398 => "0000000100010100110001",
			4399 => "0000001100010100110001",
			4400 => "0000000100010100110001",
			4401 => "0001110111010000000100",
			4402 => "1111111100010100110001",
			4403 => "0001001010110100001000",
			4404 => "0011001000011000000100",
			4405 => "0000001100010100110001",
			4406 => "0000000100010100110001",
			4407 => "0000000100010100110001",
			4408 => "0001101000010000001000",
			4409 => "0001111111011100000100",
			4410 => "0000001100010100110001",
			4411 => "0000000100010100110001",
			4412 => "0010110101110100000100",
			4413 => "0000000100010100110001",
			4414 => "0010010010101100000100",
			4415 => "0000000100010100110001",
			4416 => "0000000100010100110001",
			4417 => "0011101000000100001000",
			4418 => "0000010101011100000100",
			4419 => "0000000100010100110001",
			4420 => "1111111100010100110001",
			4421 => "0001111010010100001100",
			4422 => "0000010100110100001000",
			4423 => "0000000100000000000100",
			4424 => "0000000100010100110001",
			4425 => "0000000100010100110001",
			4426 => "0000000100010100110001",
			4427 => "0000000100010100110001",
			4428 => "0010000001010100101100",
			4429 => "0011011100010100101000",
			4430 => "0001100100110100000100",
			4431 => "0000000100010111101101",
			4432 => "0010111011011100011000",
			4433 => "0000110110111100001100",
			4434 => "0010001100011100001000",
			4435 => "0010110100000100000100",
			4436 => "0000000100010111101101",
			4437 => "0000000100010111101101",
			4438 => "0000000100010111101101",
			4439 => "0011001101010100000100",
			4440 => "0000000100010111101101",
			4441 => "0001010111100000000100",
			4442 => "0000000100010111101101",
			4443 => "0000000100010111101101",
			4444 => "0010001100011100000100",
			4445 => "0000000100010111101101",
			4446 => "0001110001101000000100",
			4447 => "0000000100010111101101",
			4448 => "0000001100010111101101",
			4449 => "0000000100010111101101",
			4450 => "0011011100010100001000",
			4451 => "0010111011110100000100",
			4452 => "1111111100010111101101",
			4453 => "0000000100010111101101",
			4454 => "0001110100010000010000",
			4455 => "0001001110111000001100",
			4456 => "0001101000010000000100",
			4457 => "0000000100010111101101",
			4458 => "0010010010101100000100",
			4459 => "0000001100010111101101",
			4460 => "0000000100010111101101",
			4461 => "0000000100010111101101",
			4462 => "0001101001111100010000",
			4463 => "0001110100010000000100",
			4464 => "0000000100010111101101",
			4465 => "0010110010110100000100",
			4466 => "0000000100010111101101",
			4467 => "0011001111011100000100",
			4468 => "0000000100010111101101",
			4469 => "0000000100010111101101",
			4470 => "0000010100110100001000",
			4471 => "0001000111011100000100",
			4472 => "0000000100010111101101",
			4473 => "0000000100010111101101",
			4474 => "0000000100010111101101",
			4475 => "0000010101011100011000",
			4476 => "0000000111000000010100",
			4477 => "0011101010000100001100",
			4478 => "0011001011000000000100",
			4479 => "1111111100011010110001",
			4480 => "0001010110100000000100",
			4481 => "0000100100011010110001",
			4482 => "1111111100011010110001",
			4483 => "0010111011110100000100",
			4484 => "0000110100011010110001",
			4485 => "0000000100011010110001",
			4486 => "1111111100011010110001",
			4487 => "0010010010101101000100",
			4488 => "0001011001010000100000",
			4489 => "0001000110111000011000",
			4490 => "0010011010100000001100",
			4491 => "0010010000001000000100",
			4492 => "1111111100011010110001",
			4493 => "0001001111100100000100",
			4494 => "0000110100011010110001",
			4495 => "0000000100011010110001",
			4496 => "0011101000001100000100",
			4497 => "0000100100011010110001",
			4498 => "0010101000100100000100",
			4499 => "1111111100011010110001",
			4500 => "0000001100011010110001",
			4501 => "0000011100011000000100",
			4502 => "1111111100011010110001",
			4503 => "0000000100011010110001",
			4504 => "0010000001010100010000",
			4505 => "0010010101010000001000",
			4506 => "0010111011110100000100",
			4507 => "0000000100011010110001",
			4508 => "0000001100011010110001",
			4509 => "0001110101110100000100",
			4510 => "1111111100011010110001",
			4511 => "1111110100011010110001",
			4512 => "0001010111011000010000",
			4513 => "0011001000000000001000",
			4514 => "0011101111101000000100",
			4515 => "0000111100011010110001",
			4516 => "0000001100011010110001",
			4517 => "0001100100111100000100",
			4518 => "0000000100011010110001",
			4519 => "0000001100011010110001",
			4520 => "1111111100011010110001",
			4521 => "0001001011110000000100",
			4522 => "0000001100011010110001",
			4523 => "1111111100011010110001",
			4524 => "0000010101011100010100",
			4525 => "0000000111000000010000",
			4526 => "0000111000100000001100",
			4527 => "0011001011000000000100",
			4528 => "1111111100011101101101",
			4529 => "0010110000011100000100",
			4530 => "0001000100011101101101",
			4531 => "1111111100011101101101",
			4532 => "0000100100011101101101",
			4533 => "1111111100011101101101",
			4534 => "0010010010101101000100",
			4535 => "0001010101110000101000",
			4536 => "0010011010100000011000",
			4537 => "0000100110111100001000",
			4538 => "0010100011101000000100",
			4539 => "1111111100011101101101",
			4540 => "0000111100011101101101",
			4541 => "0011010111111100001000",
			4542 => "0001010111100000000100",
			4543 => "1111111100011101101101",
			4544 => "0000000100011101101101",
			4545 => "0001010101001000000100",
			4546 => "1111111100011101101101",
			4547 => "1111111100011101101101",
			4548 => "0000101111100100000100",
			4549 => "0000100100011101101101",
			4550 => "0000011100011000000100",
			4551 => "1111111100011101101101",
			4552 => "0010101001000100000100",
			4553 => "0000010100011101101101",
			4554 => "1111111100011101101101",
			4555 => "0010101000010100001100",
			4556 => "0001110000011100000100",
			4557 => "0000001100011101101101",
			4558 => "0001110101110100000100",
			4559 => "1111111100011101101101",
			4560 => "1111110100011101101101",
			4561 => "0001010111011000001100",
			4562 => "0000101011110000000100",
			4563 => "0000011100011101101101",
			4564 => "0010101001000100000100",
			4565 => "1111110100011101101101",
			4566 => "0000001100011101101101",
			4567 => "1111111100011101101101",
			4568 => "0000110011000000000100",
			4569 => "0000010100011101101101",
			4570 => "1111111100011101101101",
			4571 => "0000000010101000111000",
			4572 => "0010010000001000010000",
			4573 => "0001101001100100000100",
			4574 => "0000000100100001000001",
			4575 => "0010100111110100001000",
			4576 => "0000000110001000000100",
			4577 => "0000000100100001000001",
			4578 => "0000000100100001000001",
			4579 => "0000000100100001000001",
			4580 => "0000111101101100100000",
			4581 => "0010111011011100011000",
			4582 => "0010100111110100001100",
			4583 => "0001110110100100001000",
			4584 => "0011101110110100000100",
			4585 => "0000000100100001000001",
			4586 => "0000000100100001000001",
			4587 => "0000000100100001000001",
			4588 => "0011111000001100000100",
			4589 => "0000000100100001000001",
			4590 => "0010110000011100000100",
			4591 => "0000000100100001000001",
			4592 => "0000000100100001000001",
			4593 => "0000000111000100000100",
			4594 => "0000000100100001000001",
			4595 => "0000001100100001000001",
			4596 => "0000000010101000000100",
			4597 => "0000000100100001000001",
			4598 => "0000000100100001000001",
			4599 => "0011100001011100000100",
			4600 => "1111111100100001000001",
			4601 => "0001110111110000101000",
			4602 => "0011011100010100010100",
			4603 => "0001101000010000001100",
			4604 => "0011001011000000000100",
			4605 => "0000000100100001000001",
			4606 => "0011010111111100000100",
			4607 => "0000000100100001000001",
			4608 => "0000000100100001000001",
			4609 => "0001111000011000000100",
			4610 => "0000000100100001000001",
			4611 => "0000000100100001000001",
			4612 => "0001101000010000000100",
			4613 => "0000000100100001000001",
			4614 => "0000000010011000001000",
			4615 => "0010010010101100000100",
			4616 => "0000001100100001000001",
			4617 => "0000000100100001000001",
			4618 => "0011100110001100000100",
			4619 => "0000000100100001000001",
			4620 => "0000000100100001000001",
			4621 => "0011011000001100000100",
			4622 => "0000000100100001000001",
			4623 => "0000000100100001000001",
			4624 => "0010111010011100000100",
			4625 => "1111111100100010110101",
			4626 => "0001011111010100110100",
			4627 => "0011101100001100100100",
			4628 => "0001001001001100100000",
			4629 => "0001110101100100010000",
			4630 => "0001111111011100001000",
			4631 => "0011001000000000000100",
			4632 => "0000000100100010110101",
			4633 => "1111111100100010110101",
			4634 => "0010100001010000000100",
			4635 => "0000001100100010110101",
			4636 => "0000000100100010110101",
			4637 => "0010001100000100001000",
			4638 => "0010101001000100000100",
			4639 => "1111111100100010110101",
			4640 => "0000000100100010110101",
			4641 => "0000011100011000000100",
			4642 => "0000001100100010110101",
			4643 => "0000000100100010110101",
			4644 => "1111111100100010110101",
			4645 => "0000011100011000001100",
			4646 => "0000001011000100001000",
			4647 => "0000110110001100000100",
			4648 => "0000000100100010110101",
			4649 => "0000001100100010110101",
			4650 => "0000000100100010110101",
			4651 => "0000000100100010110101",
			4652 => "1111111100100010110101",
			4653 => "0010010111101100110100",
			4654 => "0011001000000000001000",
			4655 => "0011111000000100000100",
			4656 => "1111111100100110110001",
			4657 => "0000000100100110110001",
			4658 => "0001011110110100100100",
			4659 => "0000010101011100010100",
			4660 => "0011001001110100001100",
			4661 => "0001010010011100001000",
			4662 => "0010001000010100000100",
			4663 => "0000000100100110110001",
			4664 => "0000000100100110110001",
			4665 => "0000000100100110110001",
			4666 => "0001010011001000000100",
			4667 => "0000000100100110110001",
			4668 => "0000000100100110110001",
			4669 => "0000000010101000000100",
			4670 => "0000000100100110110001",
			4671 => "0001000011010100001000",
			4672 => "0010001011010100000100",
			4673 => "0000001100100110110001",
			4674 => "0000000100100110110001",
			4675 => "0000000100100110110001",
			4676 => "0000011110010100000100",
			4677 => "0000000100100110110001",
			4678 => "0000000100100110110001",
			4679 => "0001001011110000100000",
			4680 => "0010110010001000011000",
			4681 => "0010010000001000000100",
			4682 => "0000000100100110110001",
			4683 => "0000000010101000010000",
			4684 => "0001011100100100001000",
			4685 => "0000111111010100000100",
			4686 => "0000000100100110110001",
			4687 => "0000000100100110110001",
			4688 => "0010100111110100000100",
			4689 => "0000000100100110110001",
			4690 => "0000001100100110110001",
			4691 => "0000000100100110110001",
			4692 => "0000111011101100000100",
			4693 => "0000000100100110110001",
			4694 => "0000000100100110110001",
			4695 => "0001111111011100001100",
			4696 => "0000011010011000000100",
			4697 => "1111111100100110110001",
			4698 => "0000001000110000000100",
			4699 => "0000000100100110110001",
			4700 => "0000000100100110110001",
			4701 => "0001110101100100010000",
			4702 => "0010001001101000001100",
			4703 => "0000000111000000000100",
			4704 => "0000000100100110110001",
			4705 => "0010010010101100000100",
			4706 => "0000001100100110110001",
			4707 => "0000000100100110110001",
			4708 => "0000000100100110110001",
			4709 => "0000010100110100001100",
			4710 => "0001100101010000000100",
			4711 => "0000000100100110110001",
			4712 => "0011000001011000000100",
			4713 => "0000000100100110110001",
			4714 => "0000000100100110110001",
			4715 => "0000000100100110110001",
			4716 => "0011001101010100000100",
			4717 => "1111111100101001101101",
			4718 => "0001000011001100111100",
			4719 => "0010101000010100100000",
			4720 => "0000111100111000010100",
			4721 => "0010011010100100010000",
			4722 => "0000011001011000001000",
			4723 => "0001100100110100000100",
			4724 => "0000000100101001101101",
			4725 => "0000000100101001101101",
			4726 => "0010110100000100000100",
			4727 => "0000000100101001101101",
			4728 => "0000000100101001101101",
			4729 => "0000000100101001101101",
			4730 => "0011001000000000000100",
			4731 => "0000000100101001101101",
			4732 => "0010000001010100000100",
			4733 => "0000000100101001101101",
			4734 => "0000000100101001101101",
			4735 => "0011010010000100010100",
			4736 => "0001111000011000001000",
			4737 => "0010101000010100000100",
			4738 => "0000000100101001101101",
			4739 => "0000000100101001101101",
			4740 => "0010100001010000001000",
			4741 => "0011011001011100000100",
			4742 => "0000000100101001101101",
			4743 => "0000001100101001101101",
			4744 => "0000000100101001101101",
			4745 => "0010001100000100000100",
			4746 => "0000000100101001101101",
			4747 => "0000000100101001101101",
			4748 => "0011101000110100001000",
			4749 => "0001000011001100000100",
			4750 => "0000000100101001101101",
			4751 => "1111111100101001101101",
			4752 => "0001011100010000010000",
			4753 => "0010011010100100001100",
			4754 => "0001011110010000000100",
			4755 => "0000000100101001101101",
			4756 => "0000011011111100000100",
			4757 => "0000000100101001101101",
			4758 => "0000001100101001101101",
			4759 => "0000000100101001101101",
			4760 => "0001101001111100000100",
			4761 => "0000000100101001101101",
			4762 => "0000000100101001101101",
			4763 => "0000010101011100000100",
			4764 => "1111111100101100001001",
			4765 => "0000011100011001000100",
			4766 => "0001011001010000100000",
			4767 => "0010011010100000001100",
			4768 => "0000100110111100001000",
			4769 => "0010010000001000000100",
			4770 => "1111111100101100001001",
			4771 => "0000010100101100001001",
			4772 => "1111111100101100001001",
			4773 => "0001000011000000000100",
			4774 => "0000010100101100001001",
			4775 => "0011011001011100001000",
			4776 => "0000011100011000000100",
			4777 => "1111111100101100001001",
			4778 => "0000000100101100001001",
			4779 => "0010110010001000000100",
			4780 => "0000110100101100001001",
			4781 => "0000000100101100001001",
			4782 => "0001101000010000001100",
			4783 => "0011011100010100001000",
			4784 => "0001101011001100000100",
			4785 => "0000000100101100001001",
			4786 => "0000010100101100001001",
			4787 => "1111111100101100001001",
			4788 => "0001000101010100001100",
			4789 => "0000011101111100000100",
			4790 => "0000001100101100001001",
			4791 => "0001000101000000000100",
			4792 => "0000000100101100001001",
			4793 => "0000010100101100001001",
			4794 => "0011101110100100000100",
			4795 => "1111111100101100001001",
			4796 => "0011001011011100000100",
			4797 => "0000001100101100001001",
			4798 => "0000000100101100001001",
			4799 => "0000110001011100000100",
			4800 => "0000001100101100001001",
			4801 => "1111111100101100001001",
			4802 => "0010011000010000000100",
			4803 => "1111111100101110110101",
			4804 => "0010010010101101001100",
			4805 => "0001011001010000101000",
			4806 => "0010011010100100010100",
			4807 => "0000100110111100001000",
			4808 => "0010010000001000000100",
			4809 => "1111111100101110110101",
			4810 => "0000010100101110110101",
			4811 => "0011001000000000000100",
			4812 => "1111111100101110110101",
			4813 => "0001110001101000000100",
			4814 => "0000011100101110110101",
			4815 => "1111111100101110110101",
			4816 => "0001011110000100001100",
			4817 => "0011010111111100001000",
			4818 => "0001000110111000000100",
			4819 => "0000010100101110110101",
			4820 => "1111111100101110110101",
			4821 => "0000100100101110110101",
			4822 => "0010110100010000000100",
			4823 => "1111111100101110110101",
			4824 => "0000000100101110110101",
			4825 => "0001101000010000001100",
			4826 => "0011011100010100001000",
			4827 => "0000111011101100000100",
			4828 => "0000000100101110110101",
			4829 => "0000001100101110110101",
			4830 => "1111111100101110110101",
			4831 => "0000001101010000001100",
			4832 => "0010010010101100001000",
			4833 => "0010011010100000000100",
			4834 => "0000001100101110110101",
			4835 => "0000001100101110110101",
			4836 => "1111111100101110110101",
			4837 => "0011101000011100000100",
			4838 => "1111111100101110110101",
			4839 => "0010100001010000000100",
			4840 => "0000000100101110110101",
			4841 => "0000001100101110110101",
			4842 => "0011001010111000000100",
			4843 => "0000000100101110110101",
			4844 => "1111111100101110110101",
			4845 => "0000010101011100000100",
			4846 => "1111111100110001011001",
			4847 => "0000011100011001001000",
			4848 => "0001011001010000101000",
			4849 => "0010011010100000001100",
			4850 => "0000101100000000001000",
			4851 => "0011110111011000000100",
			4852 => "1111111100110001011001",
			4853 => "0000001100110001011001",
			4854 => "1111111100110001011001",
			4855 => "0001000011000000001100",
			4856 => "0001101111000000000100",
			4857 => "0000010100110001011001",
			4858 => "0001110001101000000100",
			4859 => "1111111100110001011001",
			4860 => "0000001100110001011001",
			4861 => "0011011001011100001000",
			4862 => "0000011100011000000100",
			4863 => "1111111100110001011001",
			4864 => "0000000100110001011001",
			4865 => "0001011110000100000100",
			4866 => "0000101100110001011001",
			4867 => "0000000100110001011001",
			4868 => "0001100100111100000100",
			4869 => "1111111100110001011001",
			4870 => "0001001010110100010000",
			4871 => "0000000010101000001000",
			4872 => "0001001110000000000100",
			4873 => "0000010100110001011001",
			4874 => "1111111100110001011001",
			4875 => "0001111011011100000100",
			4876 => "0000001100110001011001",
			4877 => "0000001100110001011001",
			4878 => "0000111100001100000100",
			4879 => "1111111100110001011001",
			4880 => "0011010111010100000100",
			4881 => "0000001100110001011001",
			4882 => "0000000100110001011001",
			4883 => "0000110001011100000100",
			4884 => "0000001100110001011001",
			4885 => "1111111100110001011001",
			4886 => "0001110011100000000100",
			4887 => "1111111100110100001101",
			4888 => "0011101011111000011100",
			4889 => "0010100011101000001000",
			4890 => "0000011111001100000100",
			4891 => "0000001100110100001101",
			4892 => "1111111100110100001101",
			4893 => "0000000001110100010000",
			4894 => "0011100110010000000100",
			4895 => "0000000100110100001101",
			4896 => "0001000010010100001000",
			4897 => "0000001011010100000100",
			4898 => "0000000100110100001101",
			4899 => "0000001100110100001101",
			4900 => "0000000100110100001101",
			4901 => "0000000100110100001101",
			4902 => "0000000010101000000100",
			4903 => "1111111100110100001101",
			4904 => "0011001000011000011100",
			4905 => "0000011100011000001100",
			4906 => "0001011001010000000100",
			4907 => "1111111100110100001101",
			4908 => "0011100010010100000100",
			4909 => "0000000100110100001101",
			4910 => "0000001100110100001101",
			4911 => "0010110010001000001000",
			4912 => "0010110110110100000100",
			4913 => "0000000100110100001101",
			4914 => "0000000100110100001101",
			4915 => "0010010010101100000100",
			4916 => "0000001100110100001101",
			4917 => "0000000100110100001101",
			4918 => "0011101000011100001100",
			4919 => "0001001101001000001000",
			4920 => "0010000001110000000100",
			4921 => "0000000100110100001101",
			4922 => "0000000100110100001101",
			4923 => "1111111100110100001101",
			4924 => "0010110001000000001000",
			4925 => "0000010100110100000100",
			4926 => "0000001100110100001101",
			4927 => "0000000100110100001101",
			4928 => "0011011111100100000100",
			4929 => "0000000100110100001101",
			4930 => "1111111100110100001101",
			4931 => "0001111000000000000100",
			4932 => "1111111100111000000011",
			4933 => "0000011101111100101100",
			4934 => "0001110111010000010100",
			4935 => "0011111010001000001100",
			4936 => "0011111001011100000100",
			4937 => "0000000100111000000011",
			4938 => "0010000011101000000100",
			4939 => "0000000100111000000011",
			4940 => "0000000100111000000011",
			4941 => "0001110111010000000100",
			4942 => "1111111100111000000011",
			4943 => "0000000100111000000011",
			4944 => "0011011111010100010000",
			4945 => "0000010001111000001100",
			4946 => "0001100100111100000100",
			4947 => "0000000100111000000011",
			4948 => "0000000011010000000100",
			4949 => "0000001100111000000011",
			4950 => "0000000100111000000011",
			4951 => "0000000100111000000011",
			4952 => "0000011110010100000100",
			4953 => "1111111100111000000011",
			4954 => "0000000100111000000011",
			4955 => "0000010100110100100000",
			4956 => "0011011001011100010000",
			4957 => "0001101111000000001100",
			4958 => "0000011101111100001000",
			4959 => "0000011101111100000100",
			4960 => "0000000100111000000011",
			4961 => "0000001100111000000011",
			4962 => "0000000100111000000011",
			4963 => "0000000100111000000011",
			4964 => "0001101000010000000100",
			4965 => "0000000100111000000011",
			4966 => "0000011101111100000100",
			4967 => "0000000100111000000011",
			4968 => "0001111000011000000100",
			4969 => "0000000100111000000011",
			4970 => "0000001100111000000011",
			4971 => "0000011100011000011100",
			4972 => "0000111100111000001100",
			4973 => "0010111011011100001000",
			4974 => "0010110000011100000100",
			4975 => "0000000100111000000011",
			4976 => "0000000100111000000011",
			4977 => "0000001100111000000011",
			4978 => "0000000111000000001000",
			4979 => "0010110100010000000100",
			4980 => "0000000100111000000011",
			4981 => "1111111100111000000011",
			4982 => "0010000001110000000100",
			4983 => "0000000100111000000011",
			4984 => "0000000100111000000011",
			4985 => "0001110000011100001100",
			4986 => "0010111011011100000100",
			4987 => "0000000100111000000011",
			4988 => "0010001001101000000100",
			4989 => "0000001100111000000011",
			4990 => "0000000100111000000011",
			4991 => "0000000100111000000011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1652, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3300, initial_addr_3'length));
	end generate gen_rom_10;

	gen_rom_11: if SELECT_ROM = 11 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000011101111100000100",
			29 => "0000000000000001111101",
			30 => "0000000000000001111101",
			31 => "0010001100011100000100",
			32 => "0000000000000010001001",
			33 => "0000000000000010001001",
			34 => "0000101011111000001000",
			35 => "0011100110010000000100",
			36 => "0000000000000010011101",
			37 => "0000000000000010011101",
			38 => "0000000000000010011101",
			39 => "0010010111101100001000",
			40 => "0000000110001000000100",
			41 => "0000000000000010110001",
			42 => "0000000000000010110001",
			43 => "0000000000000010110001",
			44 => "0000010111101000001000",
			45 => "0010010111101100000100",
			46 => "0000000000000011000101",
			47 => "0000000000000011000101",
			48 => "0000000000000011000101",
			49 => "0010010000001000001000",
			50 => "0000011101111100000100",
			51 => "0000000000000011011001",
			52 => "0000000000000011011001",
			53 => "0000000000000011011001",
			54 => "0010000001010100001100",
			55 => "0000011011111100000100",
			56 => "0000000000000011110101",
			57 => "0000011100011000000100",
			58 => "0000000000000011110101",
			59 => "0000000000000011110101",
			60 => "0000000000000011110101",
			61 => "0000010100110100001100",
			62 => "0011100110010000000100",
			63 => "0000000000000100010001",
			64 => "0001000011001100000100",
			65 => "0000000000000100010001",
			66 => "0000000000000100010001",
			67 => "0000000000000100010001",
			68 => "0010011001111100001000",
			69 => "0001001100010000000100",
			70 => "0000000000000100111101",
			71 => "0000000000000100111101",
			72 => "0011101100000000001000",
			73 => "0001001111100100000100",
			74 => "0000000000000100111101",
			75 => "0000000000000100111101",
			76 => "0001001111101000000100",
			77 => "0000000000000100111101",
			78 => "0000000000000100111101",
			79 => "0011100110010000001100",
			80 => "0010010101010000000100",
			81 => "0000000000000101101001",
			82 => "0000001100000100000100",
			83 => "0000000000000101101001",
			84 => "0000000000000101101001",
			85 => "0010010111101100001000",
			86 => "0011011110101100000100",
			87 => "0000000000000101101001",
			88 => "0000000000000101101001",
			89 => "0000000000000101101001",
			90 => "0000011110010100000100",
			91 => "0000000000000110001101",
			92 => "0010011010100100001100",
			93 => "0010000001110000001000",
			94 => "0010001010110000000100",
			95 => "0000000000000110001101",
			96 => "0000000000000110001101",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0011100110010000000100",
			100 => "0000000000000110110001",
			101 => "0000011101111100001100",
			102 => "0011001011000000001000",
			103 => "0011000100001000000100",
			104 => "0000000000000110110001",
			105 => "0000000000000110110001",
			106 => "0000000000000110110001",
			107 => "0000000000000110110001",
			108 => "0010010111101100001000",
			109 => "0010110100000100000100",
			110 => "0000000000000111011101",
			111 => "0000000000000111011101",
			112 => "0011001010111000000100",
			113 => "0000000000000111011101",
			114 => "0011011111010000001000",
			115 => "0010101000010100000100",
			116 => "0000000000000111011101",
			117 => "0000000000000111011101",
			118 => "0000000000000111011101",
			119 => "0010010111101100001100",
			120 => "0000101000001100001000",
			121 => "0010001010110000000100",
			122 => "0000000000001000010001",
			123 => "0000000000001000010001",
			124 => "0000000000001000010001",
			125 => "0001101111000000001000",
			126 => "0011001011000000000100",
			127 => "0000000000001000010001",
			128 => "0000000000001000010001",
			129 => "0000101100111000000100",
			130 => "0000000000001000010001",
			131 => "0000000000001000010001",
			132 => "0000011110010100001000",
			133 => "0000001001101000000100",
			134 => "0000000000001001000101",
			135 => "0000000000001001000101",
			136 => "0011010111111100010000",
			137 => "0001000001011100000100",
			138 => "0000000000001001000101",
			139 => "0011101011111000001000",
			140 => "0000000110001000000100",
			141 => "0000000000001001000101",
			142 => "0000000000001001000101",
			143 => "0000000000001001000101",
			144 => "0000000000001001000101",
			145 => "0000101010000100010000",
			146 => "0011001000000000001100",
			147 => "0011100010000000000100",
			148 => "0000000000001010001001",
			149 => "0001101001100100000100",
			150 => "0000000000001010001001",
			151 => "0000000000001010001001",
			152 => "0000000000001010001001",
			153 => "0011111000001100001100",
			154 => "0001001011101100000100",
			155 => "0000000000001010001001",
			156 => "0010101000010100000100",
			157 => "0000000000001010001001",
			158 => "0000000000001010001001",
			159 => "0001000010010100000100",
			160 => "0000000000001010001001",
			161 => "0000000000001010001001",
			162 => "0000010100110100011000",
			163 => "0011100110010000010000",
			164 => "0011101110101000000100",
			165 => "0000000000001010111101",
			166 => "0001101010011000000100",
			167 => "0000000000001010111101",
			168 => "0011110000010000000100",
			169 => "0000000000001010111101",
			170 => "0000000000001010111101",
			171 => "0001000011001100000100",
			172 => "0000000000001010111101",
			173 => "0000000000001010111101",
			174 => "0000000000001010111101",
			175 => "0011001010111000011000",
			176 => "0011011100100100001100",
			177 => "0000011011111100000100",
			178 => "0000000000001100011001",
			179 => "0010000001110000000100",
			180 => "0000000000001100011001",
			181 => "0000000000001100011001",
			182 => "0001001101101100001000",
			183 => "0001010010110100000100",
			184 => "0000000000001100011001",
			185 => "1111111000001100011001",
			186 => "0000000000001100011001",
			187 => "0011010010011100010000",
			188 => "0010011001111100000100",
			189 => "0000000000001100011001",
			190 => "0001000001011100000100",
			191 => "0000000000001100011001",
			192 => "0011101011111000000100",
			193 => "0000000000001100011001",
			194 => "0000000000001100011001",
			195 => "0011101111010100000100",
			196 => "0000000000001100011001",
			197 => "0000000000001100011001",
			198 => "0000011110010100001100",
			199 => "0010010100101100001000",
			200 => "0001001100010000000100",
			201 => "0000000000001101011101",
			202 => "0000000000001101011101",
			203 => "0000000000001101011101",
			204 => "0011010111111100010100",
			205 => "0001000001011100000100",
			206 => "0000000000001101011101",
			207 => "0011101011111000001100",
			208 => "0001100100111100001000",
			209 => "0000000110001000000100",
			210 => "0000000000001101011101",
			211 => "0000000000001101011101",
			212 => "0000000000001101011101",
			213 => "0000000000001101011101",
			214 => "0000000000001101011101",
			215 => "0000101011111000011000",
			216 => "0010100111110100010100",
			217 => "0000111111010100010000",
			218 => "0001001111100100001000",
			219 => "0000111110110100000100",
			220 => "0000000000001110110001",
			221 => "0000000000001110110001",
			222 => "0011110110010000000100",
			223 => "0000000000001110110001",
			224 => "0000000000001110110001",
			225 => "0000000000001110110001",
			226 => "1111111000001110110001",
			227 => "0000111011111000001100",
			228 => "0001100100111100001000",
			229 => "0000010001000100000100",
			230 => "0000000000001110110001",
			231 => "0000000000001110110001",
			232 => "0000000000001110110001",
			233 => "0000011101111100000100",
			234 => "0000000000001110110001",
			235 => "0000000000001110110001",
			236 => "0000101100000000000100",
			237 => "0000000000001111100101",
			238 => "0000101111101000010100",
			239 => "0000010001000100000100",
			240 => "0000000000001111100101",
			241 => "0000011100011000001100",
			242 => "0001101101011000000100",
			243 => "0000000000001111100101",
			244 => "0001101000010000000100",
			245 => "0000000000001111100101",
			246 => "0000000000001111100101",
			247 => "0000000000001111100101",
			248 => "0000000000001111100101",
			249 => "0011001010111100001100",
			250 => "0000010111101000001000",
			251 => "0010000001010000000100",
			252 => "0000000000010001000001",
			253 => "0000000000010001000001",
			254 => "0000000000010001000001",
			255 => "0011101110110100001100",
			256 => "0010101010100000000100",
			257 => "0000000000010001000001",
			258 => "0010010101010000000100",
			259 => "0000000000010001000001",
			260 => "0000000000010001000001",
			261 => "0001000011000000001100",
			262 => "0010011010100000001000",
			263 => "0000010001111000000100",
			264 => "0000000000010001000001",
			265 => "0000000000010001000001",
			266 => "0000000000010001000001",
			267 => "0000111111100100001000",
			268 => "0000010111101000000100",
			269 => "0000000000010001000001",
			270 => "0000000000010001000001",
			271 => "0000000000010001000001",
			272 => "0011001010111000010000",
			273 => "0010001100011100000100",
			274 => "0000000000010010100101",
			275 => "0010010000001000001000",
			276 => "0001111001001000000100",
			277 => "1111111000010010100101",
			278 => "0000000000010010100101",
			279 => "0000000000010010100101",
			280 => "0011000100011000010000",
			281 => "0000001111001000000100",
			282 => "0000000000010010100101",
			283 => "0010000001010100001000",
			284 => "0011101011111000000100",
			285 => "0000000000010010100101",
			286 => "0000000000010010100101",
			287 => "0000000000010010100101",
			288 => "0011101100010000001000",
			289 => "0000011110010100000100",
			290 => "0000000000010010100101",
			291 => "0000000000010010100101",
			292 => "0001001011110000001000",
			293 => "0010001010110000000100",
			294 => "0000000000010010100101",
			295 => "1111111000010010100101",
			296 => "0000000000010010100101",
			297 => "0011001010111100010000",
			298 => "0000010111101000001100",
			299 => "0000001011010100000100",
			300 => "0000000000010100001001",
			301 => "0001111000000000000100",
			302 => "0000000000010100001001",
			303 => "0000000000010100001001",
			304 => "0000000000010100001001",
			305 => "0001111001001000001100",
			306 => "0010011010100000001000",
			307 => "0000010001000100000100",
			308 => "0000000000010100001001",
			309 => "0000000000010100001001",
			310 => "0000000000010100001001",
			311 => "0011101100010000001100",
			312 => "0000101100000000000100",
			313 => "0000000000010100001001",
			314 => "0000011110010100000100",
			315 => "0000000000010100001001",
			316 => "0000000000010100001001",
			317 => "0000011101111100001000",
			318 => "0011001000000000000100",
			319 => "0000000000010100001001",
			320 => "0000000000010100001001",
			321 => "0000000000010100001001",
			322 => "0000101010000100001100",
			323 => "0010001010110000000100",
			324 => "0000000000010101100101",
			325 => "0001101001100100000100",
			326 => "0000000000010101100101",
			327 => "0000000000010101100101",
			328 => "0011101100010000001000",
			329 => "0010010101010000000100",
			330 => "0000000000010101100101",
			331 => "0000000000010101100101",
			332 => "0010010000001000010000",
			333 => "0011001000000000001100",
			334 => "0011010001000000000100",
			335 => "0000000000010101100101",
			336 => "0000011101111100000100",
			337 => "0000000000010101100101",
			338 => "0000000000010101100101",
			339 => "0000000000010101100101",
			340 => "0010110101100100001000",
			341 => "0010101000010100000100",
			342 => "0000000000010101100101",
			343 => "0000000000010101100101",
			344 => "0000000000010101100101",
			345 => "0000011011111100001000",
			346 => "0001101001100100000100",
			347 => "0000000000010111000001",
			348 => "0000000000010111000001",
			349 => "0011101100000000001100",
			350 => "0001001111100100000100",
			351 => "0000000000010111000001",
			352 => "0011001011000000000100",
			353 => "0000000000010111000001",
			354 => "0000000000010111000001",
			355 => "0001000010010100001100",
			356 => "0000011101111100001000",
			357 => "0011110111010100000100",
			358 => "0000000000010111000001",
			359 => "0000000000010111000001",
			360 => "0000000000010111000001",
			361 => "0011010111111100001100",
			362 => "0000000111000000001000",
			363 => "0011111000101000000100",
			364 => "0000000000010111000001",
			365 => "0000000000010111000001",
			366 => "0000000000010111000001",
			367 => "0000000000010111000001",
			368 => "0000101011111000011000",
			369 => "0010100111110100010100",
			370 => "0011101100010000001100",
			371 => "0001001111100100000100",
			372 => "0000000000011000101101",
			373 => "0011110110010000000100",
			374 => "0000000000011000101101",
			375 => "0000000000011000101101",
			376 => "0001001000101000000100",
			377 => "0000000000011000101101",
			378 => "0000000000011000101101",
			379 => "1111111000011000101101",
			380 => "0000111011111000010100",
			381 => "0001100100111100010000",
			382 => "0011010010011100001100",
			383 => "0001110111001000000100",
			384 => "0000000000011000101101",
			385 => "0001101011001100000100",
			386 => "0000000000011000101101",
			387 => "0000001000011000101101",
			388 => "0000000000011000101101",
			389 => "0000000000011000101101",
			390 => "0010110111010000000100",
			391 => "0000000000011000101101",
			392 => "0001111000011000000100",
			393 => "0000000000011000101101",
			394 => "0000000000011000101101",
			395 => "0000100110111100010000",
			396 => "0011111111010100001100",
			397 => "0001101001100100001000",
			398 => "0001001100010000000100",
			399 => "0000000000011010001001",
			400 => "0000000000011010001001",
			401 => "0000000000011010001001",
			402 => "0000000000011010001001",
			403 => "0001000001011100001000",
			404 => "0011111000001100000100",
			405 => "0000000000011010001001",
			406 => "0000000000011010001001",
			407 => "0011110011000000010100",
			408 => "0001101101011000000100",
			409 => "0000000000011010001001",
			410 => "0011000100001000000100",
			411 => "0000000000011010001001",
			412 => "0001100100111100001000",
			413 => "0000010001000100000100",
			414 => "0000000000011010001001",
			415 => "0000000000011010001001",
			416 => "0000000000011010001001",
			417 => "0000000000011010001001",
			418 => "0011001010111000011000",
			419 => "0011011100100100001100",
			420 => "0000011011111100000100",
			421 => "0000000000011011111101",
			422 => "0000100011000000000100",
			423 => "0000000000011011111101",
			424 => "0000000000011011111101",
			425 => "0001001101101100001000",
			426 => "0000111001100000000100",
			427 => "0000000000011011111101",
			428 => "1111111000011011111101",
			429 => "0000000000011011111101",
			430 => "0011010010011100011100",
			431 => "0010011001111100000100",
			432 => "0000000000011011111101",
			433 => "0000101010000100001100",
			434 => "0011100110010000000100",
			435 => "0000000000011011111101",
			436 => "0010001010110000000100",
			437 => "0000000000011011111101",
			438 => "0000000000011011111101",
			439 => "0011101011111000001000",
			440 => "0000000110001000000100",
			441 => "0000000000011011111101",
			442 => "0000000000011011111101",
			443 => "0000000000011011111101",
			444 => "0011101111010100000100",
			445 => "0000000000011011111101",
			446 => "0000000000011011111101",
			447 => "0010011001111100000100",
			448 => "0000000000011100111001",
			449 => "0011010111111100011000",
			450 => "0011001010111000000100",
			451 => "0000000000011100111001",
			452 => "0001100100111100010000",
			453 => "0011101011111000001100",
			454 => "0011001000000000001000",
			455 => "0010010111101100000100",
			456 => "0000000000011100111001",
			457 => "0000000000011100111001",
			458 => "0000000000011100111001",
			459 => "0000000000011100111001",
			460 => "0000000000011100111001",
			461 => "0000000000011100111001",
			462 => "0000010001000100000100",
			463 => "0000000000011101110101",
			464 => "0010110101100100011000",
			465 => "0010101010100100000100",
			466 => "0000000000011101110101",
			467 => "0011001011000000010000",
			468 => "0001110001101000001100",
			469 => "0010011010100100001000",
			470 => "0011101011111000000100",
			471 => "0000000000011101110101",
			472 => "0000000000011101110101",
			473 => "0000000000011101110101",
			474 => "0000000000011101110101",
			475 => "0000000000011101110101",
			476 => "0000000000011101110101",
			477 => "0000011011111100001000",
			478 => "0010011001111100000100",
			479 => "1111111000011111100001",
			480 => "0000000000011111100001",
			481 => "0011100110111100010000",
			482 => "0001001111100100001000",
			483 => "0011100110010000000100",
			484 => "0000000000011111100001",
			485 => "1111111000011111100001",
			486 => "0011001011000000000100",
			487 => "0000001000011111100001",
			488 => "0000000000011111100001",
			489 => "0010010000001000001000",
			490 => "0011011110101000000100",
			491 => "0000000000011111100001",
			492 => "1111111000011111100001",
			493 => "0011010101001000001000",
			494 => "0000000111000000000100",
			495 => "0000001000011111100001",
			496 => "0000000000011111100001",
			497 => "0010011010100000001000",
			498 => "0010110110110100000100",
			499 => "0000000000011111100001",
			500 => "0000000000011111100001",
			501 => "0010110000011100000100",
			502 => "0000000000011111100001",
			503 => "1111111000011111100001",
			504 => "0011001010111000010000",
			505 => "0000000111000100000100",
			506 => "0000000000100001011101",
			507 => "0010010000001000001000",
			508 => "0001111001001000000100",
			509 => "1111111000100001011101",
			510 => "0000000000100001011101",
			511 => "0000000000100001011101",
			512 => "0001110110100100010100",
			513 => "0011010101001000010000",
			514 => "0000101100000000000100",
			515 => "0000000000100001011101",
			516 => "0010010100101100000100",
			517 => "0000000000100001011101",
			518 => "0011101011111000000100",
			519 => "0000000000100001011101",
			520 => "0000000000100001011101",
			521 => "0000000000100001011101",
			522 => "0001111000011000001100",
			523 => "0011101100010000000100",
			524 => "0000000000100001011101",
			525 => "0010110110110100000100",
			526 => "0000000000100001011101",
			527 => "0000000000100001011101",
			528 => "0001011110000100001100",
			529 => "0011111100111000001000",
			530 => "0000101010000100000100",
			531 => "0000000000100001011101",
			532 => "0000000000100001011101",
			533 => "0000000000100001011101",
			534 => "0000000000100001011101",
			535 => "0010010101010000000100",
			536 => "1111111000100011000001",
			537 => "0001000010010100100000",
			538 => "0011100110111100010100",
			539 => "0001001111100100001000",
			540 => "0011100010000000000100",
			541 => "0000000000100011000001",
			542 => "0000000000100011000001",
			543 => "0011001011000000000100",
			544 => "0000001000100011000001",
			545 => "0000001111001000000100",
			546 => "0000000000100011000001",
			547 => "0000000000100011000001",
			548 => "0011110000010000000100",
			549 => "0000000000100011000001",
			550 => "0001000010010100000100",
			551 => "1111111000100011000001",
			552 => "0000000000100011000001",
			553 => "0011101011111000001100",
			554 => "0011010010011100001000",
			555 => "0001101000010000000100",
			556 => "0000001000100011000001",
			557 => "0000000000100011000001",
			558 => "0000000000100011000001",
			559 => "0000000000100011000001",
			560 => "0000010001000100000100",
			561 => "1111111000100100000101",
			562 => "0011101011111000011100",
			563 => "0010000001110000011000",
			564 => "0011011001010000010000",
			565 => "0010101010100100000100",
			566 => "1111111000100100000101",
			567 => "0000000111000000001000",
			568 => "0011001011000000000100",
			569 => "0000001000100100000101",
			570 => "0000000000100100000101",
			571 => "0000010000100100000101",
			572 => "0000101111100100000100",
			573 => "1111111000100100000101",
			574 => "0000001000100100000101",
			575 => "1111111000100100000101",
			576 => "1111111000100100000101",
			577 => "0010000001110000101100",
			578 => "0000111011111000100100",
			579 => "0001001100111000010100",
			580 => "0011100110010000001000",
			581 => "0000011011111100000100",
			582 => "0000000000100101100001",
			583 => "0000000000100101100001",
			584 => "0010111011011100001000",
			585 => "0010110111010000000100",
			586 => "0000000000100101100001",
			587 => "0000000000100101100001",
			588 => "0000000000100101100001",
			589 => "0000010001000100000100",
			590 => "0000000000100101100001",
			591 => "0001100100111100001000",
			592 => "0010001010110000000100",
			593 => "0000000000100101100001",
			594 => "0000001000100101100001",
			595 => "0000000000100101100001",
			596 => "0000010100110100000100",
			597 => "0000000000100101100001",
			598 => "0000000000100101100001",
			599 => "1111111000100101100001",
			600 => "0010000001110000101100",
			601 => "0000111011111000100100",
			602 => "0001001100111000010000",
			603 => "0011100110010000001000",
			604 => "0000011011111100000100",
			605 => "0000000000100110111101",
			606 => "0000000000100110111101",
			607 => "0000000110001000000100",
			608 => "0000000000100110111101",
			609 => "0000000000100110111101",
			610 => "0000010001000100000100",
			611 => "0000000000100110111101",
			612 => "0001100100111100001100",
			613 => "0010001010110000000100",
			614 => "0000000000100110111101",
			615 => "0011010010011100000100",
			616 => "0000001000100110111101",
			617 => "0000000000100110111101",
			618 => "0000000000100110111101",
			619 => "0000010100110100000100",
			620 => "0000000000100110111101",
			621 => "0000000000100110111101",
			622 => "1111111000100110111101",
			623 => "0011001010111000100100",
			624 => "0000101000001100010100",
			625 => "0010100111110100010000",
			626 => "0010111010001100000100",
			627 => "0000000000101001001001",
			628 => "0001111000000000000100",
			629 => "0000000000101001001001",
			630 => "0010110000011100000100",
			631 => "0000000000101001001001",
			632 => "0000000000101001001001",
			633 => "1111111000101001001001",
			634 => "0011101010000100001100",
			635 => "0010111001001000000100",
			636 => "0000000000101001001001",
			637 => "0000101100111000000100",
			638 => "0000000000101001001001",
			639 => "0000000000101001001001",
			640 => "0000000000101001001001",
			641 => "0010010111101100001100",
			642 => "0011000100011000000100",
			643 => "0000000000101001001001",
			644 => "0011001000000000000100",
			645 => "0000000000101001001001",
			646 => "0000000000101001001001",
			647 => "0000101111010100000100",
			648 => "0000000000101001001001",
			649 => "0011101111010100000100",
			650 => "0000000000101001001001",
			651 => "0001001011110000000100",
			652 => "0000000000101001001001",
			653 => "0001110001101000001000",
			654 => "0001000101000000000100",
			655 => "0000000000101001001001",
			656 => "0000000000101001001001",
			657 => "0000000000101001001001",
			658 => "0000011011111100000100",
			659 => "1111111000101010010101",
			660 => "0000111111100100100000",
			661 => "0011100110010000000100",
			662 => "0000001000101010010101",
			663 => "0010100011101000001000",
			664 => "0001111001001000000100",
			665 => "0000000000101010010101",
			666 => "1111111000101010010101",
			667 => "0000010111101000001000",
			668 => "0001101001100100000100",
			669 => "0000000000101010010101",
			670 => "1111111000101010010101",
			671 => "0010011010100100001000",
			672 => "0000000110001000000100",
			673 => "0000000000101010010101",
			674 => "0000001000101010010101",
			675 => "1111111000101010010101",
			676 => "1111111000101010010101",
			677 => "0000010001000100000100",
			678 => "1111111000101100011001",
			679 => "0011100110111100100000",
			680 => "0010110100000100001100",
			681 => "0001001011101100001000",
			682 => "0011100110010000000100",
			683 => "0000001000101100011001",
			684 => "1111111000101100011001",
			685 => "0000001000101100011001",
			686 => "0001000001011100001100",
			687 => "0011100110010000000100",
			688 => "0000001000101100011001",
			689 => "0001010110100000000100",
			690 => "0000000000101100011001",
			691 => "1111111000101100011001",
			692 => "0000100110101100000100",
			693 => "0000001000101100011001",
			694 => "0000000000101100011001",
			695 => "0001110110100100001100",
			696 => "0001000010010100000100",
			697 => "1111111000101100011001",
			698 => "0011101011111000000100",
			699 => "0000001000101100011001",
			700 => "0000000000101100011001",
			701 => "0001000011000000001000",
			702 => "0010000110011100000100",
			703 => "1111111000101100011001",
			704 => "1111110000101100011001",
			705 => "0011111100111000001000",
			706 => "0001000010010100000100",
			707 => "0000000000101100011001",
			708 => "0000001000101100011001",
			709 => "1111111000101100011001",
			710 => "0010010101010000001100",
			711 => "0010010101010000000100",
			712 => "1111111000101110001101",
			713 => "0010010101010000000100",
			714 => "0000000000101110001101",
			715 => "1111111000101110001101",
			716 => "0011011001010000100100",
			717 => "0010000001110000100000",
			718 => "0000101101101100011100",
			719 => "0011010101001000010000",
			720 => "0011000100011000001000",
			721 => "0000101100111000000100",
			722 => "0000001000101110001101",
			723 => "0000010000101110001101",
			724 => "0000100111010100000100",
			725 => "0000000000101110001101",
			726 => "0000001000101110001101",
			727 => "0010100011101000000100",
			728 => "1111111000101110001101",
			729 => "0011100111010100000100",
			730 => "0000001000101110001101",
			731 => "1111111000101110001101",
			732 => "0000011000101110001101",
			733 => "1111111000101110001101",
			734 => "0011101111010100001000",
			735 => "0010010100101100000100",
			736 => "1111111000101110001101",
			737 => "0000001000101110001101",
			738 => "1111111000101110001101",
			739 => "0010011001111100010100",
			740 => "0000010001000100000100",
			741 => "1111111000110000110001",
			742 => "0010000001010100001100",
			743 => "0010001010110000001000",
			744 => "0000011011111100000100",
			745 => "0000000000110000110001",
			746 => "0000000000110000110001",
			747 => "0000000000110000110001",
			748 => "1111111000110000110001",
			749 => "0001110001101000100100",
			750 => "0000111011111000011000",
			751 => "0011001011000000010000",
			752 => "0000011101111100001000",
			753 => "0011101000001100000100",
			754 => "0000001000110000110001",
			755 => "0000000000110000110001",
			756 => "0000010100110100000100",
			757 => "0000000000110000110001",
			758 => "0000000000110000110001",
			759 => "0000010001111000000100",
			760 => "0000000000110000110001",
			761 => "0000000000110000110001",
			762 => "0000010100110100000100",
			763 => "1111111000110000110001",
			764 => "0001011110101000000100",
			765 => "0000000000110000110001",
			766 => "0000000000110000110001",
			767 => "0010000110011100001000",
			768 => "0000111010000100000100",
			769 => "0000000000110000110001",
			770 => "0000000000110000110001",
			771 => "0011001010111000000100",
			772 => "0000000000110000110001",
			773 => "0001000101000000000100",
			774 => "1111111000110000110001",
			775 => "0000010001111000001000",
			776 => "0000010001111000000100",
			777 => "0000000000110000110001",
			778 => "0000000000110000110001",
			779 => "0000000000110000110001",
			780 => "0000010001000100000100",
			781 => "1111111000110010010101",
			782 => "0011100110010000001000",
			783 => "0001101010011000000100",
			784 => "0000000000110010010101",
			785 => "0000001000110010010101",
			786 => "0001001100111000010100",
			787 => "0001000110101100000100",
			788 => "1111111000110010010101",
			789 => "0000111100000000000100",
			790 => "0000000000110010010101",
			791 => "0001101001100100001000",
			792 => "0001101011001100000100",
			793 => "0000000000110010010101",
			794 => "1111111000110010010101",
			795 => "0000000000110010010101",
			796 => "0011101011111000010000",
			797 => "0000010111101000000100",
			798 => "1111111000110010010101",
			799 => "0001000010010100001000",
			800 => "0011101111010100000100",
			801 => "0000001000110010010101",
			802 => "1111111000110010010101",
			803 => "0000001000110010010101",
			804 => "1111111000110010010101",
			805 => "0000010001000100000100",
			806 => "1111111000110100011001",
			807 => "0001111001001000010100",
			808 => "0001001100111000001100",
			809 => "0000001011010100000100",
			810 => "0000000000110100011001",
			811 => "0010001010110000000100",
			812 => "0000000000110100011001",
			813 => "0000000000110100011001",
			814 => "0011101000001100000100",
			815 => "0000001000110100011001",
			816 => "0000000000110100011001",
			817 => "0010010000001000010100",
			818 => "0011101100010000001100",
			819 => "0000001001101000000100",
			820 => "0000000000110100011001",
			821 => "0000001111001000000100",
			822 => "0000000000110100011001",
			823 => "0000000000110100011001",
			824 => "0011001101010100000100",
			825 => "0000000000110100011001",
			826 => "1111111000110100011001",
			827 => "0011000100011000010000",
			828 => "0000001111001000000100",
			829 => "0000000000110100011001",
			830 => "0010000001010100001000",
			831 => "0011101011111000000100",
			832 => "0000001000110100011001",
			833 => "0000000000110100011001",
			834 => "0000000000110100011001",
			835 => "0010000110011100000100",
			836 => "0000000000110100011001",
			837 => "0000000000110100011001",
			838 => "0010011001111100001000",
			839 => "0001001100000000000100",
			840 => "0000000000110110001101",
			841 => "1111111000110110001101",
			842 => "0001000010010100100100",
			843 => "0011011100100100000100",
			844 => "0000001000110110001101",
			845 => "0011001010111000000100",
			846 => "1111111000110110001101",
			847 => "0010000110011100010000",
			848 => "0011100110111100001000",
			849 => "0010001010110000000100",
			850 => "0000000000110110001101",
			851 => "0000001000110110001101",
			852 => "0001000011000000000100",
			853 => "0000000000110110001101",
			854 => "0000000000110110001101",
			855 => "0000001111001000000100",
			856 => "0000000000110110001101",
			857 => "0011000100011000000100",
			858 => "0000000000110110001101",
			859 => "0000000000110110001101",
			860 => "0011010111111100001100",
			861 => "0000010111101000000100",
			862 => "0000000000110110001101",
			863 => "0011101011111000000100",
			864 => "0000001000110110001101",
			865 => "0000000000110110001101",
			866 => "0000000000110110001101",
			867 => "0010000001010101000000",
			868 => "0011011111010000100000",
			869 => "0001101010011000000100",
			870 => "1111111000111000110001",
			871 => "0011001011000000011000",
			872 => "0001000011000000010000",
			873 => "0011101100000000001000",
			874 => "0000111100010000000100",
			875 => "0000001000111000110001",
			876 => "0000001000111000110001",
			877 => "0000101000001100000100",
			878 => "0000000000111000110001",
			879 => "1111111000111000110001",
			880 => "0000101100111000000100",
			881 => "0000001000111000110001",
			882 => "0000001000111000110001",
			883 => "0000000000111000110001",
			884 => "0001010110100000001000",
			885 => "0000000001010100000100",
			886 => "1111111000111000110001",
			887 => "0000001000111000110001",
			888 => "0011000100011000001100",
			889 => "0000000111000100000100",
			890 => "1111111000111000110001",
			891 => "0001101111000000000100",
			892 => "0000001000111000110001",
			893 => "0000000000111000110001",
			894 => "0001011100100100001000",
			895 => "0001011110101000000100",
			896 => "1111111000111000110001",
			897 => "0000000000111000110001",
			898 => "1111111000111000110001",
			899 => "0010000001110000010000",
			900 => "0011101000001100001100",
			901 => "0011000100001000000100",
			902 => "1111111000111000110001",
			903 => "0001000010110000000100",
			904 => "0000001000111000110001",
			905 => "0000001000111000110001",
			906 => "1111111000111000110001",
			907 => "1111111000111000110001",
			908 => "0000010001000100000100",
			909 => "1111111000111010111101",
			910 => "0001111001001000010100",
			911 => "0001001100111000001100",
			912 => "0000001011010100000100",
			913 => "0000000000111010111101",
			914 => "0010001010110000000100",
			915 => "0000000000111010111101",
			916 => "0000000000111010111101",
			917 => "0011101000001100000100",
			918 => "0000001000111010111101",
			919 => "0000000000111010111101",
			920 => "0010010000001000011000",
			921 => "0011101100010000010000",
			922 => "0000001001101000000100",
			923 => "0000000000111010111101",
			924 => "0000001111001000001000",
			925 => "0000101100000000000100",
			926 => "0000000000111010111101",
			927 => "0000000000111010111101",
			928 => "0000000000111010111101",
			929 => "0011001101010100000100",
			930 => "0000000000111010111101",
			931 => "1111111000111010111101",
			932 => "0011000100011000010000",
			933 => "0000001111001000000100",
			934 => "0000000000111010111101",
			935 => "0010000001010100001000",
			936 => "0011101011111000000100",
			937 => "0000001000111010111101",
			938 => "0000000000111010111101",
			939 => "0000000000111010111101",
			940 => "0010000110011100000100",
			941 => "0000000000111010111101",
			942 => "0000000000111010111101",
			943 => "0000010001000100000100",
			944 => "1111111000111100011001",
			945 => "0000111011101100101000",
			946 => "0000111100010000000100",
			947 => "0000001000111100011001",
			948 => "0001001011101100001100",
			949 => "0011110110111100001000",
			950 => "0000101100000000000100",
			951 => "1111111000111100011001",
			952 => "0000000000111100011001",
			953 => "1111111000111100011001",
			954 => "0000010111101000001000",
			955 => "0001010010110100000100",
			956 => "0000000000111100011001",
			957 => "1111111000111100011001",
			958 => "0001000011000000001000",
			959 => "0001101001100100000100",
			960 => "0000000000111100011001",
			961 => "1111111000111100011001",
			962 => "0001101000010000000100",
			963 => "0000001000111100011001",
			964 => "0000000000111100011001",
			965 => "1111111000111100011001",
			966 => "0000010001000100000100",
			967 => "1111111000111110001101",
			968 => "0011100110010000001000",
			969 => "0001101010011000000100",
			970 => "0000000000111110001101",
			971 => "0000001000111110001101",
			972 => "0001001100111000011000",
			973 => "0001001111100100000100",
			974 => "1111111000111110001101",
			975 => "0000111100000000001000",
			976 => "0010010000001000000100",
			977 => "0000000000111110001101",
			978 => "0000000000111110001101",
			979 => "0001101001100100001000",
			980 => "0001101011001100000100",
			981 => "0000000000111110001101",
			982 => "1111111000111110001101",
			983 => "0000000000111110001101",
			984 => "0011101011111000010100",
			985 => "0000010111101000000100",
			986 => "1111111000111110001101",
			987 => "0001000010010100001000",
			988 => "0011101111010100000100",
			989 => "0000001000111110001101",
			990 => "1111111000111110001101",
			991 => "0001100100111100000100",
			992 => "0000001000111110001101",
			993 => "0000000000111110001101",
			994 => "1111111000111110001101",
			995 => "0000010001000100000100",
			996 => "1111111001000000100001",
			997 => "0001111001001000011100",
			998 => "0001000011001100010100",
			999 => "0000111100010000000100",
			1000 => "0000001001000000100001",
			1001 => "0001001011101100000100",
			1002 => "1111111001000000100001",
			1003 => "0011101011111000001000",
			1004 => "0001001101101100000100",
			1005 => "0000000001000000100001",
			1006 => "0000001001000000100001",
			1007 => "0000000001000000100001",
			1008 => "0001001010110100000100",
			1009 => "0000010001000000100001",
			1010 => "0000000001000000100001",
			1011 => "0011100110111100010100",
			1012 => "0010100011101000001000",
			1013 => "0000111100010000000100",
			1014 => "0000000001000000100001",
			1015 => "1111111001000000100001",
			1016 => "0010010100101100000100",
			1017 => "0000000001000000100001",
			1018 => "0000100111011000000100",
			1019 => "0000000001000000100001",
			1020 => "0000001001000000100001",
			1021 => "0000110111010100000100",
			1022 => "1111111001000000100001",
			1023 => "0001011100100100010000",
			1024 => "0001110110100100001000",
			1025 => "0000111111100100000100",
			1026 => "0000000001000000100001",
			1027 => "0000000001000000100001",
			1028 => "0010111011011100000100",
			1029 => "0000000001000000100001",
			1030 => "0000000001000000100001",
			1031 => "1111111001000000100001",
			1032 => "0000010001000100000100",
			1033 => "1111111001000010101101",
			1034 => "0011100110010000001000",
			1035 => "0001101010011000000100",
			1036 => "0000000001000010101101",
			1037 => "0000001001000010101101",
			1038 => "0000010111101000010000",
			1039 => "0010010111101100001100",
			1040 => "0001110110100100000100",
			1041 => "1111111001000010101101",
			1042 => "0011000100011000000100",
			1043 => "0000000001000010101101",
			1044 => "0000000001000010101101",
			1045 => "0000000001000010101101",
			1046 => "0001110001101000010100",
			1047 => "0001000010010100001100",
			1048 => "0011100110111100001000",
			1049 => "0001001111100100000100",
			1050 => "1111111001000010101101",
			1051 => "0000001001000010101101",
			1052 => "1111111001000010101101",
			1053 => "0011101011111000000100",
			1054 => "0000001001000010101101",
			1055 => "0000000001000010101101",
			1056 => "0011000100011000001100",
			1057 => "0000001111001000000100",
			1058 => "0000000001000010101101",
			1059 => "0010011010100100000100",
			1060 => "0000001001000010101101",
			1061 => "0000000001000010101101",
			1062 => "0010001100011100000100",
			1063 => "0000000001000010101101",
			1064 => "0001000101000000000100",
			1065 => "1111111001000010101101",
			1066 => "0000000001000010101101",
			1067 => "0000010001000100000100",
			1068 => "1111111001000100100011",
			1069 => "0011101011111000110100",
			1070 => "0010000001110000110000",
			1071 => "0001000001011100011100",
			1072 => "0011101110110100001100",
			1073 => "0000011011111100000100",
			1074 => "1111111001000100100011",
			1075 => "0000011101111100000100",
			1076 => "0000001001000100100011",
			1077 => "0000000001000100100011",
			1078 => "0001001011101100001000",
			1079 => "0010100011101000000100",
			1080 => "1111111001000100100011",
			1081 => "1111110001000100100011",
			1082 => "0011000100011000000100",
			1083 => "0000001001000100100011",
			1084 => "1111111001000100100011",
			1085 => "0000101101101100010000",
			1086 => "0011011111010000001000",
			1087 => "0011111111100100000100",
			1088 => "0000001001000100100011",
			1089 => "0000001001000100100011",
			1090 => "0011111111100100000100",
			1091 => "0000000001000100100011",
			1092 => "0000000001000100100011",
			1093 => "0000010001000100100011",
			1094 => "1111111001000100100011",
			1095 => "1111111001000100100011",
			1096 => "0000000001000100100101",
			1097 => "0000000001000100101001",
			1098 => "0000000001000100101101",
			1099 => "0000000001000100110001",
			1100 => "0000000001000100110101",
			1101 => "0000000001000100111001",
			1102 => "0000000001000100111101",
			1103 => "0000000001000101000001",
			1104 => "0000000001000101000101",
			1105 => "0000000001000101001001",
			1106 => "0000000001000101001101",
			1107 => "0000000001000101010001",
			1108 => "0000000001000101010101",
			1109 => "0000000001000101011001",
			1110 => "0000000001000101011101",
			1111 => "0000000001000101100001",
			1112 => "0000000001000101100101",
			1113 => "0000000001000101101001",
			1114 => "0000000001000101101101",
			1115 => "0000000001000101110001",
			1116 => "0000000001000101110101",
			1117 => "0000000001000101111001",
			1118 => "0000000001000101111101",
			1119 => "0000000001000110000001",
			1120 => "0000000001000110000101",
			1121 => "0000000001000110001001",
			1122 => "0000000001000110001101",
			1123 => "0010000001010100000100",
			1124 => "0000000001000110011001",
			1125 => "0000000001000110011001",
			1126 => "0010001100011100000100",
			1127 => "0000000001000110100101",
			1128 => "0000000001000110100101",
			1129 => "0000011101111100000100",
			1130 => "0000000001000110110001",
			1131 => "0000000001000110110001",
			1132 => "0011100110010000001000",
			1133 => "0011100101001000000100",
			1134 => "0000000001000111000101",
			1135 => "0000000001000111000101",
			1136 => "0000000001000111000101",
			1137 => "0010000001010100001000",
			1138 => "0001000011000000000100",
			1139 => "0000000001000111011001",
			1140 => "0000000001000111011001",
			1141 => "0000000001000111011001",
			1142 => "0011101100000000000100",
			1143 => "0000000001000111101101",
			1144 => "0011111000001100000100",
			1145 => "0000000001000111101101",
			1146 => "0000000001000111101101",
			1147 => "0000011011111100000100",
			1148 => "0000000001001000001001",
			1149 => "0000011100011000001000",
			1150 => "0000011110010100000100",
			1151 => "0000000001001000001001",
			1152 => "0000000001001000001001",
			1153 => "0000000001001000001001",
			1154 => "0010000001010100001100",
			1155 => "0000011011111100000100",
			1156 => "0000000001001000100101",
			1157 => "0010011010100100000100",
			1158 => "0000000001001000100101",
			1159 => "0000000001001000100101",
			1160 => "0000000001001000100101",
			1161 => "0000010111101000001000",
			1162 => "0010010111101100000100",
			1163 => "0000000001001001001001",
			1164 => "0000000001001001001001",
			1165 => "0000101010000100000100",
			1166 => "0000000001001001001001",
			1167 => "0000101111101000000100",
			1168 => "0000000001001001001001",
			1169 => "0000000001001001001001",
			1170 => "0011100110010000001100",
			1171 => "0010010101010000000100",
			1172 => "0000000001001001110101",
			1173 => "0000001100000100000100",
			1174 => "0000000001001001110101",
			1175 => "0000000001001001110101",
			1176 => "0000010100110100001000",
			1177 => "0011000100001000000100",
			1178 => "0000000001001001110101",
			1179 => "0000000001001001110101",
			1180 => "0000000001001001110101",
			1181 => "0010011001111100000100",
			1182 => "0000000001001010011001",
			1183 => "0001100100111100001100",
			1184 => "0001101010011000000100",
			1185 => "0000000001001010011001",
			1186 => "0010011010100100000100",
			1187 => "0000000001001010011001",
			1188 => "0000000001001010011001",
			1189 => "0000000001001010011001",
			1190 => "0000011110010100000100",
			1191 => "0000000001001010111101",
			1192 => "0010011010100100001100",
			1193 => "0010000001110000001000",
			1194 => "0010001010110000000100",
			1195 => "0000000001001010111101",
			1196 => "0000000001001010111101",
			1197 => "0000000001001010111101",
			1198 => "0000000001001010111101",
			1199 => "0010010000001000010000",
			1200 => "0011100110010000000100",
			1201 => "0000000001001011100001",
			1202 => "0001000011110000001000",
			1203 => "0000111100010000000100",
			1204 => "0000000001001011100001",
			1205 => "0000000001001011100001",
			1206 => "0000000001001011100001",
			1207 => "0000000001001011100001",
			1208 => "0010010111101100001000",
			1209 => "0010110100000100000100",
			1210 => "0000000001001100001101",
			1211 => "0000000001001100001101",
			1212 => "0011001010111000000100",
			1213 => "0000000001001100001101",
			1214 => "0011011111010000001000",
			1215 => "0010101000010100000100",
			1216 => "0000000001001100001101",
			1217 => "0000000001001100001101",
			1218 => "0000000001001100001101",
			1219 => "0011100110010000010000",
			1220 => "0011100101001000000100",
			1221 => "0000000001001101000001",
			1222 => "0011010001000000001000",
			1223 => "0000101011101100000100",
			1224 => "0000000001001101000001",
			1225 => "0000000001001101000001",
			1226 => "0000000001001101000001",
			1227 => "0001000011000000001000",
			1228 => "0011011110101000000100",
			1229 => "0000000001001101000001",
			1230 => "0000000001001101000001",
			1231 => "0000000001001101000001",
			1232 => "0010011001111100000100",
			1233 => "0000000001001101101101",
			1234 => "0001100100111100010000",
			1235 => "0001101010011000000100",
			1236 => "0000000001001101101101",
			1237 => "0010011010100100001000",
			1238 => "0000011110010100000100",
			1239 => "0000000001001101101101",
			1240 => "0000000001001101101101",
			1241 => "0000000001001101101101",
			1242 => "0000000001001101101101",
			1243 => "0010010111101100001100",
			1244 => "0010001010110000000100",
			1245 => "0000000001001110101001",
			1246 => "0011001010111100000100",
			1247 => "0000000001001110101001",
			1248 => "0000000001001110101001",
			1249 => "0010000101000100010000",
			1250 => "0011001010111000000100",
			1251 => "0000000001001110101001",
			1252 => "0010011010100100001000",
			1253 => "0011001011000000000100",
			1254 => "0000000001001110101001",
			1255 => "0000000001001110101001",
			1256 => "0000000001001110101001",
			1257 => "0000000001001110101001",
			1258 => "0010011001111100001000",
			1259 => "0001001100010000000100",
			1260 => "0000000001001111101101",
			1261 => "0000000001001111101101",
			1262 => "0011101100000000010000",
			1263 => "0001001111100100000100",
			1264 => "0000000001001111101101",
			1265 => "0010100011101000000100",
			1266 => "0000000001001111101101",
			1267 => "0010100111110100000100",
			1268 => "0000000001001111101101",
			1269 => "0000000001001111101101",
			1270 => "0001001111101000001000",
			1271 => "0011111000001100000100",
			1272 => "0000000001001111101101",
			1273 => "0000000001001111101101",
			1274 => "0000000001001111101101",
			1275 => "0000101000001100011100",
			1276 => "0011100110010000001100",
			1277 => "0000011011111100001000",
			1278 => "0000100111011000000100",
			1279 => "0000000001010001001001",
			1280 => "0000000001010001001001",
			1281 => "0000000001010001001001",
			1282 => "0001001101101100001100",
			1283 => "0010110101100100001000",
			1284 => "0011001000000000000100",
			1285 => "0000000001010001001001",
			1286 => "0000000001010001001001",
			1287 => "0000000001010001001001",
			1288 => "0000000001010001001001",
			1289 => "0011100111010100001100",
			1290 => "0010010101010000000100",
			1291 => "0000000001010001001001",
			1292 => "0001001000101000000100",
			1293 => "0000000001010001001001",
			1294 => "0000000001010001001001",
			1295 => "0000011101111100000100",
			1296 => "0000000001010001001001",
			1297 => "0000000001010001001001",
			1298 => "0010011001111100001000",
			1299 => "0001101001100100000100",
			1300 => "0000000001010010010101",
			1301 => "0000000001010010010101",
			1302 => "0011101100000000010000",
			1303 => "0000011101111100001100",
			1304 => "0001010110100000001000",
			1305 => "0011101100010000000100",
			1306 => "0000000001010010010101",
			1307 => "0000000001010010010101",
			1308 => "0000000001010010010101",
			1309 => "0000000001010010010101",
			1310 => "0000011101111100001100",
			1311 => "0010101000100100001000",
			1312 => "0011110111010100000100",
			1313 => "0000000001010010010101",
			1314 => "0000000001010010010101",
			1315 => "0000000001010010010101",
			1316 => "0000000001010010010101",
			1317 => "0011001010111100000100",
			1318 => "0000000001010011001001",
			1319 => "0011010010011100010100",
			1320 => "0010100011101000000100",
			1321 => "0000000001010011001001",
			1322 => "0001100100111100001100",
			1323 => "0001001101101100000100",
			1324 => "0000000001010011001001",
			1325 => "0010010101010000000100",
			1326 => "0000000001010011001001",
			1327 => "0000000001010011001001",
			1328 => "0000000001010011001001",
			1329 => "0000000001010011001001",
			1330 => "0011001010111000010000",
			1331 => "0011100110010000000100",
			1332 => "0000000001010100010101",
			1333 => "0010111000011000000100",
			1334 => "0000000001010100010101",
			1335 => "0011010101001000000100",
			1336 => "0000000001010100010101",
			1337 => "0000000001010100010101",
			1338 => "0011010010011100010100",
			1339 => "0011001011000000010000",
			1340 => "0001100100111100001100",
			1341 => "0000011011111100000100",
			1342 => "0000000001010100010101",
			1343 => "0011011001010000000100",
			1344 => "0000000001010100010101",
			1345 => "0000000001010100010101",
			1346 => "0000000001010100010101",
			1347 => "0000000001010100010101",
			1348 => "0000000001010100010101",
			1349 => "0000101010000100010000",
			1350 => "0011100110010000000100",
			1351 => "0000000001010101110001",
			1352 => "0001101001100100001000",
			1353 => "0011111010000100000100",
			1354 => "0000000001010101110001",
			1355 => "0000000001010101110001",
			1356 => "0000000001010101110001",
			1357 => "0011111000001100010000",
			1358 => "0001001011101100000100",
			1359 => "0000000001010101110001",
			1360 => "0010101000010100001000",
			1361 => "0001101101011000000100",
			1362 => "0000000001010101110001",
			1363 => "0000000001010101110001",
			1364 => "0000000001010101110001",
			1365 => "0001001000000100001100",
			1366 => "0011101100010000000100",
			1367 => "0000000001010101110001",
			1368 => "0011011110101000000100",
			1369 => "0000000001010101110001",
			1370 => "0000000001010101110001",
			1371 => "0000000001010101110001",
			1372 => "0011001010111000010000",
			1373 => "0010100111110100000100",
			1374 => "0000000001010111010101",
			1375 => "0000011101111100001000",
			1376 => "0001111001001000000100",
			1377 => "1111111001010111010101",
			1378 => "0000000001010111010101",
			1379 => "0000000001010111010101",
			1380 => "0001111001001000001100",
			1381 => "0000101100000000000100",
			1382 => "0000000001010111010101",
			1383 => "0010101001000100000100",
			1384 => "0000000001010111010101",
			1385 => "0000000001010111010101",
			1386 => "0011000100011000001100",
			1387 => "0011010101001000001000",
			1388 => "0000011110010100000100",
			1389 => "0000000001010111010101",
			1390 => "0000000001010111010101",
			1391 => "0000000001010111010101",
			1392 => "0010000110011100000100",
			1393 => "0000000001010111010101",
			1394 => "0001000101000000000100",
			1395 => "0000000001010111010101",
			1396 => "0000000001010111010101",
			1397 => "0011001010111000011000",
			1398 => "0011011100100100001100",
			1399 => "0010010101010000000100",
			1400 => "0000000001011001001001",
			1401 => "0011100110111100000100",
			1402 => "0000000001011001001001",
			1403 => "0000000001011001001001",
			1404 => "0010110100000100000100",
			1405 => "0000000001011001001001",
			1406 => "0001111000000000000100",
			1407 => "0000000001011001001001",
			1408 => "0000000001011001001001",
			1409 => "0001110110100100001100",
			1410 => "0010010100101100000100",
			1411 => "0000000001011001001001",
			1412 => "0011101011111000000100",
			1413 => "0000000001011001001001",
			1414 => "0000000001011001001001",
			1415 => "0010000101000100001100",
			1416 => "0010001010110000000100",
			1417 => "0000000001011001001001",
			1418 => "0011001000000000000100",
			1419 => "0000000001011001001001",
			1420 => "0000000001011001001001",
			1421 => "0011001010111000000100",
			1422 => "0000000001011001001001",
			1423 => "0010010000001000000100",
			1424 => "0000000001011001001001",
			1425 => "0000000001011001001001",
			1426 => "0011001010111000010000",
			1427 => "0010100111110100000100",
			1428 => "0000000001011010110101",
			1429 => "0000011101111100001000",
			1430 => "0001111001001000000100",
			1431 => "1111111001011010110101",
			1432 => "0000000001011010110101",
			1433 => "0000000001011010110101",
			1434 => "0001111001001000010000",
			1435 => "0000101100000000000100",
			1436 => "0000000001011010110101",
			1437 => "0010101001000100001000",
			1438 => "0000011110010100000100",
			1439 => "0000000001011010110101",
			1440 => "0000000001011010110101",
			1441 => "0000000001011010110101",
			1442 => "0011000100011000001100",
			1443 => "0011010101001000001000",
			1444 => "0000011110010100000100",
			1445 => "0000000001011010110101",
			1446 => "0000000001011010110101",
			1447 => "0000000001011010110101",
			1448 => "0010000110011100000100",
			1449 => "0000000001011010110101",
			1450 => "0001000101000000000100",
			1451 => "0000000001011010110101",
			1452 => "0000000001011010110101",
			1453 => "0000100110111100001100",
			1454 => "0001101001100100001000",
			1455 => "0001001100010000000100",
			1456 => "0000000001011100000001",
			1457 => "0000000001011100000001",
			1458 => "0000000001011100000001",
			1459 => "0001000001011100000100",
			1460 => "0000000001011100000001",
			1461 => "0001100100111100010100",
			1462 => "0011000100001000000100",
			1463 => "0000000001011100000001",
			1464 => "0010100011101000000100",
			1465 => "0000000001011100000001",
			1466 => "0000101111101000001000",
			1467 => "0000010001000100000100",
			1468 => "0000000001011100000001",
			1469 => "0000000001011100000001",
			1470 => "0000000001011100000001",
			1471 => "0000000001011100000001",
			1472 => "0011111000001100100000",
			1473 => "0001111110110000001100",
			1474 => "0000011011111100001000",
			1475 => "0011011110101100000100",
			1476 => "0000000001011101101101",
			1477 => "0000000001011101101101",
			1478 => "0000000001011101101101",
			1479 => "0001001111100100001100",
			1480 => "0000111110110100000100",
			1481 => "0000000001011101101101",
			1482 => "0011100110010000000100",
			1483 => "0000000001011101101101",
			1484 => "0000000001011101101101",
			1485 => "0000010001000100000100",
			1486 => "0000000001011101101101",
			1487 => "0000000001011101101101",
			1488 => "0011001011000000010100",
			1489 => "0000011101111100010000",
			1490 => "0011101100010000000100",
			1491 => "0000000001011101101101",
			1492 => "0011011110101000000100",
			1493 => "0000000001011101101101",
			1494 => "0010010000001000000100",
			1495 => "0000000001011101101101",
			1496 => "0000000001011101101101",
			1497 => "0000000001011101101101",
			1498 => "0000000001011101101101",
			1499 => "0010000001110000101000",
			1500 => "0001000011000000011000",
			1501 => "0011101100010000010000",
			1502 => "0010101010100100000100",
			1503 => "0000000001011111000001",
			1504 => "0011011110000100001000",
			1505 => "0000011011111100000100",
			1506 => "0000000001011111000001",
			1507 => "0000000001011111000001",
			1508 => "0000000001011111000001",
			1509 => "0010011010100000000100",
			1510 => "0000000001011111000001",
			1511 => "0000000001011111000001",
			1512 => "0011010111111100001100",
			1513 => "0000010001000100000100",
			1514 => "0000000001011111000001",
			1515 => "0011101011111000000100",
			1516 => "0000000001011111000001",
			1517 => "0000000001011111000001",
			1518 => "0000000001011111000001",
			1519 => "0000000001011111000001",
			1520 => "0011001010111100001100",
			1521 => "0000010111101000001000",
			1522 => "0010000001010000000100",
			1523 => "0000000001100000101101",
			1524 => "0000000001100000101101",
			1525 => "0000000001100000101101",
			1526 => "0011101110110100001100",
			1527 => "0010101010100000000100",
			1528 => "0000000001100000101101",
			1529 => "0010010101010000000100",
			1530 => "0000000001100000101101",
			1531 => "0000000001100000101101",
			1532 => "0001000011000000010000",
			1533 => "0010011010100000001100",
			1534 => "0011000111001000000100",
			1535 => "0000000001100000101101",
			1536 => "0000010001111000000100",
			1537 => "0000000001100000101101",
			1538 => "0000000001100000101101",
			1539 => "0000000001100000101101",
			1540 => "0000111111100100001100",
			1541 => "0000010111101000000100",
			1542 => "0000000001100000101101",
			1543 => "0011001010111000000100",
			1544 => "0000000001100000101101",
			1545 => "0000000001100000101101",
			1546 => "0000000001100000101101",
			1547 => "0010011001111100000100",
			1548 => "0000000001100001101001",
			1549 => "0001010001000000011000",
			1550 => "0000001001101000000100",
			1551 => "0000000001100001101001",
			1552 => "0001100100111100010000",
			1553 => "0011101011111000001100",
			1554 => "0001110011100000000100",
			1555 => "0000000001100001101001",
			1556 => "0001111000011000000100",
			1557 => "0000000001100001101001",
			1558 => "0000000001100001101001",
			1559 => "0000000001100001101001",
			1560 => "0000000001100001101001",
			1561 => "0000000001100001101001",
			1562 => "0011001010111000011000",
			1563 => "0000000111000100010000",
			1564 => "0011011100100100000100",
			1565 => "0000000001100011011101",
			1566 => "0001010010110100001000",
			1567 => "0001010010110100000100",
			1568 => "0000000001100011011101",
			1569 => "0000000001100011011101",
			1570 => "0000000001100011011101",
			1571 => "0000101000001100000100",
			1572 => "0000000001100011011101",
			1573 => "0000000001100011011101",
			1574 => "0011010010011100011100",
			1575 => "0010011001111100000100",
			1576 => "0000000001100011011101",
			1577 => "0000101010000100001100",
			1578 => "0011100110010000000100",
			1579 => "0000000001100011011101",
			1580 => "0000010001111000000100",
			1581 => "0000000001100011011101",
			1582 => "0000000001100011011101",
			1583 => "0011101011111000001000",
			1584 => "0000000110001000000100",
			1585 => "0000000001100011011101",
			1586 => "0000000001100011011101",
			1587 => "0000000001100011011101",
			1588 => "0011101111010100000100",
			1589 => "0000000001100011011101",
			1590 => "0000000001100011011101",
			1591 => "0010011001111100001100",
			1592 => "0001101001100100001000",
			1593 => "0001001100010000000100",
			1594 => "0000000001100101001001",
			1595 => "0000000001100101001001",
			1596 => "0000000001100101001001",
			1597 => "0011101100000000010000",
			1598 => "0001001111100100000100",
			1599 => "0000000001100101001001",
			1600 => "0010000110011100001000",
			1601 => "0010001010110000000100",
			1602 => "0000000001100101001001",
			1603 => "0000000001100101001001",
			1604 => "0000000001100101001001",
			1605 => "0001000011000000001000",
			1606 => "0011110111010100000100",
			1607 => "0000000001100101001001",
			1608 => "0000000001100101001001",
			1609 => "0010000001010100010000",
			1610 => "0001000010010100000100",
			1611 => "0000000001100101001001",
			1612 => "0011010111111100001000",
			1613 => "0011111000101000000100",
			1614 => "0000000001100101001001",
			1615 => "0000000001100101001001",
			1616 => "0000000001100101001001",
			1617 => "0000000001100101001001",
			1618 => "0011001010111000010000",
			1619 => "0010100111110100000100",
			1620 => "0000000001100111000101",
			1621 => "0010010000001000001000",
			1622 => "0001111001001000000100",
			1623 => "1111111001100111000101",
			1624 => "0000000001100111000101",
			1625 => "0000000001100111000101",
			1626 => "0001110110100100010100",
			1627 => "0011010101001000010000",
			1628 => "0000101100000000000100",
			1629 => "0000000001100111000101",
			1630 => "0010010100101100000100",
			1631 => "0000000001100111000101",
			1632 => "0011101011111000000100",
			1633 => "0000000001100111000101",
			1634 => "0000000001100111000101",
			1635 => "0000000001100111000101",
			1636 => "0001111000011000001100",
			1637 => "0011101100010000000100",
			1638 => "0000000001100111000101",
			1639 => "0001010111100000000100",
			1640 => "0000000001100111000101",
			1641 => "0000000001100111000101",
			1642 => "0001011110000100001100",
			1643 => "0011111100111000001000",
			1644 => "0000101010000100000100",
			1645 => "0000000001100111000101",
			1646 => "0000000001100111000101",
			1647 => "0000000001100111000101",
			1648 => "0000000001100111000101",
			1649 => "0010010101010000000100",
			1650 => "1111111001101000011001",
			1651 => "0011101111010100011000",
			1652 => "0011100110010000000100",
			1653 => "0000001001101000011001",
			1654 => "0001001111100100000100",
			1655 => "1111111001101000011001",
			1656 => "0010010111101100000100",
			1657 => "1111111001101000011001",
			1658 => "0001101111000000001000",
			1659 => "0010001010110000000100",
			1660 => "0000000001101000011001",
			1661 => "0000001001101000011001",
			1662 => "0000000001101000011001",
			1663 => "0011101011111000001100",
			1664 => "0010011010100000000100",
			1665 => "1111111001101000011001",
			1666 => "0001000010010100000100",
			1667 => "1111111001101000011001",
			1668 => "0000001001101000011001",
			1669 => "1111111001101000011001",
			1670 => "0000101011111000100100",
			1671 => "0010100111110100100000",
			1672 => "0010001010110000010100",
			1673 => "0010110111010000000100",
			1674 => "0000000001101010000101",
			1675 => "0001110001101000001100",
			1676 => "0000111110110100000100",
			1677 => "0000000001101010000101",
			1678 => "0011100010000000000100",
			1679 => "0000000001101010000101",
			1680 => "0000000001101010000101",
			1681 => "0000000001101010000101",
			1682 => "0011101111010100001000",
			1683 => "0000011011111100000100",
			1684 => "0000000001101010000101",
			1685 => "0000000001101010000101",
			1686 => "0000000001101010000101",
			1687 => "0000000001101010000101",
			1688 => "0011010111111100010000",
			1689 => "0010000001110000001100",
			1690 => "0001001011110000000100",
			1691 => "0000000001101010000101",
			1692 => "0011101011111000000100",
			1693 => "0000001001101010000101",
			1694 => "0000000001101010000101",
			1695 => "0000000001101010000101",
			1696 => "0000000001101010000101",
			1697 => "0010000001110000110100",
			1698 => "0011101110110100010100",
			1699 => "0000100010000100001000",
			1700 => "0000011011111100000100",
			1701 => "0000000001101011110001",
			1702 => "0000000001101011110001",
			1703 => "0000111100000000001000",
			1704 => "0000010001000100000100",
			1705 => "0000000001101011110001",
			1706 => "0000001001101011110001",
			1707 => "0000000001101011110001",
			1708 => "0000011101111100010000",
			1709 => "0010110111010000000100",
			1710 => "0000000001101011110001",
			1711 => "0001110001101000001000",
			1712 => "0001101011001100000100",
			1713 => "0000000001101011110001",
			1714 => "1111111001101011110001",
			1715 => "0000000001101011110001",
			1716 => "0010000101000100001100",
			1717 => "0001001101101100000100",
			1718 => "0000000001101011110001",
			1719 => "0010110101100100000100",
			1720 => "0000001001101011110001",
			1721 => "0000000001101011110001",
			1722 => "0000000001101011110001",
			1723 => "1111111001101011110001",
			1724 => "0000011011111100001000",
			1725 => "0010011001111100000100",
			1726 => "1111111001101101100101",
			1727 => "0000000001101101100101",
			1728 => "0011100110111100010000",
			1729 => "0001001111100100001000",
			1730 => "0011100110010000000100",
			1731 => "0000000001101101100101",
			1732 => "1111111001101101100101",
			1733 => "0011001011000000000100",
			1734 => "0000001001101101100101",
			1735 => "0000000001101101100101",
			1736 => "0010010000001000001000",
			1737 => "0001010000110100000100",
			1738 => "0000000001101101100101",
			1739 => "1111111001101101100101",
			1740 => "0010110101100100001100",
			1741 => "0011000100011000001000",
			1742 => "0001101000010000000100",
			1743 => "0000001001101101100101",
			1744 => "0000000001101101100101",
			1745 => "0000000001101101100101",
			1746 => "0000011101111100001100",
			1747 => "0001111000011000000100",
			1748 => "0000000001101101100101",
			1749 => "0010110010001000000100",
			1750 => "0000000001101101100101",
			1751 => "0000000001101101100101",
			1752 => "0000000001101101100101",
			1753 => "0010011001111100010100",
			1754 => "0000001010101100010000",
			1755 => "0010010101010000000100",
			1756 => "0000000001101111101001",
			1757 => "0010001010110000001000",
			1758 => "0000001001101000000100",
			1759 => "0000000001101111101001",
			1760 => "0000000001101111101001",
			1761 => "0000000001101111101001",
			1762 => "1111111001101111101001",
			1763 => "0000111011111000100100",
			1764 => "0001000010010100011100",
			1765 => "0011100110111100010100",
			1766 => "0011001011000000001100",
			1767 => "0010011010100000001000",
			1768 => "0001011101000100000100",
			1769 => "0000001001101111101001",
			1770 => "0000000001101111101001",
			1771 => "0000000001101111101001",
			1772 => "0010001010110000000100",
			1773 => "0000000001101111101001",
			1774 => "0000000001101111101001",
			1775 => "0011111000001100000100",
			1776 => "0000000001101111101001",
			1777 => "1111111001101111101001",
			1778 => "0001100100111100000100",
			1779 => "0000001001101111101001",
			1780 => "0000000001101111101001",
			1781 => "0001010110100000001000",
			1782 => "0010011010100100000100",
			1783 => "0000000001101111101001",
			1784 => "0000000001101111101001",
			1785 => "1111111001101111101001",
			1786 => "0000010001000100000100",
			1787 => "1111111001110001010101",
			1788 => "0011011111010000100000",
			1789 => "0011101011111000011100",
			1790 => "0000011101111100010100",
			1791 => "0011011110000100001100",
			1792 => "0010000110011000000100",
			1793 => "0000011001110001010101",
			1794 => "0010110101100100000100",
			1795 => "0000010001110001010101",
			1796 => "0000010001110001010101",
			1797 => "0001001101101100000100",
			1798 => "0000000001110001010101",
			1799 => "0000010001110001010101",
			1800 => "0010011010100000000100",
			1801 => "0000011001110001010101",
			1802 => "0000010001110001010101",
			1803 => "1111111001110001010101",
			1804 => "0011100111010100001000",
			1805 => "0000010001111000000100",
			1806 => "1111111001110001010101",
			1807 => "0000010001110001010101",
			1808 => "0011101011111000001000",
			1809 => "0011111011101100000100",
			1810 => "1111111001110001010101",
			1811 => "0000001001110001010101",
			1812 => "1111111001110001010101",
			1813 => "0000011011111100000100",
			1814 => "1111111001110010100001",
			1815 => "0000111111100100100000",
			1816 => "0011100110010000000100",
			1817 => "0000001001110010100001",
			1818 => "0001001011101100001000",
			1819 => "0000111100010000000100",
			1820 => "0000000001110010100001",
			1821 => "1111111001110010100001",
			1822 => "0010010111101100000100",
			1823 => "0000000001110010100001",
			1824 => "0011101000001100001000",
			1825 => "0001110001101000000100",
			1826 => "0000001001110010100001",
			1827 => "0000000001110010100001",
			1828 => "0001001110000000000100",
			1829 => "1111111001110010100001",
			1830 => "0000001001110010100001",
			1831 => "1111111001110010100001",
			1832 => "0010000001110000111000",
			1833 => "0001001000000100101000",
			1834 => "0011101100010000011000",
			1835 => "0001101010011000001000",
			1836 => "0000100010000100000100",
			1837 => "0000000001110100010101",
			1838 => "0000000001110100010101",
			1839 => "0010100111110100001100",
			1840 => "0010011010100000001000",
			1841 => "0010011001111100000100",
			1842 => "0000000001110100010101",
			1843 => "0000001001110100010101",
			1844 => "0000000001110100010101",
			1845 => "0000000001110100010101",
			1846 => "0010010000001000001100",
			1847 => "0001011110101000001000",
			1848 => "0011011100100100000100",
			1849 => "0000000001110100010101",
			1850 => "1111111001110100010101",
			1851 => "0000000001110100010101",
			1852 => "0000000001110100010101",
			1853 => "0001010001000000001100",
			1854 => "0010010101010000000100",
			1855 => "0000000001110100010101",
			1856 => "0011101111100100000100",
			1857 => "0000001001110100010101",
			1858 => "0000000001110100010101",
			1859 => "0000000001110100010101",
			1860 => "1111111001110100010101",
			1861 => "0010011001111100010100",
			1862 => "0000001010101100010000",
			1863 => "0000010001000100000100",
			1864 => "1111111001110111000001",
			1865 => "0000001111001000001000",
			1866 => "0000011011111100000100",
			1867 => "0000000001110111000001",
			1868 => "0000000001110111000001",
			1869 => "0000000001110111000001",
			1870 => "1111111001110111000001",
			1871 => "0001110001101000100100",
			1872 => "0000111011111000011000",
			1873 => "0011001011000000010000",
			1874 => "0000011101111100001000",
			1875 => "0011101000001100000100",
			1876 => "0000001001110111000001",
			1877 => "0000000001110111000001",
			1878 => "0000010100110100000100",
			1879 => "0000000001110111000001",
			1880 => "0000000001110111000001",
			1881 => "0011001000000000000100",
			1882 => "0000000001110111000001",
			1883 => "0000000001110111000001",
			1884 => "0000010100110100000100",
			1885 => "1111111001110111000001",
			1886 => "0001011110101000000100",
			1887 => "0000000001110111000001",
			1888 => "0000000001110111000001",
			1889 => "0010100111110100001100",
			1890 => "0000111000001100001000",
			1891 => "0000001001101000000100",
			1892 => "0000000001110111000001",
			1893 => "0000000001110111000001",
			1894 => "0000000001110111000001",
			1895 => "0001000101000000000100",
			1896 => "1111111001110111000001",
			1897 => "0000000111000000001000",
			1898 => "0010010010101100000100",
			1899 => "0000000001110111000001",
			1900 => "0000000001110111000001",
			1901 => "0011001010111000000100",
			1902 => "0000000001110111000001",
			1903 => "0000000001110111000001",
			1904 => "0010000001110000111000",
			1905 => "0011100110010000001100",
			1906 => "0001101010011000000100",
			1907 => "0000000001111000110101",
			1908 => "0000010001000100000100",
			1909 => "0000000001111000110101",
			1910 => "0000001001111000110101",
			1911 => "0011000100011000011100",
			1912 => "0001001100111000001100",
			1913 => "0010001010110000001000",
			1914 => "0001101011001100000100",
			1915 => "0000000001111000110101",
			1916 => "1111111001111000110101",
			1917 => "0000000001111000110101",
			1918 => "0011101010000100000100",
			1919 => "0000001001111000110101",
			1920 => "0000011101111100000100",
			1921 => "1111111001111000110101",
			1922 => "0001001011110000000100",
			1923 => "0000000001111000110101",
			1924 => "0000000001111000110101",
			1925 => "0001110110100100000100",
			1926 => "0000000001111000110101",
			1927 => "0001000110001100001000",
			1928 => "0001101011001100000100",
			1929 => "0000000001111000110101",
			1930 => "1111111001111000110101",
			1931 => "0000000001111000110101",
			1932 => "1111111001111000110101",
			1933 => "0000010001000100000100",
			1934 => "1111111001111011001001",
			1935 => "0001111001001000100000",
			1936 => "0001000010010100010100",
			1937 => "0000110111011000001000",
			1938 => "0000011101111100000100",
			1939 => "0000000001111011001001",
			1940 => "0000000001111011001001",
			1941 => "0011000100011000001000",
			1942 => "0011011100100100000100",
			1943 => "0000000001111011001001",
			1944 => "0000000001111011001001",
			1945 => "0000000001111011001001",
			1946 => "0011101011111000001000",
			1947 => "0011000000001100000100",
			1948 => "0000000001111011001001",
			1949 => "0000001001111011001001",
			1950 => "0000000001111011001001",
			1951 => "0011000100011000010000",
			1952 => "0010001100011100001000",
			1953 => "0000111100000000000100",
			1954 => "0000000001111011001001",
			1955 => "0000000001111011001001",
			1956 => "0010000001010100000100",
			1957 => "0000000001111011001001",
			1958 => "0000000001111011001001",
			1959 => "0011101100010000001100",
			1960 => "0011011110000100000100",
			1961 => "0000000001111011001001",
			1962 => "0010100011101000000100",
			1963 => "0000000001111011001001",
			1964 => "0000000001111011001001",
			1965 => "0001110110100100000100",
			1966 => "0000000001111011001001",
			1967 => "0010000110011100000100",
			1968 => "0000000001111011001001",
			1969 => "1111111001111011001001",
			1970 => "0000011011111100000100",
			1971 => "1111111001111100011101",
			1972 => "0000111111100100100100",
			1973 => "0011100110010000000100",
			1974 => "0000001001111100011101",
			1975 => "0001001011101100001100",
			1976 => "0000111100010000000100",
			1977 => "0000000001111100011101",
			1978 => "0000110110111100000100",
			1979 => "1111111001111100011101",
			1980 => "1111111001111100011101",
			1981 => "0010010111101100000100",
			1982 => "1111111001111100011101",
			1983 => "0011101000001100001000",
			1984 => "0001110001101000000100",
			1985 => "0000001001111100011101",
			1986 => "0000000001111100011101",
			1987 => "0001001110000000000100",
			1988 => "1111111001111100011101",
			1989 => "0000001001111100011101",
			1990 => "1111111001111100011101",
			1991 => "0000010001000100000100",
			1992 => "1111111001111110000001",
			1993 => "0011011001010000100100",
			1994 => "0010000001110000100000",
			1995 => "0000101101101100011100",
			1996 => "0011010101001000010000",
			1997 => "0011000100011000001000",
			1998 => "0001001101101100000100",
			1999 => "0000001001111110000001",
			2000 => "0000001001111110000001",
			2001 => "0000100111010100000100",
			2002 => "0000000001111110000001",
			2003 => "0000001001111110000001",
			2004 => "0000001111001000000100",
			2005 => "1111111001111110000001",
			2006 => "0001101111000000000100",
			2007 => "0000001001111110000001",
			2008 => "1111111001111110000001",
			2009 => "0000010001111110000001",
			2010 => "1111111001111110000001",
			2011 => "0000111011111000001000",
			2012 => "0000010001111000000100",
			2013 => "1111111001111110000001",
			2014 => "0000001001111110000001",
			2015 => "1111111001111110000001",
			2016 => "0000010001000100000100",
			2017 => "1111111001111111100101",
			2018 => "0011101011111000101100",
			2019 => "0000111100010000001000",
			2020 => "0000011011111100000100",
			2021 => "0000001001111111100101",
			2022 => "0000001001111111100101",
			2023 => "0001001011101100001100",
			2024 => "0011101110110100000100",
			2025 => "0000000001111111100101",
			2026 => "0001110110100100000100",
			2027 => "1111110001111111100101",
			2028 => "1111111001111111100101",
			2029 => "0010010111101100001000",
			2030 => "0001101011001100000100",
			2031 => "0000000001111111100101",
			2032 => "1111111001111111100101",
			2033 => "0001000011000000001000",
			2034 => "0010100111110100000100",
			2035 => "0000001001111111100101",
			2036 => "1111110001111111100101",
			2037 => "0000101101101100000100",
			2038 => "0000001001111111100101",
			2039 => "0000001001111111100101",
			2040 => "1111111001111111100101",
			2041 => "0000010001000100000100",
			2042 => "1111111010000000111001",
			2043 => "0011101011111000100100",
			2044 => "0010000001110000100000",
			2045 => "0011100110010000000100",
			2046 => "0000001010000000111001",
			2047 => "0000101111010100001100",
			2048 => "0000111100010000000100",
			2049 => "0000000010000000111001",
			2050 => "0010100010101100000100",
			2051 => "1111111010000000111001",
			2052 => "1111111010000000111001",
			2053 => "0010010111101100001000",
			2054 => "0011000100011000000100",
			2055 => "0000000010000000111001",
			2056 => "1111111010000000111001",
			2057 => "0010010111101100000100",
			2058 => "0000100010000000111001",
			2059 => "0000001010000000111001",
			2060 => "1111111010000000111001",
			2061 => "1111111010000000111001",
			2062 => "0010000001110000111000",
			2063 => "0001101010011000000100",
			2064 => "1111111010000010101101",
			2065 => "0011010111100000010100",
			2066 => "0001111110110000001100",
			2067 => "0000011011111100001000",
			2068 => "0000100110111100000100",
			2069 => "0000000010000010101101",
			2070 => "0000000010000010101101",
			2071 => "0000000010000010101101",
			2072 => "0001101111000000000100",
			2073 => "0000001010000010101101",
			2074 => "0000000010000010101101",
			2075 => "0001001000000100010100",
			2076 => "0011100111010100010000",
			2077 => "0000100111010100001000",
			2078 => "0011100010000100000100",
			2079 => "0000000010000010101101",
			2080 => "1111111010000010101101",
			2081 => "0011011111010000000100",
			2082 => "0000001010000010101101",
			2083 => "0000000010000010101101",
			2084 => "1111111010000010101101",
			2085 => "0001010001000000001000",
			2086 => "0011101111100100000100",
			2087 => "0000001010000010101101",
			2088 => "0000000010000010101101",
			2089 => "0000000010000010101101",
			2090 => "1111111010000010101101",
			2091 => "0010000001110000110100",
			2092 => "0001101010011000000100",
			2093 => "1111111010000100011001",
			2094 => "0011010111100000010100",
			2095 => "0000010001000100000100",
			2096 => "0000000010000100011001",
			2097 => "0001101111000000001100",
			2098 => "0011000100001000001000",
			2099 => "0011000100001000000100",
			2100 => "0000000010000100011001",
			2101 => "0000000010000100011001",
			2102 => "0000001010000100011001",
			2103 => "0000000010000100011001",
			2104 => "0011001010111000000100",
			2105 => "1111111010000100011001",
			2106 => "0010010111101100001100",
			2107 => "0011000100011000000100",
			2108 => "0000000010000100011001",
			2109 => "0000101111010100000100",
			2110 => "0000000010000100011001",
			2111 => "1111111010000100011001",
			2112 => "0011010111111100001000",
			2113 => "0001001110000000000100",
			2114 => "0000000010000100011001",
			2115 => "0000001010000100011001",
			2116 => "0000000010000100011001",
			2117 => "1111111010000100011001",
			2118 => "0000010001000100000100",
			2119 => "1111111010000110010101",
			2120 => "0011100110010000000100",
			2121 => "0000001010000110010101",
			2122 => "0011000100011000011100",
			2123 => "0001000110101100000100",
			2124 => "1111111010000110010101",
			2125 => "0011101100000000001000",
			2126 => "0000100110111100000100",
			2127 => "0000000010000110010101",
			2128 => "0000001010000110010101",
			2129 => "0001000010010100001000",
			2130 => "0011000100011000000100",
			2131 => "1111111010000110010101",
			2132 => "0000000010000110010101",
			2133 => "0011101011111000000100",
			2134 => "0000001010000110010101",
			2135 => "1111111010000110010101",
			2136 => "0001110110100100001000",
			2137 => "0000110000010000000100",
			2138 => "0000001010000110010101",
			2139 => "0000000010000110010101",
			2140 => "0011000100011000001000",
			2141 => "0000011101111100000100",
			2142 => "1111110010000110010101",
			2143 => "0000000010000110010101",
			2144 => "0011100111010100001000",
			2145 => "0010010111101100000100",
			2146 => "1111111010000110010101",
			2147 => "0000001010000110010101",
			2148 => "1111111010000110010101",
			2149 => "0000010001000100000100",
			2150 => "1111111010001000111011",
			2151 => "0011100110010000001000",
			2152 => "0001101010011000000100",
			2153 => "0000000010001000111011",
			2154 => "0000001010001000111011",
			2155 => "0011001010111000010100",
			2156 => "0011011100100100001100",
			2157 => "0000010111101000000100",
			2158 => "0000000010001000111011",
			2159 => "0001001110100100000100",
			2160 => "0000001010001000111011",
			2161 => "0000000010001000111011",
			2162 => "0000011101111100000100",
			2163 => "1111111010001000111011",
			2164 => "0000000010001000111011",
			2165 => "0001110001101000011100",
			2166 => "0010100011101000001100",
			2167 => "0000101100000000000100",
			2168 => "0000000010001000111011",
			2169 => "0011011110000100000100",
			2170 => "0000001010001000111011",
			2171 => "0000000010001000111011",
			2172 => "0001100100111100001000",
			2173 => "0001001100111000000100",
			2174 => "0000000010001000111011",
			2175 => "0000001010001000111011",
			2176 => "0011010101001000000100",
			2177 => "0000000010001000111011",
			2178 => "0000000010001000111011",
			2179 => "0011000100011000001100",
			2180 => "0010100011101000000100",
			2181 => "0000000010001000111011",
			2182 => "0001101000010000000100",
			2183 => "0000001010001000111011",
			2184 => "0000000010001000111011",
			2185 => "0010001100011100000100",
			2186 => "0000000010001000111011",
			2187 => "0001000101000000000100",
			2188 => "1111111010001000111011",
			2189 => "0000000010001000111011",
			2190 => "0000000010001000111101",
			2191 => "0000000010001001000001",
			2192 => "0000000010001001000101",
			2193 => "0000000010001001001001",
			2194 => "0000000010001001001101",
			2195 => "0000000010001001010001",
			2196 => "0000000010001001010101",
			2197 => "0000000010001001011001",
			2198 => "0000000010001001011101",
			2199 => "0000000010001001100001",
			2200 => "0000000010001001100101",
			2201 => "0000000010001001101001",
			2202 => "0000000010001001101101",
			2203 => "0000000010001001110001",
			2204 => "0000000010001001110101",
			2205 => "0000000010001001111001",
			2206 => "0000000010001001111101",
			2207 => "0000000010001010000001",
			2208 => "0000000010001010000101",
			2209 => "0000000010001010001001",
			2210 => "0000000010001010001101",
			2211 => "0000000010001010010001",
			2212 => "0000000010001010010101",
			2213 => "0000000010001010011001",
			2214 => "0000000010001010011101",
			2215 => "0000000010001010100001",
			2216 => "0000000010001010100101",
			2217 => "0011101100000000000100",
			2218 => "0000000010001010110001",
			2219 => "0000000010001010110001",
			2220 => "0010001100011100000100",
			2221 => "0000000010001010111101",
			2222 => "0000000010001010111101",
			2223 => "0010010000001000000100",
			2224 => "0000000010001011001001",
			2225 => "0000000010001011001001",
			2226 => "0011100110010000001000",
			2227 => "0011100101001000000100",
			2228 => "0000000010001011011101",
			2229 => "0000000010001011011101",
			2230 => "0000000010001011011101",
			2231 => "0000010111101000001000",
			2232 => "0010010111101100000100",
			2233 => "0000000010001011110001",
			2234 => "0000000010001011110001",
			2235 => "0000000010001011110001",
			2236 => "0000011011111100000100",
			2237 => "0000000010001100000101",
			2238 => "0010011010100100000100",
			2239 => "0000000010001100000101",
			2240 => "0000000010001100000101",
			2241 => "0011100110010000001100",
			2242 => "0011100101001000000100",
			2243 => "0000000010001100100001",
			2244 => "0000111100000000000100",
			2245 => "0000000010001100100001",
			2246 => "0000000010001100100001",
			2247 => "0000000010001100100001",
			2248 => "0000011101111100001100",
			2249 => "0011001011000000001000",
			2250 => "0010001010110000000100",
			2251 => "0000000010001100111101",
			2252 => "0000000010001100111101",
			2253 => "0000000010001100111101",
			2254 => "0000000010001100111101",
			2255 => "0011101100000000001100",
			2256 => "0011111100010000000100",
			2257 => "0000000010001101100001",
			2258 => "0011111000001100000100",
			2259 => "0000000010001101100001",
			2260 => "0000000010001101100001",
			2261 => "0011111000001100000100",
			2262 => "0000000010001101100001",
			2263 => "0000000010001101100001",
			2264 => "0011100110010000001100",
			2265 => "0010010101010000000100",
			2266 => "0000000010001110001101",
			2267 => "0000001100000100000100",
			2268 => "0000000010001110001101",
			2269 => "0000000010001110001101",
			2270 => "0000010100110100001000",
			2271 => "0011000100001000000100",
			2272 => "0000000010001110001101",
			2273 => "0000000010001110001101",
			2274 => "0000000010001110001101",
			2275 => "0000011110010100000100",
			2276 => "0000000010001110110001",
			2277 => "0010011010100100001100",
			2278 => "0010000001110000001000",
			2279 => "0010001010110000000100",
			2280 => "0000000010001110110001",
			2281 => "0000000010001110110001",
			2282 => "0000000010001110110001",
			2283 => "0000000010001110110001",
			2284 => "0010000001010100010000",
			2285 => "0011011111010000001100",
			2286 => "0010001000010100000100",
			2287 => "0000000010001111010101",
			2288 => "0011010101110100000100",
			2289 => "0000000010001111010101",
			2290 => "0000000010001111010101",
			2291 => "0000000010001111010101",
			2292 => "0000000010001111010101",
			2293 => "0010010000001000010000",
			2294 => "0011100110010000000100",
			2295 => "0000000010001111111001",
			2296 => "0000100011000000001000",
			2297 => "0000111100010000000100",
			2298 => "0000000010001111111001",
			2299 => "0000000010001111111001",
			2300 => "0000000010001111111001",
			2301 => "0000000010001111111001",
			2302 => "0011100110010000010000",
			2303 => "0011100101001000000100",
			2304 => "0000000010010000100101",
			2305 => "0000101110010000000100",
			2306 => "0000000010010000100101",
			2307 => "0000101100111000000100",
			2308 => "0000000010010000100101",
			2309 => "0000000010010000100101",
			2310 => "0001000011000000000100",
			2311 => "0000000010010000100101",
			2312 => "0000000010010000100101",
			2313 => "0010010111101100001000",
			2314 => "0010110100000100000100",
			2315 => "0000000010010001011001",
			2316 => "0000000010010001011001",
			2317 => "0001001101101100000100",
			2318 => "0000000010010001011001",
			2319 => "0011111100111000001100",
			2320 => "0011001000000000001000",
			2321 => "0010101000010100000100",
			2322 => "0000000010010001011001",
			2323 => "0000000010010001011001",
			2324 => "0000000010010001011001",
			2325 => "0000000010010001011001",
			2326 => "0011100110010000000100",
			2327 => "0000000010010010000101",
			2328 => "0010010000001000010000",
			2329 => "0011001011000000001100",
			2330 => "0011000100001000000100",
			2331 => "0000000010010010000101",
			2332 => "0000011101111100000100",
			2333 => "0000000010010010000101",
			2334 => "0000000010010010000101",
			2335 => "0000000010010010000101",
			2336 => "0000000010010010000101",
			2337 => "0000101000001100010100",
			2338 => "0011100110010000001000",
			2339 => "0000011011111100000100",
			2340 => "0000000010010011010001",
			2341 => "0000000010010011010001",
			2342 => "0001001101101100001000",
			2343 => "0011001000000000000100",
			2344 => "0000000010010011010001",
			2345 => "0000000010010011010001",
			2346 => "0000000010010011010001",
			2347 => "0011100111010100001100",
			2348 => "0000001111000100001000",
			2349 => "0000010001000100000100",
			2350 => "0000000010010011010001",
			2351 => "0000000010010011010001",
			2352 => "0000000010010011010001",
			2353 => "0000011101111100000100",
			2354 => "0000000010010011010001",
			2355 => "0000000010010011010001",
			2356 => "0000101010000100010000",
			2357 => "0011001000000000001100",
			2358 => "0001101001100100001000",
			2359 => "0011100010000000000100",
			2360 => "0000000010010100011101",
			2361 => "0000000010010100011101",
			2362 => "0000000010010100011101",
			2363 => "0000000010010100011101",
			2364 => "0011101100000000010000",
			2365 => "0001101101011000000100",
			2366 => "0000000010010100011101",
			2367 => "0011001011000000001000",
			2368 => "0010101000010100000100",
			2369 => "0000000010010100011101",
			2370 => "0000000010010100011101",
			2371 => "0000000010010100011101",
			2372 => "0001000010010100000100",
			2373 => "0000000010010100011101",
			2374 => "0000000010010100011101",
			2375 => "0000011110010100001100",
			2376 => "0010010100101100001000",
			2377 => "0001001100010000000100",
			2378 => "0000000010010101100001",
			2379 => "0000000010010101100001",
			2380 => "0000000010010101100001",
			2381 => "0011010111111100010100",
			2382 => "0001000001011100000100",
			2383 => "0000000010010101100001",
			2384 => "0011101011111000001100",
			2385 => "0001100100111100001000",
			2386 => "0000000110001000000100",
			2387 => "0000000010010101100001",
			2388 => "0000000010010101100001",
			2389 => "0000000010010101100001",
			2390 => "0000000010010101100001",
			2391 => "0000000010010101100001",
			2392 => "0011001010111100001100",
			2393 => "0010001010110000000100",
			2394 => "0000000010010110101101",
			2395 => "0000010111101000000100",
			2396 => "0000000010010110101101",
			2397 => "0000000010010110101101",
			2398 => "0001000011000000001000",
			2399 => "0010001100011100000100",
			2400 => "0000000010010110101101",
			2401 => "0000000010010110101101",
			2402 => "0001100100111100010000",
			2403 => "0010000001110000001100",
			2404 => "0000101111101000001000",
			2405 => "0011001001110100000100",
			2406 => "0000000010010110101101",
			2407 => "0000000010010110101101",
			2408 => "0000000010010110101101",
			2409 => "0000000010010110101101",
			2410 => "0000000010010110101101",
			2411 => "0011001010111000000100",
			2412 => "0000000010010111100001",
			2413 => "0011010010011100010100",
			2414 => "0011001011000000010000",
			2415 => "0011101011111000001100",
			2416 => "0000011011111100000100",
			2417 => "0000000010010111100001",
			2418 => "0011011001010000000100",
			2419 => "0000000010010111100001",
			2420 => "0000000010010111100001",
			2421 => "0000000010010111100001",
			2422 => "0000000010010111100001",
			2423 => "0000000010010111100001",
			2424 => "0000010111101000010000",
			2425 => "0011001010111100001100",
			2426 => "0001111000000000001000",
			2427 => "0001000110101100000100",
			2428 => "0000000010011000110101",
			2429 => "0000000010011000110101",
			2430 => "0000000010011000110101",
			2431 => "0000000010011000110101",
			2432 => "0001000001011100001000",
			2433 => "0000010001111000000100",
			2434 => "0000000010011000110101",
			2435 => "0000000010011000110101",
			2436 => "0011110011000000010000",
			2437 => "0001100100111100001100",
			2438 => "0000011100011000001000",
			2439 => "0011001000000000000100",
			2440 => "0000000010011000110101",
			2441 => "0000000010011000110101",
			2442 => "0000000010011000110101",
			2443 => "0000000010011000110101",
			2444 => "0000000010011000110101",
			2445 => "0000011011111100001000",
			2446 => "0000010001000100000100",
			2447 => "1100100010011010010001",
			2448 => "1100110010011010010001",
			2449 => "0000111111010100010100",
			2450 => "0010110101100100001100",
			2451 => "0010000110011000000100",
			2452 => "1110010010011010010001",
			2453 => "0000011101111100000100",
			2454 => "1111011010011010010001",
			2455 => "1110011010011010010001",
			2456 => "0000001011010100000100",
			2457 => "1100101010011010010001",
			2458 => "1110100010011010010001",
			2459 => "0011100111010100001000",
			2460 => "0001000011000000000100",
			2461 => "1100101010011010010001",
			2462 => "1111010010011010010001",
			2463 => "0011101011111000001000",
			2464 => "0000011101111100000100",
			2465 => "1100101010011010010001",
			2466 => "1101010010011010010001",
			2467 => "1100100010011010010001",
			2468 => "0000101011111000100000",
			2469 => "0010100111110100011000",
			2470 => "0011101100010000010000",
			2471 => "0010011010100000001100",
			2472 => "0000011110010100000100",
			2473 => "0000000010011011110101",
			2474 => "0001010110100000000100",
			2475 => "0000000010011011110101",
			2476 => "0000000010011011110101",
			2477 => "0000000010011011110101",
			2478 => "0000011101111100000100",
			2479 => "0000000010011011110101",
			2480 => "0000000010011011110101",
			2481 => "0000100000010000000100",
			2482 => "1111111010011011110101",
			2483 => "0000000010011011110101",
			2484 => "0000111011111000001100",
			2485 => "0001100100111100001000",
			2486 => "0000010001000100000100",
			2487 => "0000000010011011110101",
			2488 => "0000001010011011110101",
			2489 => "0000000010011011110101",
			2490 => "0000011101111100000100",
			2491 => "0000000010011011110101",
			2492 => "0000000010011011110101",
			2493 => "0011001010111000001100",
			2494 => "0010001100011100000100",
			2495 => "0000000010011101011001",
			2496 => "0010010000001000000100",
			2497 => "1111111010011101011001",
			2498 => "0000000010011101011001",
			2499 => "0001111001001000010000",
			2500 => "0001000110101100000100",
			2501 => "0000000010011101011001",
			2502 => "0011101111100100001000",
			2503 => "0000011011111100000100",
			2504 => "0000000010011101011001",
			2505 => "0000000010011101011001",
			2506 => "0000000010011101011001",
			2507 => "0011000100011000001100",
			2508 => "0011010101001000001000",
			2509 => "0000011110010100000100",
			2510 => "0000000010011101011001",
			2511 => "0000000010011101011001",
			2512 => "0000000010011101011001",
			2513 => "0010000110011100000100",
			2514 => "0000000010011101011001",
			2515 => "0001000101000000000100",
			2516 => "0000000010011101011001",
			2517 => "0000000010011101011001",
			2518 => "0011001010111100001100",
			2519 => "0000010111101000001000",
			2520 => "0000001001101000000100",
			2521 => "0000000010011110111101",
			2522 => "0000000010011110111101",
			2523 => "0000000010011110111101",
			2524 => "0001111001001000001100",
			2525 => "0001100100111100001000",
			2526 => "0000010001000100000100",
			2527 => "0000000010011110111101",
			2528 => "0000000010011110111101",
			2529 => "0000000010011110111101",
			2530 => "0010010000001000010000",
			2531 => "0011101110110100000100",
			2532 => "0000000010011110111101",
			2533 => "0001101011001100000100",
			2534 => "0000000010011110111101",
			2535 => "0000011101111100000100",
			2536 => "0000000010011110111101",
			2537 => "0000000010011110111101",
			2538 => "0011000100011000001000",
			2539 => "0011101011111000000100",
			2540 => "0000000010011110111101",
			2541 => "0000000010011110111101",
			2542 => "0000000010011110111101",
			2543 => "0000010111101000100000",
			2544 => "0010000110011100011000",
			2545 => "0010001001000100001000",
			2546 => "0010101010100100000100",
			2547 => "0000000010100000110001",
			2548 => "0000000010100000110001",
			2549 => "0011101100000000001100",
			2550 => "0010010101010000000100",
			2551 => "0000000010100000110001",
			2552 => "0001011101000100000100",
			2553 => "0000000010100000110001",
			2554 => "0000000010100000110001",
			2555 => "0000000010100000110001",
			2556 => "0000010111101000000100",
			2557 => "1111111010100000110001",
			2558 => "0000000010100000110001",
			2559 => "0011101000001100010100",
			2560 => "0010100011101000001100",
			2561 => "0000110111011000001000",
			2562 => "0000011101111100000100",
			2563 => "0000000010100000110001",
			2564 => "0000000010100000110001",
			2565 => "0000000010100000110001",
			2566 => "0000110000010000000100",
			2567 => "0000001010100000110001",
			2568 => "0000000010100000110001",
			2569 => "0001010110100000000100",
			2570 => "0000000010100000110001",
			2571 => "0000000010100000110001",
			2572 => "0011001010111100010000",
			2573 => "0000010111101000001100",
			2574 => "0010000001010000000100",
			2575 => "0000000010100010011101",
			2576 => "0001111000000000000100",
			2577 => "0000000010100010011101",
			2578 => "0000000010100010011101",
			2579 => "0000000010100010011101",
			2580 => "0001111001001000001100",
			2581 => "0010011010100000001000",
			2582 => "0000010001000100000100",
			2583 => "0000000010100010011101",
			2584 => "0000000010100010011101",
			2585 => "0000000010100010011101",
			2586 => "0011111000001100010000",
			2587 => "0010100010101100000100",
			2588 => "0000000010100010011101",
			2589 => "0010000110011100001000",
			2590 => "0000101100000000000100",
			2591 => "0000000010100010011101",
			2592 => "0000000010100010011101",
			2593 => "0000000010100010011101",
			2594 => "0000011101111100001000",
			2595 => "0011101100010000000100",
			2596 => "0000000010100010011101",
			2597 => "0000000010100010011101",
			2598 => "0000000010100010011101",
			2599 => "0011001010111000011100",
			2600 => "0000101000001100010000",
			2601 => "0010110101100100001100",
			2602 => "0011010101001000001000",
			2603 => "0001111001001000000100",
			2604 => "1111111010100100011001",
			2605 => "0000000010100100011001",
			2606 => "0000000010100100011001",
			2607 => "0000000010100100011001",
			2608 => "0011101010000100001000",
			2609 => "0011011011110100000100",
			2610 => "0000000010100100011001",
			2611 => "0000000010100100011001",
			2612 => "0000000010100100011001",
			2613 => "0011010101001000010100",
			2614 => "0011000100011000010000",
			2615 => "0000101100000000000100",
			2616 => "0000000010100100011001",
			2617 => "0011101011111000001000",
			2618 => "0001101101011000000100",
			2619 => "0000000010100100011001",
			2620 => "0000000010100100011001",
			2621 => "0000000010100100011001",
			2622 => "0000000010100100011001",
			2623 => "0001001011110000001100",
			2624 => "0011001010111000000100",
			2625 => "0000000010100100011001",
			2626 => "0010110100000100000100",
			2627 => "0000000010100100011001",
			2628 => "0000000010100100011001",
			2629 => "0000000010100100011001",
			2630 => "0010011001111100000100",
			2631 => "0000000010100101010101",
			2632 => "0001010001000000011000",
			2633 => "0000001001101000000100",
			2634 => "0000000010100101010101",
			2635 => "0001100100111100010000",
			2636 => "0011101011111000001100",
			2637 => "0001110011100000000100",
			2638 => "0000000010100101010101",
			2639 => "0010100011101000000100",
			2640 => "0000000010100101010101",
			2641 => "0000000010100101010101",
			2642 => "0000000010100101010101",
			2643 => "0000000010100101010101",
			2644 => "0000000010100101010101",
			2645 => "0000101100000000000100",
			2646 => "0000000010100110010001",
			2647 => "0010110101100100011000",
			2648 => "0010001010110000000100",
			2649 => "0000000010100110010001",
			2650 => "0001110001101000010000",
			2651 => "0001001011101100000100",
			2652 => "0000000010100110010001",
			2653 => "0010000001110000001000",
			2654 => "0011101011111000000100",
			2655 => "0000000010100110010001",
			2656 => "0000000010100110010001",
			2657 => "0000000010100110010001",
			2658 => "0000000010100110010001",
			2659 => "0000000010100110010001",
			2660 => "0010010101010000001100",
			2661 => "0010010101010000000100",
			2662 => "1111111010100111111101",
			2663 => "0010010101010000000100",
			2664 => "0000000010100111111101",
			2665 => "1111111010100111111101",
			2666 => "0011011111010000011000",
			2667 => "0011101011111000010100",
			2668 => "0011111001100000000100",
			2669 => "0000011010100111111101",
			2670 => "0000001001101000000100",
			2671 => "0000001010100111111101",
			2672 => "0011111011101100001000",
			2673 => "0010011010100000000100",
			2674 => "0000010010100111111101",
			2675 => "0000001010100111111101",
			2676 => "0000011010100111111101",
			2677 => "1111111010100111111101",
			2678 => "0011100111010100001000",
			2679 => "0010010000001000000100",
			2680 => "1111111010100111111101",
			2681 => "0000010010100111111101",
			2682 => "0011101011111000001000",
			2683 => "0011000100011000000100",
			2684 => "0000001010100111111101",
			2685 => "1111111010100111111101",
			2686 => "1111111010100111111101",
			2687 => "0010010101010000000100",
			2688 => "1111111010101001010001",
			2689 => "0011101111010100010100",
			2690 => "0011100110010000000100",
			2691 => "0000001010101001010001",
			2692 => "0001001111100100000100",
			2693 => "1111111010101001010001",
			2694 => "0010010111101100000100",
			2695 => "1111111010101001010001",
			2696 => "0001101111000000000100",
			2697 => "0000001010101001010001",
			2698 => "0000000010101001010001",
			2699 => "0011000100011000010000",
			2700 => "0001000010010100000100",
			2701 => "1111111010101001010001",
			2702 => "0011101011111000001000",
			2703 => "0000101100111000000100",
			2704 => "0000000010101001010001",
			2705 => "0000001010101001010001",
			2706 => "1111111010101001010001",
			2707 => "1111111010101001010001",
			2708 => "0011001010111000100000",
			2709 => "0000101000001100010000",
			2710 => "0010110101100100001100",
			2711 => "0011010101001000001000",
			2712 => "0001111001001000000100",
			2713 => "1111111010101011100101",
			2714 => "0000000010101011100101",
			2715 => "0000000010101011100101",
			2716 => "0000000010101011100101",
			2717 => "0011101010000100001100",
			2718 => "0010111001001000000100",
			2719 => "0000000010101011100101",
			2720 => "0000101100111000000100",
			2721 => "0000000010101011100101",
			2722 => "0000000010101011100101",
			2723 => "0000000010101011100101",
			2724 => "0010010111101100001100",
			2725 => "0011000100011000000100",
			2726 => "0000000010101011100101",
			2727 => "0011001000000000000100",
			2728 => "0000000010101011100101",
			2729 => "0000000010101011100101",
			2730 => "0011010101001000001100",
			2731 => "0000101100000000000100",
			2732 => "0000000010101011100101",
			2733 => "0011101011111000000100",
			2734 => "0000000010101011100101",
			2735 => "0000000010101011100101",
			2736 => "0001001011110000001100",
			2737 => "0000010001111000000100",
			2738 => "0000000010101011100101",
			2739 => "0001110110100100000100",
			2740 => "0000000010101011100101",
			2741 => "0000000010101011100101",
			2742 => "0011101111100100000100",
			2743 => "0000000010101011100101",
			2744 => "0000000010101011100101",
			2745 => "0000010001000100000100",
			2746 => "1111111010101100111001",
			2747 => "0011100110010000001000",
			2748 => "0010110000011100000100",
			2749 => "0000001010101100111001",
			2750 => "0000000010101100111001",
			2751 => "0001001100111000001100",
			2752 => "0001000110101100000100",
			2753 => "1111111010101100111001",
			2754 => "0000111100000000000100",
			2755 => "0000000010101100111001",
			2756 => "1111111010101100111001",
			2757 => "0011101011111000010000",
			2758 => "0000010111101000000100",
			2759 => "1111111010101100111001",
			2760 => "0001000010010100001000",
			2761 => "0011101111010100000100",
			2762 => "0000001010101100111001",
			2763 => "1111111010101100111001",
			2764 => "0000001010101100111001",
			2765 => "1111111010101100111001",
			2766 => "0000010001000100000100",
			2767 => "1111111010101110010101",
			2768 => "0011011111010000011000",
			2769 => "0010000001110000010100",
			2770 => "0000101101101100010000",
			2771 => "0011001011000000001100",
			2772 => "0000101100111000001000",
			2773 => "0000111000001100000100",
			2774 => "0000001010101110010101",
			2775 => "0000001010101110010101",
			2776 => "0000010010101110010101",
			2777 => "0000001010101110010101",
			2778 => "0000100010101110010101",
			2779 => "1111111010101110010101",
			2780 => "0001010110100000001000",
			2781 => "0000001000110000000100",
			2782 => "0000010010101110010101",
			2783 => "0000000010101110010101",
			2784 => "0011101111010100001000",
			2785 => "0000010111101000000100",
			2786 => "1111111010101110010101",
			2787 => "0000001010101110010101",
			2788 => "1111111010101110010101",
			2789 => "0010000001110000101100",
			2790 => "0001001000000100011100",
			2791 => "0011100111010100011000",
			2792 => "0000011011111100001000",
			2793 => "0010011001111100000100",
			2794 => "1111111010101111110001",
			2795 => "0000000010101111110001",
			2796 => "0001000001011100001100",
			2797 => "0001010010110100000100",
			2798 => "0000001010101111110001",
			2799 => "0011100110010000000100",
			2800 => "0000000010101111110001",
			2801 => "0000000010101111110001",
			2802 => "0000001010101111110001",
			2803 => "1111111010101111110001",
			2804 => "0001010001000000001100",
			2805 => "0000010001000100000100",
			2806 => "0000000010101111110001",
			2807 => "0011101111100100000100",
			2808 => "0000001010101111110001",
			2809 => "0000000010101111110001",
			2810 => "0000000010101111110001",
			2811 => "1111111010101111110001",
			2812 => "0010000001110000111000",
			2813 => "0011101110110100011000",
			2814 => "0000100010000100001100",
			2815 => "0000001011010100001000",
			2816 => "0000011011111100000100",
			2817 => "0000000010110001100101",
			2818 => "0000000010110001100101",
			2819 => "0000000010110001100101",
			2820 => "0000111100000000001000",
			2821 => "0000010001000100000100",
			2822 => "0000000010110001100101",
			2823 => "0000001010110001100101",
			2824 => "0000000010110001100101",
			2825 => "0000011101111100010000",
			2826 => "0011011100100100000100",
			2827 => "0000000010110001100101",
			2828 => "0001110001101000001000",
			2829 => "0001101011001100000100",
			2830 => "0000000010110001100101",
			2831 => "1111111010110001100101",
			2832 => "0000000010110001100101",
			2833 => "0011010101001000001000",
			2834 => "0000101000001100000100",
			2835 => "0000000010110001100101",
			2836 => "0000001010110001100101",
			2837 => "0011100111010100000100",
			2838 => "0000000010110001100101",
			2839 => "0000000010110001100101",
			2840 => "1111111010110001100101",
			2841 => "0000011011111100001000",
			2842 => "0010011001111100000100",
			2843 => "1111111010110011101001",
			2844 => "0000000010110011101001",
			2845 => "0011110000010000011100",
			2846 => "0001001111100100001100",
			2847 => "0000111110110100000100",
			2848 => "0000000010110011101001",
			2849 => "0011000100011000000100",
			2850 => "1111111010110011101001",
			2851 => "0000000010110011101001",
			2852 => "0011001011000000001000",
			2853 => "0000111010000100000100",
			2854 => "0000001010110011101001",
			2855 => "0000000010110011101001",
			2856 => "0010010111101100000100",
			2857 => "0000000010110011101001",
			2858 => "0000000010110011101001",
			2859 => "0010010000001000001000",
			2860 => "0010110111010000000100",
			2861 => "0000000010110011101001",
			2862 => "1111111010110011101001",
			2863 => "0011010101001000001000",
			2864 => "0000000111000000000100",
			2865 => "0000001010110011101001",
			2866 => "0000000010110011101001",
			2867 => "0010011010100000001000",
			2868 => "0010110110110100000100",
			2869 => "0000000010110011101001",
			2870 => "0000000010110011101001",
			2871 => "0010110000011100000100",
			2872 => "0000000010110011101001",
			2873 => "0000000010110011101001",
			2874 => "0010010101010000000100",
			2875 => "1111111010110101010101",
			2876 => "0011101111010100011000",
			2877 => "0011100110010000000100",
			2878 => "0000001010110101010101",
			2879 => "0001001111100100000100",
			2880 => "1111111010110101010101",
			2881 => "0010010111101100000100",
			2882 => "1111111010110101010101",
			2883 => "0001101111000000001000",
			2884 => "0010010111101100000100",
			2885 => "0000000010110101010101",
			2886 => "0000001010110101010101",
			2887 => "0000000010110101010101",
			2888 => "0011000100011000010000",
			2889 => "0001000010010100000100",
			2890 => "1111111010110101010101",
			2891 => "0011101011111000001000",
			2892 => "0000101100111000000100",
			2893 => "0000000010110101010101",
			2894 => "0000001010110101010101",
			2895 => "1111111010110101010101",
			2896 => "0011111111100100001000",
			2897 => "0001101001100100000100",
			2898 => "0000000010110101010101",
			2899 => "0000000010110101010101",
			2900 => "1111111010110101010101",
			2901 => "0010000001110000110000",
			2902 => "0001001000000100100000",
			2903 => "0011101010000100011100",
			2904 => "0000100111010100010100",
			2905 => "0011100010000100010000",
			2906 => "0001101010011000001000",
			2907 => "0000100010000100000100",
			2908 => "0000000010110110111001",
			2909 => "0000000010110110111001",
			2910 => "0001111110110000000100",
			2911 => "0000000010110110111001",
			2912 => "0000000010110110111001",
			2913 => "1111111010110110111001",
			2914 => "0001011101000100000100",
			2915 => "0000001010110110111001",
			2916 => "0000000010110110111001",
			2917 => "1111111010110110111001",
			2918 => "0011010111111100001100",
			2919 => "0001101101011000000100",
			2920 => "0000000010110110111001",
			2921 => "0011101111100100000100",
			2922 => "0000001010110110111001",
			2923 => "0000000010110110111001",
			2924 => "0000000010110110111001",
			2925 => "1111111010110110111001",
			2926 => "0010000001110000111000",
			2927 => "0001001000000100101000",
			2928 => "0010000110011100011100",
			2929 => "0011011100100100001000",
			2930 => "0010010101010000000100",
			2931 => "0000000010111000101101",
			2932 => "0000000010111000101101",
			2933 => "0001001111100100001000",
			2934 => "0011100010000000000100",
			2935 => "0000000010111000101101",
			2936 => "0000000010111000101101",
			2937 => "0000111111010100000100",
			2938 => "0000000010111000101101",
			2939 => "0010100111110100000100",
			2940 => "0000000010111000101101",
			2941 => "0000000010111000101101",
			2942 => "0010010000001000001000",
			2943 => "0001011110101000000100",
			2944 => "1111111010111000101101",
			2945 => "0000000010111000101101",
			2946 => "0000000010111000101101",
			2947 => "0001010001000000001100",
			2948 => "0010010101010000000100",
			2949 => "0000000010111000101101",
			2950 => "0011101111100100000100",
			2951 => "0000001010111000101101",
			2952 => "0000000010111000101101",
			2953 => "0000000010111000101101",
			2954 => "1111111010111000101101",
			2955 => "0010010101010000000100",
			2956 => "1111111010111010000001",
			2957 => "0011101011111000100100",
			2958 => "0011011001010000011100",
			2959 => "0000101101101100011000",
			2960 => "0011011111010000010000",
			2961 => "0000111100010000001000",
			2962 => "0010000110011000000100",
			2963 => "0000010010111010000001",
			2964 => "0000001010111010000001",
			2965 => "0001001011101100000100",
			2966 => "1111111010111010000001",
			2967 => "0000001010111010000001",
			2968 => "0000010001111000000100",
			2969 => "1111111010111010000001",
			2970 => "0000001010111010000001",
			2971 => "0000010010111010000001",
			2972 => "0011111011101100000100",
			2973 => "1111111010111010000001",
			2974 => "0000001010111010000001",
			2975 => "1111111010111010000001",
			2976 => "0000010001000100000100",
			2977 => "1111111010111011111101",
			2978 => "0001000010010100101100",
			2979 => "0011110000010000100000",
			2980 => "0001001111100100001100",
			2981 => "0000111110110100000100",
			2982 => "0000000010111011111101",
			2983 => "0001110001101000000100",
			2984 => "0000000010111011111101",
			2985 => "0000000010111011111101",
			2986 => "0011001011000000001000",
			2987 => "0000111000001100000100",
			2988 => "0000001010111011111101",
			2989 => "0000000010111011111101",
			2990 => "0000001111001000001000",
			2991 => "0000111010000100000100",
			2992 => "0000000010111011111101",
			2993 => "0000000010111011111101",
			2994 => "0000000010111011111101",
			2995 => "0001000010010100001000",
			2996 => "0010011010100100000100",
			2997 => "1111111010111011111101",
			2998 => "0000000010111011111101",
			2999 => "0000000010111011111101",
			3000 => "0000111111100100001000",
			3001 => "0001101000010000000100",
			3002 => "0000001010111011111101",
			3003 => "0000000010111011111101",
			3004 => "0010000101000100000100",
			3005 => "0000000010111011111101",
			3006 => "0000000010111011111101",
			3007 => "0000011011111100001000",
			3008 => "0010011001111100000100",
			3009 => "1111111010111110001001",
			3010 => "0000000010111110001001",
			3011 => "0001111001001000010000",
			3012 => "0000111011111000001100",
			3013 => "0010011010100000001000",
			3014 => "0011001101111000000100",
			3015 => "0000000010111110001001",
			3016 => "0000001010111110001001",
			3017 => "0000000010111110001001",
			3018 => "0000000010111110001001",
			3019 => "0000010001111000010000",
			3020 => "0011100110010000000100",
			3021 => "0000000010111110001001",
			3022 => "0010010111101100001000",
			3023 => "0001111000011000000100",
			3024 => "1111111010111110001001",
			3025 => "0000000010111110001001",
			3026 => "0000000010111110001001",
			3027 => "0011010101001000001100",
			3028 => "0000101111010100000100",
			3029 => "0000000010111110001001",
			3030 => "0011101011111000000100",
			3031 => "0000001010111110001001",
			3032 => "0000000010111110001001",
			3033 => "0011000100011000001100",
			3034 => "0010010000001000000100",
			3035 => "0000000010111110001001",
			3036 => "0001100100111100000100",
			3037 => "0000000010111110001001",
			3038 => "0000000010111110001001",
			3039 => "0010010000001000000100",
			3040 => "0000000010111110001001",
			3041 => "0000000010111110001001",
			3042 => "0010000001110000111100",
			3043 => "0001000010010100101000",
			3044 => "0011100110111100100000",
			3045 => "0001001100111000010100",
			3046 => "0011100110010000001100",
			3047 => "0001101010011000000100",
			3048 => "0000000011000000000101",
			3049 => "0011010000110100000100",
			3050 => "0000000011000000000101",
			3051 => "0000000011000000000101",
			3052 => "0011111010000100000100",
			3053 => "1111111011000000000101",
			3054 => "0000000011000000000101",
			3055 => "0000011110010100000100",
			3056 => "0000000011000000000101",
			3057 => "0010001010110000000100",
			3058 => "0000000011000000000101",
			3059 => "0000001011000000000101",
			3060 => "0000011101111100000100",
			3061 => "1111111011000000000101",
			3062 => "0000000011000000000101",
			3063 => "0011010111111100010000",
			3064 => "0000010001000100000100",
			3065 => "0000000011000000000101",
			3066 => "0001100100111100001000",
			3067 => "0011101011111000000100",
			3068 => "0000001011000000000101",
			3069 => "0000000011000000000101",
			3070 => "0000000011000000000101",
			3071 => "0000000011000000000101",
			3072 => "1111111011000000000101",
			3073 => "0000010001000100000100",
			3074 => "1111111011000010010001",
			3075 => "0001111001001000011000",
			3076 => "0001001101101100001100",
			3077 => "0000111100010000000100",
			3078 => "0000001011000010010001",
			3079 => "0001001011101100000100",
			3080 => "1111111011000010010001",
			3081 => "0000000011000010010001",
			3082 => "0011101011111000001000",
			3083 => "0001000010110000000100",
			3084 => "0000001011000010010001",
			3085 => "0000010011000010010001",
			3086 => "0000000011000010010001",
			3087 => "0011100110111100010100",
			3088 => "0010100011101000001000",
			3089 => "0000111100010000000100",
			3090 => "0000000011000010010001",
			3091 => "1111111011000010010001",
			3092 => "0010010100101100000100",
			3093 => "0000000011000010010001",
			3094 => "0000000110001000000100",
			3095 => "0000000011000010010001",
			3096 => "0000001011000010010001",
			3097 => "0000110111010100000100",
			3098 => "1111111011000010010001",
			3099 => "0001011100100100010000",
			3100 => "0001110110100100001000",
			3101 => "0000111111100100000100",
			3102 => "0000000011000010010001",
			3103 => "0000000011000010010001",
			3104 => "0001110001101000000100",
			3105 => "0000000011000010010001",
			3106 => "0000000011000010010001",
			3107 => "1111111011000010010001",
			3108 => "0000010001000100000100",
			3109 => "1111111011000011101101",
			3110 => "0011101011111000101000",
			3111 => "0000111100010000000100",
			3112 => "0000001011000011101101",
			3113 => "0001001011101100001100",
			3114 => "0011110110111100001000",
			3115 => "0011101110110100000100",
			3116 => "0000000011000011101101",
			3117 => "1111111011000011101101",
			3118 => "1111111011000011101101",
			3119 => "0000010111101000001000",
			3120 => "0011101111010100000100",
			3121 => "0000000011000011101101",
			3122 => "1111111011000011101101",
			3123 => "0001000011000000001000",
			3124 => "0010100111110100000100",
			3125 => "0000000011000011101101",
			3126 => "1111110011000011101101",
			3127 => "0000101101101100000100",
			3128 => "0000001011000011101101",
			3129 => "0000001011000011101101",
			3130 => "1111111011000011101101",
			3131 => "0010010101010000000100",
			3132 => "1111111011000101011001",
			3133 => "0011101011111000110000",
			3134 => "0011001011000000011100",
			3135 => "0000101101101100011000",
			3136 => "0011011111010000010000",
			3137 => "0011100110111100001000",
			3138 => "0001001011101100000100",
			3139 => "0000001011000101011001",
			3140 => "0000001011000101011001",
			3141 => "0001000011000000000100",
			3142 => "1111111011000101011001",
			3143 => "0000001011000101011001",
			3144 => "0001000011000000000100",
			3145 => "1111111011000101011001",
			3146 => "0000000011000101011001",
			3147 => "0000010011000101011001",
			3148 => "0011001000000000001000",
			3149 => "0010010111101100000100",
			3150 => "1111110011000101011001",
			3151 => "0000000011000101011001",
			3152 => "0011011001010000000100",
			3153 => "0000001011000101011001",
			3154 => "0000010001111000000100",
			3155 => "1111111011000101011001",
			3156 => "0000000011000101011001",
			3157 => "1111111011000101011001",
			3158 => "0000010001000100000100",
			3159 => "1111111011000111110101",
			3160 => "0001111001001000011100",
			3161 => "0001000011001100010100",
			3162 => "0000111100010000000100",
			3163 => "0000001011000111110101",
			3164 => "0001001011101100000100",
			3165 => "1111111011000111110101",
			3166 => "0011101011111000001000",
			3167 => "0001001101101100000100",
			3168 => "0000000011000111110101",
			3169 => "0000001011000111110101",
			3170 => "0000000011000111110101",
			3171 => "0011111110000000000100",
			3172 => "0000010011000111110101",
			3173 => "0000000011000111110101",
			3174 => "0011100110111100010000",
			3175 => "0010100011101000001000",
			3176 => "0000111100010000000100",
			3177 => "0000000011000111110101",
			3178 => "1111111011000111110101",
			3179 => "0000010111101000000100",
			3180 => "0000000011000111110101",
			3181 => "0000001011000111110101",
			3182 => "0011000100011000010000",
			3183 => "0001110110100100001000",
			3184 => "0000111111100100000100",
			3185 => "0000000011000111110101",
			3186 => "0000000011000111110101",
			3187 => "0011000100011000000100",
			3188 => "1111111011000111110101",
			3189 => "0000000011000111110101",
			3190 => "0010110000011100000100",
			3191 => "1111111011000111110101",
			3192 => "0000111000001100001000",
			3193 => "0001011100100100000100",
			3194 => "0000000011000111110101",
			3195 => "0000000011000111110101",
			3196 => "1111111011000111110101",
			3197 => "0010000001110000111100",
			3198 => "0001101010011000000100",
			3199 => "1111111011001001110001",
			3200 => "0011101100010000011000",
			3201 => "0011100110010000001000",
			3202 => "0011100101001000000100",
			3203 => "0000000011001001110001",
			3204 => "0000001011001001110001",
			3205 => "0000101010000100001100",
			3206 => "0000111100010000001000",
			3207 => "0010100011101000000100",
			3208 => "0000001011001001110001",
			3209 => "0000000011001001110001",
			3210 => "1111111011001001110001",
			3211 => "0000001011001001110001",
			3212 => "0001000011000000010000",
			3213 => "0010100111110100001100",
			3214 => "0010100011101000000100",
			3215 => "1111111011001001110001",
			3216 => "0010001100011100000100",
			3217 => "0000000011001001110001",
			3218 => "0000000011001001110001",
			3219 => "1111111011001001110001",
			3220 => "0011101011111000001100",
			3221 => "0001000010010100001000",
			3222 => "0000110111010100000100",
			3223 => "0000001011001001110001",
			3224 => "1111111011001001110001",
			3225 => "0000001011001001110001",
			3226 => "1111111011001001110001",
			3227 => "1111111011001001110001",
			3228 => "0000010001000100000100",
			3229 => "1111111011001011111101",
			3230 => "0011100110010000001000",
			3231 => "0011111000001100000100",
			3232 => "0000000011001011111101",
			3233 => "0000000011001011111101",
			3234 => "0000010111101000001100",
			3235 => "0011011101000100000100",
			3236 => "0000000011001011111101",
			3237 => "0010010111101100000100",
			3238 => "1111111011001011111101",
			3239 => "0000000011001011111101",
			3240 => "0001110110100100011000",
			3241 => "0011001010111000001100",
			3242 => "0000110111011000000100",
			3243 => "0000000011001011111101",
			3244 => "0011011100100100000100",
			3245 => "0000000011001011111101",
			3246 => "0000000011001011111101",
			3247 => "0001100100111100001000",
			3248 => "0000111011111000000100",
			3249 => "0000001011001011111101",
			3250 => "0000000011001011111101",
			3251 => "0000000011001011111101",
			3252 => "0001110001101000001100",
			3253 => "0011001010111000000100",
			3254 => "0000000011001011111101",
			3255 => "0010110110110100000100",
			3256 => "0000000011001011111101",
			3257 => "0000000011001011111101",
			3258 => "0011111100111000001000",
			3259 => "0001111000011000000100",
			3260 => "0000000011001011111101",
			3261 => "0000000011001011111101",
			3262 => "0000000011001011111101",
			3263 => "0000010001000100000100",
			3264 => "1111111011001110110011",
			3265 => "0011100110010000001000",
			3266 => "0010110000011100000100",
			3267 => "0000001011001110110011",
			3268 => "0000000011001110110011",
			3269 => "0011001010111000011100",
			3270 => "0001010010110100001100",
			3271 => "0000010111101000000100",
			3272 => "0000000011001110110011",
			3273 => "0010001100000100000100",
			3274 => "0000000011001110110011",
			3275 => "0000000011001110110011",
			3276 => "0000010001111000001000",
			3277 => "0011010101001000000100",
			3278 => "1111111011001110110011",
			3279 => "0000000011001110110011",
			3280 => "0010010000001000000100",
			3281 => "0000000011001110110011",
			3282 => "0000000011001110110011",
			3283 => "0001110001101000100000",
			3284 => "0010100011101000010000",
			3285 => "0011011110000100001000",
			3286 => "0001111001001000000100",
			3287 => "0000000011001110110011",
			3288 => "0000000011001110110011",
			3289 => "0010110101100100000100",
			3290 => "0000000011001110110011",
			3291 => "0000000011001110110011",
			3292 => "0011001011000000001000",
			3293 => "0011101000001100000100",
			3294 => "0000001011001110110011",
			3295 => "0000000011001110110011",
			3296 => "0011001000000000000100",
			3297 => "0000000011001110110011",
			3298 => "0000000011001110110011",
			3299 => "0011000100011000001100",
			3300 => "0010100011101000000100",
			3301 => "0000000011001110110011",
			3302 => "0010000001010100000100",
			3303 => "0000000011001110110011",
			3304 => "0000000011001110110011",
			3305 => "0010001100011100000100",
			3306 => "0000000011001110110011",
			3307 => "1111111011001110110011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1096, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2190, initial_addr_3'length));
	end generate gen_rom_11;

	gen_rom_12: if SELECT_ROM = 12 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0000000000000001010001",
			20 => "0000000000000001010101",
			21 => "0000000000000001011001",
			22 => "0000000000000001011101",
			23 => "0000000000000001100001",
			24 => "0000000000000001100101",
			25 => "0000000000000001101001",
			26 => "0000000000000001101101",
			27 => "0000000000000001110001",
			28 => "0000000000000001110101",
			29 => "0001000001001100000100",
			30 => "0000000000000010000001",
			31 => "0000000000000010000001",
			32 => "0001000011011000000100",
			33 => "0000000000000010001101",
			34 => "0000000000000010001101",
			35 => "0001000100111000000100",
			36 => "0000000000000010011001",
			37 => "0000000000000010011001",
			38 => "0001000011111000000100",
			39 => "0000000000000010100101",
			40 => "0000000000000010100101",
			41 => "0001000100111000000100",
			42 => "0000000000000010110001",
			43 => "0000000000000010110001",
			44 => "0000011111001100000100",
			45 => "0000000000000010111101",
			46 => "0000000000000010111101",
			47 => "0001000011111000000100",
			48 => "0000000000000011001001",
			49 => "0000000000000011001001",
			50 => "0001000000010100000100",
			51 => "0000000000000011011101",
			52 => "0001001010010000000100",
			53 => "0000000000000011011101",
			54 => "0000000000000011011101",
			55 => "0001000101100000001000",
			56 => "0010011010011000000100",
			57 => "0000000000000011110001",
			58 => "0000000000000011110001",
			59 => "0000000000000011110001",
			60 => "0000100110101100000100",
			61 => "0000000000000100000101",
			62 => "0000101101101100000100",
			63 => "0000000000000100000101",
			64 => "0000000000000100000101",
			65 => "0000101011111000000100",
			66 => "0000000000000100011001",
			67 => "0000101101101100000100",
			68 => "0000000000000100011001",
			69 => "0000000000000100011001",
			70 => "0000100110101100000100",
			71 => "0000000000000100101101",
			72 => "0000101111101000000100",
			73 => "0000000000000100101101",
			74 => "0000000000000100101101",
			75 => "0001000100111000001000",
			76 => "0010011010011000000100",
			77 => "0000000000000101000001",
			78 => "0000000000000101000001",
			79 => "0000000000000101000001",
			80 => "0000011101011100001000",
			81 => "0000101011101100000100",
			82 => "0000000000000101010101",
			83 => "0000000000000101010101",
			84 => "0000000000000101010101",
			85 => "0000101011111000001100",
			86 => "0001101001100100001000",
			87 => "0000010000111100000100",
			88 => "0000000000000101110001",
			89 => "0000000000000101110001",
			90 => "0000000000000101110001",
			91 => "0000000000000101110001",
			92 => "0011100111110000001100",
			93 => "0001001001000000000100",
			94 => "0000000000000110001101",
			95 => "0001001010010000000100",
			96 => "0000000000000110001101",
			97 => "0000000000000110001101",
			98 => "0000000000000110001101",
			99 => "0001000010100100000100",
			100 => "0000000000000110101001",
			101 => "0000100000010000000100",
			102 => "0000000000000110101001",
			103 => "0000101111101000000100",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0000011101011100001100",
			107 => "0000101011101100001000",
			108 => "0010011101011000000100",
			109 => "0000000000000111000101",
			110 => "0000000000000111000101",
			111 => "0000000000000111000101",
			112 => "0000000000000111000101",
			113 => "0000011101011100001000",
			114 => "0000101011101100000100",
			115 => "0000000000000111101001",
			116 => "0000000000000111101001",
			117 => "0001010111110000001000",
			118 => "0001001110111000000100",
			119 => "0000000000000111101001",
			120 => "0000000000000111101001",
			121 => "0000000000000111101001",
			122 => "0000011101101000000100",
			123 => "0000000000001000001101",
			124 => "0011101110101100001100",
			125 => "0001101011001100001000",
			126 => "0001110111001000000100",
			127 => "0000000000001000001101",
			128 => "0000000000001000001101",
			129 => "0000000000001000001101",
			130 => "0000000000001000001101",
			131 => "0001000011010100000100",
			132 => "0000000000001000110001",
			133 => "0000100110101100000100",
			134 => "0000000000001000110001",
			135 => "0000100011000000001000",
			136 => "0001001010010000000100",
			137 => "0000000000001000110001",
			138 => "0000000000001000110001",
			139 => "0000000000001000110001",
			140 => "0001000011011000000100",
			141 => "0000000000001001010101",
			142 => "0011010100010000001100",
			143 => "0011100110000100000100",
			144 => "0000000000001001010101",
			145 => "0011011000011000000100",
			146 => "0000000000001001010101",
			147 => "0000000000001001010101",
			148 => "0000000000001001010101",
			149 => "0000011011101000001000",
			150 => "0001000011111000000100",
			151 => "0000000000001010000001",
			152 => "0000000000001010000001",
			153 => "0011101001010100001100",
			154 => "0001111101111000000100",
			155 => "0000000000001010000001",
			156 => "0000011111001100000100",
			157 => "0000000000001010000001",
			158 => "0000000000001010000001",
			159 => "0000000000001010000001",
			160 => "0000011111001100001000",
			161 => "0001000100111000000100",
			162 => "0000000000001010101101",
			163 => "0000000000001010101101",
			164 => "0011100111110000001100",
			165 => "0001111101111000000100",
			166 => "0000000000001010101101",
			167 => "0001101001100100000100",
			168 => "0000000000001010101101",
			169 => "0000000000001010101101",
			170 => "0000000000001010101101",
			171 => "0000100110101100001100",
			172 => "0000000011111100000100",
			173 => "0000000000001011100001",
			174 => "0011001110001100000100",
			175 => "0000000000001011100001",
			176 => "0000000000001011100001",
			177 => "0011111100010000001100",
			178 => "0010100001110000001000",
			179 => "0011000011011100000100",
			180 => "0000000000001011100001",
			181 => "0000000000001011100001",
			182 => "0000000000001011100001",
			183 => "0000000000001011100001",
			184 => "0001000011110100000100",
			185 => "0000000000001100010101",
			186 => "0010110011100000001100",
			187 => "0000011111001100000100",
			188 => "0000000000001100010101",
			189 => "0001111101111000000100",
			190 => "0000000000001100010101",
			191 => "0000000000001100010101",
			192 => "0010001011010100000100",
			193 => "0000000000001100010101",
			194 => "0011100111110000000100",
			195 => "0000000000001100010101",
			196 => "0000000000001100010101",
			197 => "0010010001111000001000",
			198 => "0000101011101100000100",
			199 => "0000000000001101001001",
			200 => "0000000000001101001001",
			201 => "0011101001010100010000",
			202 => "0011001100110000000100",
			203 => "0000000000001101001001",
			204 => "0000100111011000000100",
			205 => "0000000000001101001001",
			206 => "0001101111000000000100",
			207 => "0000000000001101001001",
			208 => "0000000000001101001001",
			209 => "0000000000001101001001",
			210 => "0010011011111100000100",
			211 => "0000000000001101110101",
			212 => "0011101110101100010000",
			213 => "0001101011001100001100",
			214 => "0010110001111100000100",
			215 => "0000000000001101110101",
			216 => "0011110001000000000100",
			217 => "0000000000001101110101",
			218 => "0000000000001101110101",
			219 => "0000000000001101110101",
			220 => "0000000000001101110101",
			221 => "0000101000001100001100",
			222 => "0001111100101000001000",
			223 => "0011001110001100000100",
			224 => "1111111000001110111001",
			225 => "0000000000001110111001",
			226 => "0000000000001110111001",
			227 => "0011110010000000010000",
			228 => "0010001010101100001100",
			229 => "0011100111110000001000",
			230 => "0000011011101000000100",
			231 => "0000000000001110111001",
			232 => "0000000000001110111001",
			233 => "0000000000001110111001",
			234 => "0000000000001110111001",
			235 => "0011101110101100000100",
			236 => "0000000000001110111001",
			237 => "0000000000001110111001",
			238 => "0001000011010100000100",
			239 => "0000000000001111110101",
			240 => "0000011111001100001000",
			241 => "0001000101100000000100",
			242 => "0000000000001111110101",
			243 => "0000000000001111110101",
			244 => "0001101011001100001100",
			245 => "0000111101000100001000",
			246 => "0010101010110000000100",
			247 => "0000000000001111110101",
			248 => "0000000000001111110101",
			249 => "0000000000001111110101",
			250 => "0011101110101000000100",
			251 => "0000000000001111110101",
			252 => "0000000000001111110101",
			253 => "0001000011010100000100",
			254 => "0000000000010000101001",
			255 => "0001101001100100010100",
			256 => "0000010110101000000100",
			257 => "0000000000010000101001",
			258 => "0000111101000100001100",
			259 => "0011110010000000001000",
			260 => "0001110110000100000100",
			261 => "0000000000010000101001",
			262 => "0000000000010000101001",
			263 => "0000000000010000101001",
			264 => "0000000000010000101001",
			265 => "0000000000010000101001",
			266 => "0001000011010100000100",
			267 => "0000000000010001101101",
			268 => "0000011111001100001000",
			269 => "0001000101100000000100",
			270 => "0000000000010001101101",
			271 => "0000000000010001101101",
			272 => "0001101011001100010000",
			273 => "0011111100010100001000",
			274 => "0010101010110000000100",
			275 => "0000000000010001101101",
			276 => "0000000000010001101101",
			277 => "0010100110011000000100",
			278 => "0000000000010001101101",
			279 => "0000000000010001101101",
			280 => "0011110111011000000100",
			281 => "0000000000010001101101",
			282 => "0000000000010001101101",
			283 => "0000100111011000000100",
			284 => "1111111000010010111001",
			285 => "0001101011001100001100",
			286 => "0000010110101000000100",
			287 => "0000000000010010111001",
			288 => "0011111110110100000100",
			289 => "0000001000010010111001",
			290 => "0000000000010010111001",
			291 => "0000011101011100001100",
			292 => "0001110011100000001000",
			293 => "0010100001010000000100",
			294 => "0000000000010010111001",
			295 => "1111111000010010111001",
			296 => "0000000000010010111001",
			297 => "0011101110101000001000",
			298 => "0010100001010000000100",
			299 => "0000000000010010111001",
			300 => "0000000000010010111001",
			301 => "0000000000010010111001",
			302 => "0001000010100100001000",
			303 => "0001000011110100000100",
			304 => "1111111000010100000101",
			305 => "0000000000010100000101",
			306 => "0000010110101000000100",
			307 => "0000000000010100000101",
			308 => "0001010101100100001100",
			309 => "0001101111000000001000",
			310 => "0010101100000100000100",
			311 => "0000001000010100000101",
			312 => "0000000000010100000101",
			313 => "0000000000010100000101",
			314 => "0000011101011100000100",
			315 => "0000000000010100000101",
			316 => "0011110111011000001000",
			317 => "0000101011111000000100",
			318 => "0000000000010100000101",
			319 => "0000001000010100000101",
			320 => "0000000000010100000101",
			321 => "0000100000010000010100",
			322 => "0000011111001100000100",
			323 => "1111111000010101101001",
			324 => "0001011011011100001100",
			325 => "0000100000010000001000",
			326 => "0011101110101100000100",
			327 => "0000000000010101101001",
			328 => "0000000000010101101001",
			329 => "0000000000010101101001",
			330 => "1111111000010101101001",
			331 => "0001101011001100001100",
			332 => "0000010110101000000100",
			333 => "0000000000010101101001",
			334 => "0000110011001000000100",
			335 => "0000001000010101101001",
			336 => "0000000000010101101001",
			337 => "0011111100000000010000",
			338 => "0010011010011000000100",
			339 => "0000000000010101101001",
			340 => "0000101011111000001000",
			341 => "0000111101000100000100",
			342 => "0000000000010101101001",
			343 => "0000000000010101101001",
			344 => "0000001000010101101001",
			345 => "1111111000010101101001",
			346 => "0000100000010000001100",
			347 => "0011001110001100001000",
			348 => "0001110001111100000100",
			349 => "1111111000010110110101",
			350 => "0000000000010110110101",
			351 => "0000000000010110110101",
			352 => "0011000100001000011000",
			353 => "0011001100110000000100",
			354 => "0000000000010110110101",
			355 => "0000101101101100010000",
			356 => "0000101011111000000100",
			357 => "0000000000010110110101",
			358 => "0001000011110100000100",
			359 => "0000000000010110110101",
			360 => "0000001100101100000100",
			361 => "0000000000010110110101",
			362 => "0000000000010110110101",
			363 => "0000000000010110110101",
			364 => "0000000000010110110101",
			365 => "0000100111011000000100",
			366 => "1111111000010111111001",
			367 => "0011111100000000011100",
			368 => "0000100110101100010000",
			369 => "0010100001010000001100",
			370 => "0011101110101100001000",
			371 => "0000011111001100000100",
			372 => "0000000000010111111001",
			373 => "0000000000010111111001",
			374 => "0000000000010111111001",
			375 => "0000000000010111111001",
			376 => "0010101100000100001000",
			377 => "0011000011011100000100",
			378 => "0000000000010111111001",
			379 => "0000001000010111111001",
			380 => "0000000000010111111001",
			381 => "1111111000010111111001",
			382 => "0000100000010000011000",
			383 => "0000011111001100000100",
			384 => "1111111000011001011101",
			385 => "0010110011100000001100",
			386 => "0000100000010000001000",
			387 => "0011101110101000000100",
			388 => "0000000000011001011101",
			389 => "0000000000011001011101",
			390 => "0000000000011001011101",
			391 => "0011100111110000000100",
			392 => "0000000000011001011101",
			393 => "1111111000011001011101",
			394 => "0011111100000000011000",
			395 => "0001101011001100001000",
			396 => "0000010110101000000100",
			397 => "0000000000011001011101",
			398 => "0000001000011001011101",
			399 => "0010011010011000000100",
			400 => "0000000000011001011101",
			401 => "0000101011111000001000",
			402 => "0011010101110100000100",
			403 => "0000000000011001011101",
			404 => "0000000000011001011101",
			405 => "0000001000011001011101",
			406 => "1111111000011001011101",
			407 => "0001000000010100000100",
			408 => "0000000000011010011001",
			409 => "0000010110101000000100",
			410 => "0000000000011010011001",
			411 => "0000101101101100010100",
			412 => "0001101111000000010000",
			413 => "0011000100001000001100",
			414 => "0001110110000100000100",
			415 => "0000000000011010011001",
			416 => "0011001100110000000100",
			417 => "0000000000011010011001",
			418 => "0000000000011010011001",
			419 => "0000000000011010011001",
			420 => "0000000000011010011001",
			421 => "0000000000011010011001",
			422 => "0000010110101000000100",
			423 => "0000000000011011101101",
			424 => "0001101011001100001100",
			425 => "0001001110111000000100",
			426 => "0000000000011011101101",
			427 => "0001101011001100000100",
			428 => "0000000000011011101101",
			429 => "0000000000011011101101",
			430 => "0010000110001000010100",
			431 => "0011000100001000010000",
			432 => "0001101011001100000100",
			433 => "0000000000011011101101",
			434 => "0001101001100100001000",
			435 => "0000000010011000000100",
			436 => "0000000000011011101101",
			437 => "0000000000011011101101",
			438 => "0000000000011011101101",
			439 => "0000000000011011101101",
			440 => "0000011101011100000100",
			441 => "0000000000011011101101",
			442 => "0000000000011011101101",
			443 => "0000011101101000000100",
			444 => "1111111000011101001001",
			445 => "0011000100001000100100",
			446 => "0011101001010100010100",
			447 => "0011010010001000001100",
			448 => "0011111001010000000100",
			449 => "0000000000011101001001",
			450 => "0010110001111100000100",
			451 => "0000000000011101001001",
			452 => "0000001000011101001001",
			453 => "0010011010011000000100",
			454 => "1111111000011101001001",
			455 => "0000001000011101001001",
			456 => "0011001110001100001000",
			457 => "0010100110011000000100",
			458 => "0000000000011101001001",
			459 => "1111111000011101001001",
			460 => "0011101110101000000100",
			461 => "0000001000011101001001",
			462 => "0000000000011101001001",
			463 => "0011100111110000000100",
			464 => "0000000000011101001001",
			465 => "1111111000011101001001",
			466 => "0010011110010100000100",
			467 => "1111111000011110100101",
			468 => "0000110110100000010100",
			469 => "0001000000010100000100",
			470 => "0000000000011110100101",
			471 => "0010001000101100001100",
			472 => "0011001100110000000100",
			473 => "0000000000011110100101",
			474 => "0000101111100100000100",
			475 => "0000000000011110100101",
			476 => "0000001000011110100101",
			477 => "0000000000011110100101",
			478 => "0011010000110100010100",
			479 => "0000101011111000001100",
			480 => "0010100110011000001000",
			481 => "0001001110111000000100",
			482 => "0000000000011110100101",
			483 => "0000000000011110100101",
			484 => "1111111000011110100101",
			485 => "0011110111011000000100",
			486 => "0000001000011110100101",
			487 => "0000000000011110100101",
			488 => "1111111000011110100101",
			489 => "0001000010100100001000",
			490 => "0001000011110100000100",
			491 => "1111111000100000011001",
			492 => "0000000000100000011001",
			493 => "0000100110101100010100",
			494 => "0010001011010100001100",
			495 => "0011111100010100001000",
			496 => "0000011111001100000100",
			497 => "0000000000100000011001",
			498 => "0000000000100000011001",
			499 => "0000000000100000011001",
			500 => "0010100110011000000100",
			501 => "0000000000100000011001",
			502 => "1111111000100000011001",
			503 => "0000110010110100010100",
			504 => "0010101100000100010000",
			505 => "0000100110101100000100",
			506 => "0000000000100000011001",
			507 => "0000101101101100001000",
			508 => "0001110110000100000100",
			509 => "0000000000100000011001",
			510 => "0000001000100000011001",
			511 => "0000000000100000011001",
			512 => "0000000000100000011001",
			513 => "0000011101011100000100",
			514 => "0000000000100000011001",
			515 => "0011011110101100000100",
			516 => "0000000000100000011001",
			517 => "0000000000100000011001",
			518 => "0000011101101000000100",
			519 => "1111111000100001100101",
			520 => "0011010000110100100000",
			521 => "0001001110111000000100",
			522 => "1111111000100001100101",
			523 => "0001010101100100001100",
			524 => "0011001100110000000100",
			525 => "0000000000100001100101",
			526 => "0000001100001000000100",
			527 => "0000001000100001100101",
			528 => "0000001000100001100101",
			529 => "0010011010011000000100",
			530 => "1111111000100001100101",
			531 => "0011000110000100000100",
			532 => "0000000000100001100101",
			533 => "0000011101011100000100",
			534 => "0000000000100001100101",
			535 => "0000001000100001100101",
			536 => "1111111000100001100101",
			537 => "0000011101101000000100",
			538 => "1111111000100011000001",
			539 => "0011010000110100101000",
			540 => "0000101011111000011100",
			541 => "0011101001010100001100",
			542 => "0010101010110000001000",
			543 => "0000100111011000000100",
			544 => "0000000000100011000001",
			545 => "0000001000100011000001",
			546 => "0000000000100011000001",
			547 => "0011001110001100001000",
			548 => "0010100110011000000100",
			549 => "0000000000100011000001",
			550 => "1111111000100011000001",
			551 => "0000110111100000000100",
			552 => "0000000000100011000001",
			553 => "0000000000100011000001",
			554 => "0001100100111100001000",
			555 => "0010100001010100000100",
			556 => "0000001000100011000001",
			557 => "0000000000100011000001",
			558 => "0000000000100011000001",
			559 => "1111111000100011000001",
			560 => "0000101111010100001000",
			561 => "0000100111011000000100",
			562 => "1111111000100100110101",
			563 => "0000000000100100110101",
			564 => "0011101010111000010000",
			565 => "0000010110101000000100",
			566 => "0000000000100100110101",
			567 => "0010110000001100000100",
			568 => "0000011000100100110101",
			569 => "0000010111100100000100",
			570 => "0000000000100100110101",
			571 => "0000001000100100110101",
			572 => "0011101110101000100000",
			573 => "0010001011010100001100",
			574 => "0001111101010100000100",
			575 => "0000001000100100110101",
			576 => "0001110111001000000100",
			577 => "0000000000100100110101",
			578 => "0000000000100100110101",
			579 => "0000100110101100001100",
			580 => "0010111010111000001000",
			581 => "0000011101101000000100",
			582 => "0000000000100100110101",
			583 => "0000000000100100110101",
			584 => "1111111000100100110101",
			585 => "0010000001110100000100",
			586 => "0000001000100100110101",
			587 => "0000000000100100110101",
			588 => "1111111000100100110101",
			589 => "0000100111011000000100",
			590 => "1111111000100110010001",
			591 => "0011111100000000101000",
			592 => "0010001011010100001100",
			593 => "0001001110111000000100",
			594 => "0000000000100110010001",
			595 => "0000011111001100000100",
			596 => "0000000000100110010001",
			597 => "0000001000100110010001",
			598 => "0001101101011000001000",
			599 => "0000010110101000000100",
			600 => "0000000000100110010001",
			601 => "0000000000100110010001",
			602 => "0000101000100000001000",
			603 => "0001101011001100000100",
			604 => "0000000000100110010001",
			605 => "0000000000100110010001",
			606 => "0010011010011000001000",
			607 => "0001101011001100000100",
			608 => "0000000000100110010001",
			609 => "0000000000100110010001",
			610 => "0000000000100110010001",
			611 => "0000000000100110010001",
			612 => "0000101111010100001000",
			613 => "0000100111011000000100",
			614 => "1111111000101000010101",
			615 => "1111111000101000010101",
			616 => "0011000100001000101000",
			617 => "0000011101101000001100",
			618 => "0011000110000100000100",
			619 => "1111111000101000010101",
			620 => "0000001100101100000100",
			621 => "0000011000101000010101",
			622 => "1111111000101000010101",
			623 => "0000110001011000000100",
			624 => "0001011000101000010101",
			625 => "0000110111110000001000",
			626 => "0010100101000100000100",
			627 => "0000011000101000010101",
			628 => "0000000000101000010101",
			629 => "0010011010011000001000",
			630 => "0010100001010000000100",
			631 => "0000000000101000010101",
			632 => "1111111000101000010101",
			633 => "0000111001011100000100",
			634 => "0000001000101000010101",
			635 => "1111111000101000010101",
			636 => "0001110111001000001100",
			637 => "0001010101100100000100",
			638 => "0000000000101000010101",
			639 => "0011000100001000000100",
			640 => "0000000000101000010101",
			641 => "0000001000101000010101",
			642 => "0011000100001000000100",
			643 => "0000000000101000010101",
			644 => "1111111000101000010101",
			645 => "0000101111010100001100",
			646 => "0000100111011000000100",
			647 => "1111111000101010000001",
			648 => "0000100110111100000100",
			649 => "0000000000101010000001",
			650 => "0000000000101010000001",
			651 => "0011111100000000101000",
			652 => "0010011110010100000100",
			653 => "1111111000101010000001",
			654 => "0001010101100100001100",
			655 => "0011000011011100000100",
			656 => "0000000000101010000001",
			657 => "0010100001010100000100",
			658 => "0000001000101010000001",
			659 => "0000000000101010000001",
			660 => "0000100110101100001100",
			661 => "0010001011010100001000",
			662 => "0000110111100000000100",
			663 => "0000001000101010000001",
			664 => "0000000000101010000001",
			665 => "1111111000101010000001",
			666 => "0010011010011000000100",
			667 => "0000000000101010000001",
			668 => "0001110100001000000100",
			669 => "0000000000101010000001",
			670 => "0000001000101010000001",
			671 => "1111111000101010000001",
			672 => "0000011101101000000100",
			673 => "1111111000101011011101",
			674 => "0011010000110100101000",
			675 => "0001001110111000000100",
			676 => "1111111000101011011101",
			677 => "0001010101100100001100",
			678 => "0000000100000000001000",
			679 => "0010100110011100000100",
			680 => "0000001000101011011101",
			681 => "0000000000101011011101",
			682 => "0000010000101011011101",
			683 => "0000011101011100001100",
			684 => "0010101010110000000100",
			685 => "0000000000101011011101",
			686 => "0011110010000000000100",
			687 => "1111111000101011011101",
			688 => "0000000000101011011101",
			689 => "0011001110001100001000",
			690 => "0000101011111000000100",
			691 => "0000000000101011011101",
			692 => "0000000000101011011101",
			693 => "0000001000101011011101",
			694 => "1111111000101011011101",
			695 => "0000101111010100000100",
			696 => "1111111000101101011011",
			697 => "0011000100001000101100",
			698 => "0000011101101000000100",
			699 => "1111111000101101011011",
			700 => "0011101001010100010000",
			701 => "0010001000101100001100",
			702 => "0000011111001100000100",
			703 => "0000010000101101011011",
			704 => "0000011101011100000100",
			705 => "0000000000101101011011",
			706 => "0000001000101101011011",
			707 => "1111111000101101011011",
			708 => "0000011001011000001100",
			709 => "0001001101110100001000",
			710 => "0001000000010100000100",
			711 => "1111111000101101011011",
			712 => "0000000000101101011011",
			713 => "1111110000101101011011",
			714 => "0011101110101000001000",
			715 => "0000100110101100000100",
			716 => "0000000000101101011011",
			717 => "0000010000101101011011",
			718 => "1111111000101101011011",
			719 => "0001110111001000001100",
			720 => "0011100111110000001000",
			721 => "0011101000110000000100",
			722 => "0000000000101101011011",
			723 => "0000000000101101011011",
			724 => "1111111000101101011011",
			725 => "1111111000101101011011",
			726 => "0000000000101101011101",
			727 => "0000000000101101100001",
			728 => "0000000000101101100101",
			729 => "0000000000101101101001",
			730 => "0000000000101101101101",
			731 => "0000000000101101110001",
			732 => "0000000000101101110101",
			733 => "0000000000101101111001",
			734 => "0000000000101101111101",
			735 => "0000000000101110000001",
			736 => "0000000000101110000101",
			737 => "0000000000101110001001",
			738 => "0000000000101110001101",
			739 => "0000000000101110010001",
			740 => "0000000000101110010101",
			741 => "0000000000101110011001",
			742 => "0000000000101110011101",
			743 => "0000000000101110100001",
			744 => "0000000000101110100101",
			745 => "0000000000101110101001",
			746 => "0000000000101110101101",
			747 => "0000000000101110110001",
			748 => "0000000000101110110101",
			749 => "0000000000101110111001",
			750 => "0000000000101110111101",
			751 => "0000000000101111000001",
			752 => "0000000000101111000101",
			753 => "0000000000101111001001",
			754 => "0000000000101111001101",
			755 => "0001000100111000000100",
			756 => "0000000000101111011001",
			757 => "0000000000101111011001",
			758 => "0001000011011000000100",
			759 => "0000000000101111100101",
			760 => "0000000000101111100101",
			761 => "0000100110101100000100",
			762 => "0000000000101111110001",
			763 => "0000000000101111110001",
			764 => "0001000011111000000100",
			765 => "0000000000101111111101",
			766 => "0000000000101111111101",
			767 => "0000011111001100000100",
			768 => "0000000000110000001001",
			769 => "0000000000110000001001",
			770 => "0000101011101100000100",
			771 => "0000000000110000010101",
			772 => "0000000000110000010101",
			773 => "0001000011111000000100",
			774 => "0000000000110000100001",
			775 => "0000000000110000100001",
			776 => "0001000000010100000100",
			777 => "0000000000110000110101",
			778 => "0001001010010000000100",
			779 => "0000000000110000110101",
			780 => "0000000000110000110101",
			781 => "0001000011010100000100",
			782 => "0000000000110001001001",
			783 => "0001001010010000000100",
			784 => "0000000000110001001001",
			785 => "0000000000110001001001",
			786 => "0001000010100100000100",
			787 => "0000000000110001011101",
			788 => "0001001010010000000100",
			789 => "0000000000110001011101",
			790 => "0000000000110001011101",
			791 => "0000101011111000000100",
			792 => "0000000000110001110001",
			793 => "0000101101101100000100",
			794 => "0000000000110001110001",
			795 => "0000000000110001110001",
			796 => "0000100110101100000100",
			797 => "0000000000110010000101",
			798 => "0000101111101000000100",
			799 => "0000000000110010000101",
			800 => "0000000000110010000101",
			801 => "0001000011011000001000",
			802 => "0010100110011000000100",
			803 => "0000000000110010011001",
			804 => "0000000000110010011001",
			805 => "0000000000110010011001",
			806 => "0000011111001100000100",
			807 => "0000000000110010110101",
			808 => "0011101001010100001000",
			809 => "0001111101111000000100",
			810 => "0000000000110010110101",
			811 => "0000000000110010110101",
			812 => "0000000000110010110101",
			813 => "0001000101100000001100",
			814 => "0000011101011100001000",
			815 => "0010011101011000000100",
			816 => "0000000000110011010001",
			817 => "0000000000110011010001",
			818 => "0000000000110011010001",
			819 => "0000000000110011010001",
			820 => "0001000011010100000100",
			821 => "0000000000110011101101",
			822 => "0000100000010000000100",
			823 => "0000000000110011101101",
			824 => "0000101111101000000100",
			825 => "0000000000110011101101",
			826 => "0000000000110011101101",
			827 => "0010011101011000001100",
			828 => "0001000100111000001000",
			829 => "0000011101011100000100",
			830 => "0000000000110100001001",
			831 => "0000000000110100001001",
			832 => "0000000000110100001001",
			833 => "0000000000110100001001",
			834 => "0000011101011100001100",
			835 => "0000101011101100001000",
			836 => "0010011101011000000100",
			837 => "0000000000110100100101",
			838 => "0000000000110100100101",
			839 => "0000000000110100100101",
			840 => "0000000000110100100101",
			841 => "0000011111001100000100",
			842 => "0000000000110101001001",
			843 => "0011011001010100001100",
			844 => "0011000000001100001000",
			845 => "0011101110101000000100",
			846 => "0000000000110101001001",
			847 => "0000000000110101001001",
			848 => "0000000000110101001001",
			849 => "0000000000110101001001",
			850 => "0001000000010100000100",
			851 => "0000000000110101101101",
			852 => "0010011011111100000100",
			853 => "0000000000110101101101",
			854 => "0000101111101000001000",
			855 => "0001111110001100000100",
			856 => "0000000000110101101101",
			857 => "0000000000110101101101",
			858 => "0000000000110101101101",
			859 => "0001000011010100000100",
			860 => "0000000000110110010001",
			861 => "0000100110101100000100",
			862 => "0000000000110110010001",
			863 => "0000100011000000001000",
			864 => "0001001010010000000100",
			865 => "0000000000110110010001",
			866 => "0000000000110110010001",
			867 => "0000000000110110010001",
			868 => "0001000011011000000100",
			869 => "0000000000110110110101",
			870 => "0011010100010000001100",
			871 => "0011011000011000000100",
			872 => "0000000000110110110101",
			873 => "0010111000000000000100",
			874 => "0000000000110110110101",
			875 => "0000000000110110110101",
			876 => "0000000000110110110101",
			877 => "0000011111001100001000",
			878 => "0001000100111000000100",
			879 => "0000000000110111100001",
			880 => "0000000000110111100001",
			881 => "0011100111110000001100",
			882 => "0001111101111000000100",
			883 => "0000000000110111100001",
			884 => "0001101001100100000100",
			885 => "0000000000110111100001",
			886 => "0000000000110111100001",
			887 => "0000000000110111100001",
			888 => "0000011101011100001000",
			889 => "0000101011101100000100",
			890 => "0000000000111000001101",
			891 => "0000000000111000001101",
			892 => "0010110001101000001100",
			893 => "0001111100101000000100",
			894 => "0000000000111000001101",
			895 => "0001001110111000000100",
			896 => "0000000000111000001101",
			897 => "0000000000111000001101",
			898 => "0000000000111000001101",
			899 => "0000100110101100001100",
			900 => "0000000011111100000100",
			901 => "0000000000111001000001",
			902 => "0001101001100100000100",
			903 => "0000000000111001000001",
			904 => "0000000000111001000001",
			905 => "0011111100010000001100",
			906 => "0000011111001100000100",
			907 => "0000000000111001000001",
			908 => "0000100001011100000100",
			909 => "0000000000111001000001",
			910 => "0000000000111001000001",
			911 => "0000000000111001000001",
			912 => "0001000011110100000100",
			913 => "0000000000111001110101",
			914 => "0010110011100000001100",
			915 => "0000011111001100000100",
			916 => "0000000000111001110101",
			917 => "0001111101111000000100",
			918 => "0000000000111001110101",
			919 => "0000000000111001110101",
			920 => "0010001011010100000100",
			921 => "0000000000111001110101",
			922 => "0011010101110100000100",
			923 => "0000000000111001110101",
			924 => "0000000000111001110101",
			925 => "0010010100110100000100",
			926 => "0000000000111010100001",
			927 => "0011011001010100010000",
			928 => "0011000000001100001100",
			929 => "0001111110001100000100",
			930 => "0000000000111010100001",
			931 => "0011101110101000000100",
			932 => "0000000000111010100001",
			933 => "0000000000111010100001",
			934 => "0000000000111010100001",
			935 => "0000000000111010100001",
			936 => "0001000000010100000100",
			937 => "0000000000111011001101",
			938 => "0011001100110000000100",
			939 => "0000000000111011001101",
			940 => "0000101101101100001100",
			941 => "0001001010010000001000",
			942 => "0011000100001000000100",
			943 => "0000000000111011001101",
			944 => "0000000000111011001101",
			945 => "0000000000111011001101",
			946 => "0000000000111011001101",
			947 => "0001110110000100001000",
			948 => "0000011111001100000100",
			949 => "1111111000111100010001",
			950 => "0000000000111100010001",
			951 => "0000111101000100010000",
			952 => "0000011111001100000100",
			953 => "0000000000111100010001",
			954 => "0001111101111000000100",
			955 => "0000000000111100010001",
			956 => "0011000000001100000100",
			957 => "0000001000111100010001",
			958 => "0000000000111100010001",
			959 => "0001010101100100000100",
			960 => "0000000000111100010001",
			961 => "0010100001010000000100",
			962 => "0000000000111100010001",
			963 => "0000000000111100010001",
			964 => "0001000011111000011000",
			965 => "0010011100011000000100",
			966 => "1111111000111101011101",
			967 => "0011100111110000001000",
			968 => "0010011010011000000100",
			969 => "0000000000111101011101",
			970 => "0000001000111101011101",
			971 => "0010110011100000000100",
			972 => "0000000000111101011101",
			973 => "0011000110000100000100",
			974 => "0000000000111101011101",
			975 => "1111111000111101011101",
			976 => "0010101100000100001100",
			977 => "0011010001011000001000",
			978 => "0000101111100100000100",
			979 => "0000000000111101011101",
			980 => "0000001000111101011101",
			981 => "0000000000111101011101",
			982 => "0000000000111101011101",
			983 => "0001000000010100000100",
			984 => "0000000000111110011001",
			985 => "0000100110101100001000",
			986 => "0010001011010100000100",
			987 => "0000000000111110011001",
			988 => "0000000000111110011001",
			989 => "0001100100111100010000",
			990 => "0011000011011100000100",
			991 => "0000000000111110011001",
			992 => "0010101100000100001000",
			993 => "0011000100001000000100",
			994 => "0000000000111110011001",
			995 => "0000000000111110011001",
			996 => "0000000000111110011001",
			997 => "0000000000111110011001",
			998 => "0000101000001100001100",
			999 => "0011001110001100001000",
			1000 => "0001111100101000000100",
			1001 => "1111111000111111100101",
			1002 => "0000000000111111100101",
			1003 => "0000000000111111100101",
			1004 => "0011111100000000011000",
			1005 => "0000011111001100010000",
			1006 => "0011111110000100001100",
			1007 => "0000001100101100001000",
			1008 => "0000001001110000000100",
			1009 => "0000000000111111100101",
			1010 => "0000000000111111100101",
			1011 => "0000000000111111100101",
			1012 => "0000000000111111100101",
			1013 => "0000101011111000000100",
			1014 => "0000000000111111100101",
			1015 => "0000000000111111100101",
			1016 => "0000000000111111100101",
			1017 => "0000011111001100100000",
			1018 => "0000011111001100011000",
			1019 => "0000101011111000000100",
			1020 => "1011111001000000111001",
			1021 => "0000100110101100001000",
			1022 => "0000010110000000000100",
			1023 => "1011111001000000111001",
			1024 => "1100110001000000111001",
			1025 => "0001101011001100001000",
			1026 => "0000010110101000000100",
			1027 => "1011111001000000111001",
			1028 => "1100110001000000111001",
			1029 => "1011111001000000111001",
			1030 => "0011100100010000000100",
			1031 => "1110011001000000111001",
			1032 => "1011111001000000111001",
			1033 => "0011101110101100000100",
			1034 => "0001101001000000111001",
			1035 => "0011101110101000000100",
			1036 => "1101100001000000111001",
			1037 => "1011111001000000111001",
			1038 => "0001000010100100001000",
			1039 => "0001000011110100000100",
			1040 => "1111111001000010000101",
			1041 => "0000000001000010000101",
			1042 => "0000010110101000000100",
			1043 => "0000000001000010000101",
			1044 => "0011010101110100001100",
			1045 => "0001101111000000001000",
			1046 => "0010101100000100000100",
			1047 => "0000001001000010000101",
			1048 => "0000000001000010000101",
			1049 => "0000000001000010000101",
			1050 => "0000011101011100000100",
			1051 => "0000000001000010000101",
			1052 => "0001100100111100001000",
			1053 => "0000101011111000000100",
			1054 => "0000000001000010000101",
			1055 => "0000000001000010000101",
			1056 => "0000000001000010000101",
			1057 => "0000100000010000001100",
			1058 => "0010011111000000001000",
			1059 => "0011001110001100000100",
			1060 => "1111111001000011011001",
			1061 => "0000000001000011011001",
			1062 => "0000000001000011011001",
			1063 => "0011110010000100011000",
			1064 => "0000100110101100000100",
			1065 => "0000000001000011011001",
			1066 => "0011001100110000000100",
			1067 => "0000000001000011011001",
			1068 => "0010101100000100001100",
			1069 => "0000100001011100001000",
			1070 => "0001101111000000000100",
			1071 => "0000001001000011011001",
			1072 => "0000000001000011011001",
			1073 => "0000000001000011011001",
			1074 => "0000000001000011011001",
			1075 => "0011111100000000000100",
			1076 => "0000000001000011011001",
			1077 => "0000000001000011011001",
			1078 => "0000101000001100001100",
			1079 => "0001111100101000001000",
			1080 => "0011001110001100000100",
			1081 => "1111111001000100100101",
			1082 => "0000000001000100100101",
			1083 => "0000000001000100100101",
			1084 => "0011000100001000011000",
			1085 => "0011001100110000000100",
			1086 => "0000000001000100100101",
			1087 => "0000101011111000000100",
			1088 => "0000000001000100100101",
			1089 => "0000101101101100001100",
			1090 => "0001000011110100000100",
			1091 => "0000000001000100100101",
			1092 => "0000001100101100000100",
			1093 => "0000000001000100100101",
			1094 => "0000000001000100100101",
			1095 => "0000000001000100100101",
			1096 => "0000000001000100100101",
			1097 => "0000101000001100001000",
			1098 => "0011001110001100000100",
			1099 => "0000000001000101101001",
			1100 => "0000000001000101101001",
			1101 => "0011000100001000011000",
			1102 => "0011001100110000000100",
			1103 => "0000000001000101101001",
			1104 => "0000101011111000000100",
			1105 => "0000000001000101101001",
			1106 => "0000101101101100001100",
			1107 => "0001000011110100000100",
			1108 => "0000000001000101101001",
			1109 => "0000001100101100000100",
			1110 => "0000000001000101101001",
			1111 => "0000000001000101101001",
			1112 => "0000000001000101101001",
			1113 => "0000000001000101101001",
			1114 => "0001110110000100000100",
			1115 => "0000000001000110111101",
			1116 => "0000111101000100010100",
			1117 => "0010100101000100010000",
			1118 => "0010011110010100000100",
			1119 => "0000000001000110111101",
			1120 => "0011001100110000000100",
			1121 => "0000000001000110111101",
			1122 => "0001000000010100000100",
			1123 => "0000000001000110111101",
			1124 => "0000000001000110111101",
			1125 => "0000000001000110111101",
			1126 => "0001101001100100001000",
			1127 => "0010110011100000000100",
			1128 => "0000000001000110111101",
			1129 => "0000000001000110111101",
			1130 => "0001101001100100001000",
			1131 => "0010110110100100000100",
			1132 => "0000000001000110111101",
			1133 => "0000000001000110111101",
			1134 => "0000000001000110111101",
			1135 => "0001000000010100000100",
			1136 => "0000000001000111111001",
			1137 => "0000010110101000000100",
			1138 => "0000000001000111111001",
			1139 => "0000101101101100010100",
			1140 => "0001101111000000010000",
			1141 => "0011000100001000001100",
			1142 => "0001110110000100000100",
			1143 => "0000000001000111111001",
			1144 => "0011001100110000000100",
			1145 => "0000000001000111111001",
			1146 => "0000000001000111111001",
			1147 => "0000000001000111111001",
			1148 => "0000000001000111111001",
			1149 => "0000000001000111111001",
			1150 => "0001110110000100001000",
			1151 => "0000011111001100000100",
			1152 => "1111111001001001011101",
			1153 => "0000000001001001011101",
			1154 => "0011000100001000100100",
			1155 => "0000011101011100011000",
			1156 => "0001101011001100001100",
			1157 => "0011111110101000000100",
			1158 => "0000000001001001011101",
			1159 => "0000001101010000000100",
			1160 => "0000000001001001011101",
			1161 => "0000001001001001011101",
			1162 => "0001010110110100001000",
			1163 => "0010011101011000000100",
			1164 => "0000000001001001011101",
			1165 => "0000000001001001011101",
			1166 => "0000000001001001011101",
			1167 => "0011101110101000001000",
			1168 => "0010000110001000000100",
			1169 => "0000001001001001011101",
			1170 => "0000000001001001011101",
			1171 => "0000000001001001011101",
			1172 => "0001111101010100000100",
			1173 => "0000000001001001011101",
			1174 => "0000000001001001011101",
			1175 => "0000011101101000000100",
			1176 => "1111111001001010100001",
			1177 => "0011010000110100011100",
			1178 => "0001001110111000000100",
			1179 => "1111111001001010100001",
			1180 => "0001010101100100001000",
			1181 => "0011001100110000000100",
			1182 => "0000000001001010100001",
			1183 => "0000001001001010100001",
			1184 => "0010011010011000000100",
			1185 => "1111111001001010100001",
			1186 => "0011000110000100000100",
			1187 => "0000000001001010100001",
			1188 => "0000011101011100000100",
			1189 => "0000000001001010100001",
			1190 => "0000001001001010100001",
			1191 => "1111111001001010100001",
			1192 => "0000011101101000000100",
			1193 => "1111111001001011111101",
			1194 => "0011100111110000010100",
			1195 => "0010001000101100010000",
			1196 => "0000100111011000000100",
			1197 => "0000000001001011111101",
			1198 => "0000101011101100001000",
			1199 => "0011110010000000000100",
			1200 => "0000001001001011111101",
			1201 => "0000000001001011111101",
			1202 => "0000001001001011111101",
			1203 => "0000000001001011111101",
			1204 => "0011010000110100010100",
			1205 => "0000101011111000001100",
			1206 => "0010100110011000001000",
			1207 => "0001001110111000000100",
			1208 => "0000000001001011111101",
			1209 => "0000000001001011111101",
			1210 => "1111111001001011111101",
			1211 => "0011110111011000000100",
			1212 => "0000001001001011111101",
			1213 => "0000000001001011111101",
			1214 => "1111111001001011111101",
			1215 => "0001000010100100000100",
			1216 => "1111111001001101100001",
			1217 => "0011100111110000011100",
			1218 => "0000010110101000000100",
			1219 => "0000000001001101100001",
			1220 => "0011010001011000001100",
			1221 => "0001101001100100001000",
			1222 => "0011001100110000000100",
			1223 => "0000000001001101100001",
			1224 => "0000001001001101100001",
			1225 => "0000000001001101100001",
			1226 => "0010101100011100001000",
			1227 => "0011111001011100000100",
			1228 => "0000000001001101100001",
			1229 => "0000000001001101100001",
			1230 => "0000000001001101100001",
			1231 => "0010001011010100001000",
			1232 => "0001111101010100000100",
			1233 => "0000000001001101100001",
			1234 => "0000000001001101100001",
			1235 => "0011010101110100000100",
			1236 => "0000000001001101100001",
			1237 => "0010111000000000000100",
			1238 => "1111111001001101100001",
			1239 => "0000000001001101100001",
			1240 => "0000100111011000000100",
			1241 => "1111111001001110101101",
			1242 => "0011111100000000100000",
			1243 => "0010011110010100000100",
			1244 => "1111111001001110101101",
			1245 => "0000101011111000010100",
			1246 => "0010001011010100001000",
			1247 => "0011101110101100000100",
			1248 => "0000001001001110101101",
			1249 => "0000000001001110101101",
			1250 => "0001010101100100001000",
			1251 => "0010010100110100000100",
			1252 => "0000000001001110101101",
			1253 => "0000000001001110101101",
			1254 => "1111111001001110101101",
			1255 => "0010100001010100000100",
			1256 => "0000001001001110101101",
			1257 => "0000000001001110101101",
			1258 => "1111111001001110101101",
			1259 => "0000011101101000000100",
			1260 => "1111111001010000010001",
			1261 => "0011010000110100101000",
			1262 => "0000101011111000011000",
			1263 => "0010001011010100010000",
			1264 => "0000001000110000000100",
			1265 => "0000000001010000010001",
			1266 => "0011110010000000001000",
			1267 => "0000011111001100000100",
			1268 => "0000000001010000010001",
			1269 => "0000001001010000010001",
			1270 => "0000000001010000010001",
			1271 => "0001010101100100000100",
			1272 => "0000000001010000010001",
			1273 => "1111111001010000010001",
			1274 => "0011001100110000000100",
			1275 => "0000000001010000010001",
			1276 => "0010001000101100001000",
			1277 => "0011110111011000000100",
			1278 => "0000001001010000010001",
			1279 => "0000000001010000010001",
			1280 => "0000000001010000010001",
			1281 => "0001011011110100000100",
			1282 => "0000000001010000010001",
			1283 => "1111111001010000010001",
			1284 => "0000101111010100001000",
			1285 => "0000100111011000000100",
			1286 => "1111111001010010000101",
			1287 => "0000000001010010000101",
			1288 => "0001101011001100010000",
			1289 => "0001111101010100001100",
			1290 => "0000010110101000000100",
			1291 => "0000000001010010000101",
			1292 => "0011001100110000000100",
			1293 => "0000000001010010000101",
			1294 => "0000001001010010000101",
			1295 => "0000000001010010000101",
			1296 => "0011111100000000100000",
			1297 => "0000011101011100010000",
			1298 => "0011111100010100001000",
			1299 => "0010100001010000000100",
			1300 => "0000000001010010000101",
			1301 => "1111111001010010000101",
			1302 => "0010011010011000000100",
			1303 => "0000000001010010000101",
			1304 => "0000000001010010000101",
			1305 => "0000101011111000001100",
			1306 => "0000111101000100000100",
			1307 => "0000000001010010000101",
			1308 => "0011001110001100000100",
			1309 => "0000000001010010000101",
			1310 => "0000000001010010000101",
			1311 => "0000001001010010000101",
			1312 => "1111111001010010000101",
			1313 => "0000100111011000000100",
			1314 => "1111111001010011110001",
			1315 => "0011001010111100101100",
			1316 => "0000101011111000011100",
			1317 => "0010001011010100001100",
			1318 => "0011101110101100001000",
			1319 => "0000011111001100000100",
			1320 => "0000000001010011110001",
			1321 => "0000001001010011110001",
			1322 => "0000000001010011110001",
			1323 => "0011001110001100001000",
			1324 => "0010100110011000000100",
			1325 => "0000000001010011110001",
			1326 => "1111111001010011110001",
			1327 => "0000110010001000000100",
			1328 => "0000000001010011110001",
			1329 => "0000000001010011110001",
			1330 => "0010100001010100001100",
			1331 => "0001000011110100000100",
			1332 => "0000000001010011110001",
			1333 => "0011000011011100000100",
			1334 => "0000000001010011110001",
			1335 => "0000001001010011110001",
			1336 => "0000000001010011110001",
			1337 => "0011001010111100000100",
			1338 => "0000000001010011110001",
			1339 => "1111111001010011110001",
			1340 => "0001000011110100001100",
			1341 => "0001000011010100000100",
			1342 => "1111111001010101110101",
			1343 => "0001000011010100000100",
			1344 => "0000000001010101110101",
			1345 => "1111111001010101110101",
			1346 => "0010000010101000100100",
			1347 => "0010011110010100000100",
			1348 => "1111111001010101110101",
			1349 => "0011100111110000001100",
			1350 => "0001010101100100000100",
			1351 => "0000001001010101110101",
			1352 => "0001010101100100000100",
			1353 => "0000000001010101110101",
			1354 => "0000001001010101110101",
			1355 => "0010001011010100001000",
			1356 => "0001101011001100000100",
			1357 => "0000000001010101110101",
			1358 => "0000001001010101110101",
			1359 => "0001101001100100000100",
			1360 => "1111111001010101110101",
			1361 => "0011101110101100000100",
			1362 => "0000001001010101110101",
			1363 => "0000000001010101110101",
			1364 => "0010100001110000010000",
			1365 => "0010011011111100000100",
			1366 => "1111111001010101110101",
			1367 => "0001111101111000000100",
			1368 => "0000010001010101110101",
			1369 => "0010100101000100000100",
			1370 => "0000000001010101110101",
			1371 => "0000000001010101110101",
			1372 => "1111111001010101110101",
			1373 => "0000100110111100000100",
			1374 => "1111111001010111101001",
			1375 => "0011000100001000100100",
			1376 => "0011000011011100001000",
			1377 => "0001111101111000000100",
			1378 => "1111111001010111101001",
			1379 => "0000000001010111101001",
			1380 => "0010101100000100011000",
			1381 => "0011100001101000001000",
			1382 => "0000100110101100000100",
			1383 => "0000001001010111101001",
			1384 => "0000100001010111101001",
			1385 => "0001010101100100001000",
			1386 => "0000011111001100000100",
			1387 => "0000000001010111101001",
			1388 => "0000001001010111101001",
			1389 => "0010011010011000000100",
			1390 => "1111111001010111101001",
			1391 => "0000001001010111101001",
			1392 => "1111111001010111101001",
			1393 => "0001110111001000001100",
			1394 => "0001010101100100000100",
			1395 => "0000000001010111101001",
			1396 => "0011000100001000000100",
			1397 => "0000000001010111101001",
			1398 => "0000001001010111101001",
			1399 => "0011000100001000000100",
			1400 => "0000000001010111101001",
			1401 => "1111111001010111101001",
			1402 => "0000011101101000000100",
			1403 => "1111111001011001110101",
			1404 => "0011101001010100100000",
			1405 => "0001010101100100010000",
			1406 => "0011101001001000000100",
			1407 => "0000010001011001110101",
			1408 => "0001000000010100000100",
			1409 => "0000000001011001110101",
			1410 => "0010100110011100000100",
			1411 => "0000001001011001110101",
			1412 => "0000000001011001110101",
			1413 => "0000011101011100001100",
			1414 => "0011111100010100001000",
			1415 => "0011101011011100000100",
			1416 => "0000000001011001110101",
			1417 => "1111111001011001110101",
			1418 => "0000000001011001110101",
			1419 => "0000001001011001110101",
			1420 => "0011010000110100100000",
			1421 => "0011001110001100010100",
			1422 => "0010001011010100001000",
			1423 => "0001000110001100000100",
			1424 => "0000000001011001110101",
			1425 => "0000000001011001110101",
			1426 => "0011010100010000001000",
			1427 => "0001010100000100000100",
			1428 => "0000000001011001110101",
			1429 => "0000000001011001110101",
			1430 => "1111111001011001110101",
			1431 => "0001000000010100000100",
			1432 => "0000000001011001110101",
			1433 => "0010011111000000000100",
			1434 => "0000000001011001110101",
			1435 => "0000001001011001110101",
			1436 => "1111111001011001110101",
			1437 => "0000101111010100000100",
			1438 => "1111111001011011111011",
			1439 => "0011000100001000110000",
			1440 => "0010011110010100000100",
			1441 => "1111111001011011111011",
			1442 => "0011101001010100010100",
			1443 => "0010001000101100010000",
			1444 => "0000011111001100001000",
			1445 => "0011111110010000000100",
			1446 => "0000010001011011111011",
			1447 => "0000001001011011111011",
			1448 => "0000011101011100000100",
			1449 => "0000000001011011111011",
			1450 => "0000001001011011111011",
			1451 => "1111111001011011111011",
			1452 => "0000011001011000001100",
			1453 => "0010001100000100000100",
			1454 => "0000000001011011111011",
			1455 => "0010110100011000000100",
			1456 => "1111111001011011111011",
			1457 => "1111110001011011111011",
			1458 => "0011101110101000001000",
			1459 => "0011001110001100000100",
			1460 => "0000000001011011111011",
			1461 => "0000001001011011111011",
			1462 => "1111111001011011111011",
			1463 => "0001110111001000001100",
			1464 => "0011100111110000001000",
			1465 => "0011101000110000000100",
			1466 => "0000000001011011111011",
			1467 => "0000000001011011111011",
			1468 => "1111111001011011111011",
			1469 => "1111111001011011111011",
			1470 => "0000000001011011111101",
			1471 => "0000000001011100000001",
			1472 => "0000000001011100000101",
			1473 => "0000000001011100001001",
			1474 => "0000000001011100001101",
			1475 => "0000000001011100010001",
			1476 => "0000000001011100010101",
			1477 => "0000000001011100011001",
			1478 => "0000000001011100011101",
			1479 => "0000000001011100100001",
			1480 => "0000000001011100100101",
			1481 => "0000000001011100101001",
			1482 => "0000000001011100101101",
			1483 => "0000000001011100110001",
			1484 => "0000000001011100110101",
			1485 => "0000000001011100111001",
			1486 => "0000000001011100111101",
			1487 => "0000000001011101000001",
			1488 => "0000000001011101000101",
			1489 => "0000000001011101001001",
			1490 => "0000000001011101001101",
			1491 => "0000000001011101010001",
			1492 => "0000000001011101010101",
			1493 => "0000000001011101011001",
			1494 => "0000000001011101011101",
			1495 => "0000000001011101100001",
			1496 => "0000000001011101100101",
			1497 => "0000000001011101101001",
			1498 => "0000000001011101101101",
			1499 => "0001000100111000000100",
			1500 => "0000000001011101111001",
			1501 => "0000000001011101111001",
			1502 => "0001000011011000000100",
			1503 => "0000000001011110000101",
			1504 => "0000000001011110000101",
			1505 => "0000100110101100000100",
			1506 => "0000000001011110010001",
			1507 => "0000000001011110010001",
			1508 => "0000001100001000000100",
			1509 => "0000000001011110011101",
			1510 => "0000000001011110011101",
			1511 => "0000011111001100000100",
			1512 => "0000000001011110101001",
			1513 => "0000000001011110101001",
			1514 => "0001000011111000000100",
			1515 => "0000000001011110110101",
			1516 => "0000000001011110110101",
			1517 => "0000101011111000001000",
			1518 => "0000010000111100000100",
			1519 => "0000000001011111001001",
			1520 => "0000000001011111001001",
			1521 => "0000000001011111001001",
			1522 => "0001000000010100000100",
			1523 => "0000000001011111011101",
			1524 => "0001001010010000000100",
			1525 => "0000000001011111011101",
			1526 => "0000000001011111011101",
			1527 => "0000100110101100000100",
			1528 => "0000000001011111110001",
			1529 => "0000101101101100000100",
			1530 => "0000000001011111110001",
			1531 => "0000000001011111110001",
			1532 => "0001000010100100000100",
			1533 => "0000000001100000000101",
			1534 => "0001001010010000000100",
			1535 => "0000000001100000000101",
			1536 => "0000000001100000000101",
			1537 => "0000101011111000000100",
			1538 => "0000000001100000011001",
			1539 => "0000101100111000000100",
			1540 => "0000000001100000011001",
			1541 => "0000000001100000011001",
			1542 => "0000100110101100000100",
			1543 => "0000000001100000101101",
			1544 => "0000101111101000000100",
			1545 => "0000000001100000101101",
			1546 => "0000000001100000101101",
			1547 => "0000011101011100001000",
			1548 => "0001000100111000000100",
			1549 => "0000000001100001000001",
			1550 => "0000000001100001000001",
			1551 => "0000000001100001000001",
			1552 => "0001000011111000001100",
			1553 => "0000011101011100001000",
			1554 => "0010011101011000000100",
			1555 => "0000000001100001011101",
			1556 => "0000000001100001011101",
			1557 => "0000000001100001011101",
			1558 => "0000000001100001011101",
			1559 => "0001000101100000001100",
			1560 => "0000011101011100001000",
			1561 => "0010011101011000000100",
			1562 => "0000000001100001111001",
			1563 => "0000000001100001111001",
			1564 => "0000000001100001111001",
			1565 => "0000000001100001111001",
			1566 => "0001000010100100000100",
			1567 => "0000000001100010010101",
			1568 => "0000100000010000000100",
			1569 => "0000000001100010010101",
			1570 => "0000101111101000000100",
			1571 => "0000000001100010010101",
			1572 => "0000000001100010010101",
			1573 => "0010011101011000001100",
			1574 => "0001000100111000001000",
			1575 => "0000011101011100000100",
			1576 => "0000000001100010110001",
			1577 => "0000000001100010110001",
			1578 => "0000000001100010110001",
			1579 => "0000000001100010110001",
			1580 => "0010011010011000001000",
			1581 => "0001000100111000000100",
			1582 => "0000000001100011010101",
			1583 => "0000000001100011010101",
			1584 => "0011101001010100001000",
			1585 => "0001010100010000000100",
			1586 => "0000000001100011010101",
			1587 => "0000000001100011010101",
			1588 => "0000000001100011010101",
			1589 => "0000011111001100000100",
			1590 => "0000000001100011111001",
			1591 => "0001111101010100001100",
			1592 => "0011101110101000001000",
			1593 => "0011000000001100000100",
			1594 => "0000000001100011111001",
			1595 => "0000000001100011111001",
			1596 => "0000000001100011111001",
			1597 => "0000000001100011111001",
			1598 => "0001000011010100000100",
			1599 => "0000000001100100011101",
			1600 => "0000100110101100000100",
			1601 => "0000000001100100011101",
			1602 => "0000100011000000001000",
			1603 => "0001001010010000000100",
			1604 => "0000000001100100011101",
			1605 => "0000000001100100011101",
			1606 => "0000000001100100011101",
			1607 => "0001000010100100000100",
			1608 => "0000000001100101000001",
			1609 => "0000101100111000001100",
			1610 => "0000100000010000000100",
			1611 => "0000000001100101000001",
			1612 => "0001001010010000000100",
			1613 => "0000000001100101000001",
			1614 => "0000000001100101000001",
			1615 => "0000000001100101000001",
			1616 => "0010011010011000001000",
			1617 => "0001000100111000000100",
			1618 => "0000000001100101101101",
			1619 => "0000000001100101101101",
			1620 => "0011101110101000001100",
			1621 => "0000101011111000000100",
			1622 => "0000000001100101101101",
			1623 => "0011000100001000000100",
			1624 => "0000000001100101101101",
			1625 => "0000000001100101101101",
			1626 => "0000000001100101101101",
			1627 => "0000011111001100001000",
			1628 => "0001000100111000000100",
			1629 => "0000000001100110011001",
			1630 => "0000000001100110011001",
			1631 => "0011100111110000001100",
			1632 => "0001111101111000000100",
			1633 => "0000000001100110011001",
			1634 => "0001101001100100000100",
			1635 => "0000000001100110011001",
			1636 => "0000000001100110011001",
			1637 => "0000000001100110011001",
			1638 => "0001000011110100000100",
			1639 => "0000000001100111000101",
			1640 => "0010110011100000001000",
			1641 => "0000011111001100000100",
			1642 => "0000000001100111000101",
			1643 => "0000000001100111000101",
			1644 => "0010001011010100000100",
			1645 => "0000000001100111000101",
			1646 => "0011110011001000000100",
			1647 => "0000000001100111000101",
			1648 => "0000000001100111000101",
			1649 => "0000100110101100010000",
			1650 => "0000000011111100000100",
			1651 => "0000000001101000000001",
			1652 => "0001101001100100001000",
			1653 => "0011000000001100000100",
			1654 => "0000000001101000000001",
			1655 => "0000000001101000000001",
			1656 => "0000000001101000000001",
			1657 => "0011111100010000001100",
			1658 => "0010100001110000001000",
			1659 => "0001111110001100000100",
			1660 => "0000000001101000000001",
			1661 => "0000000001101000000001",
			1662 => "0000000001101000000001",
			1663 => "0000000001101000000001",
			1664 => "0000101011111000001000",
			1665 => "0010001011010100000100",
			1666 => "0000000001101000110101",
			1667 => "0000000001101000110101",
			1668 => "0011111100000000010000",
			1669 => "0001110110000100000100",
			1670 => "0000000001101000110101",
			1671 => "0010101100000100001000",
			1672 => "0000100110101100000100",
			1673 => "0000000001101000110101",
			1674 => "0000000001101000110101",
			1675 => "0000000001101000110101",
			1676 => "0000000001101000110101",
			1677 => "0000011101101000000100",
			1678 => "0000000001101001100001",
			1679 => "0011101110101100010000",
			1680 => "0011000100001000001100",
			1681 => "0011111111010000000100",
			1682 => "0000000001101001100001",
			1683 => "0011000110000100000100",
			1684 => "0000000001101001100001",
			1685 => "0000000001101001100001",
			1686 => "0000000001101001100001",
			1687 => "0000000001101001100001",
			1688 => "0000101000001100001100",
			1689 => "0001111100101000001000",
			1690 => "0011001110001100000100",
			1691 => "1111111001101010100101",
			1692 => "0000000001101010100101",
			1693 => "0000000001101010100101",
			1694 => "0011110011001000001100",
			1695 => "0010001010101100001000",
			1696 => "0000011011101000000100",
			1697 => "0000000001101010100101",
			1698 => "0000000001101010100101",
			1699 => "0000000001101010100101",
			1700 => "0011101110101100001000",
			1701 => "0000011101011100000100",
			1702 => "0000000001101010100101",
			1703 => "0000000001101010100101",
			1704 => "0000000001101010100101",
			1705 => "0000100111011000000100",
			1706 => "1111111001101011100001",
			1707 => "0001101011001100001100",
			1708 => "0000010110101000000100",
			1709 => "0000000001101011100001",
			1710 => "0011101110101100000100",
			1711 => "0000000001101011100001",
			1712 => "0000000001101011100001",
			1713 => "0010011010011000000100",
			1714 => "0000000001101011100001",
			1715 => "0011101001010100000100",
			1716 => "0000000001101011100001",
			1717 => "0001101011001100000100",
			1718 => "0000000001101011100001",
			1719 => "0000000001101011100001",
			1720 => "0000101011111000001100",
			1721 => "0010001011010100000100",
			1722 => "0000000001101100100101",
			1723 => "0011000000001100000100",
			1724 => "0000000001101100100101",
			1725 => "0000000001101100100101",
			1726 => "0011111100000000010100",
			1727 => "0011000110000100000100",
			1728 => "0000000001101100100101",
			1729 => "0011000100001000001100",
			1730 => "0001101001100100001000",
			1731 => "0000010110101000000100",
			1732 => "0000000001101100100101",
			1733 => "0000000001101100100101",
			1734 => "0000000001101100100101",
			1735 => "0000000001101100100101",
			1736 => "0000000001101100100101",
			1737 => "0001001011100000000100",
			1738 => "1111111001101101101001",
			1739 => "0000100110101100010000",
			1740 => "0010001011010100001100",
			1741 => "0011110010000000001000",
			1742 => "0000011111001100000100",
			1743 => "0000000001101101101001",
			1744 => "0000000001101101101001",
			1745 => "0000000001101101101001",
			1746 => "0000000001101101101001",
			1747 => "0001100100111100001100",
			1748 => "0010101100000100001000",
			1749 => "0000010110101000000100",
			1750 => "0000000001101101101001",
			1751 => "0000000001101101101001",
			1752 => "0000000001101101101001",
			1753 => "0000000001101101101001",
			1754 => "0000101000001100001100",
			1755 => "0011001110001100001000",
			1756 => "0001111100101000000100",
			1757 => "1111111001101110110101",
			1758 => "0000000001101110110101",
			1759 => "0000000001101110110101",
			1760 => "0011111100000000011000",
			1761 => "0000011111001100010000",
			1762 => "0001101101011000001100",
			1763 => "0001001111101100001000",
			1764 => "0001000011111000000100",
			1765 => "0000000001101110110101",
			1766 => "0000000001101110110101",
			1767 => "0000000001101110110101",
			1768 => "0000000001101110110101",
			1769 => "0000101011111000000100",
			1770 => "0000000001101110110101",
			1771 => "0000000001101110110101",
			1772 => "0000000001101110110101",
			1773 => "0001001001000000001000",
			1774 => "0010011010011000000100",
			1775 => "1111111001110000010001",
			1776 => "0000000001110000010001",
			1777 => "0000100110101100010000",
			1778 => "0010001011010100001100",
			1779 => "0011110010000000001000",
			1780 => "0011110101110000000100",
			1781 => "0000000001110000010001",
			1782 => "0000000001110000010001",
			1783 => "0000000001110000010001",
			1784 => "0000000001110000010001",
			1785 => "0011000110000100001100",
			1786 => "0000011101011100001000",
			1787 => "0000011101101000000100",
			1788 => "0000000001110000010001",
			1789 => "0000000001110000010001",
			1790 => "0000000001110000010001",
			1791 => "0011110111011000001000",
			1792 => "0010101100000100000100",
			1793 => "0000000001110000010001",
			1794 => "0000000001110000010001",
			1795 => "0000000001110000010001",
			1796 => "0000010110101000000100",
			1797 => "0000000001110001011101",
			1798 => "0000111101000100010100",
			1799 => "0011000100001000010000",
			1800 => "0001110110000100000100",
			1801 => "0000000001110001011101",
			1802 => "0001000000010100000100",
			1803 => "0000000001110001011101",
			1804 => "0010101100000100000100",
			1805 => "0000000001110001011101",
			1806 => "0000000001110001011101",
			1807 => "0000000001110001011101",
			1808 => "0010011111000000001000",
			1809 => "0011010101110100000100",
			1810 => "0000000001110001011101",
			1811 => "0000000001110001011101",
			1812 => "0010110110100100000100",
			1813 => "0000000001110001011101",
			1814 => "0000000001110001011101",
			1815 => "0000100000010000001100",
			1816 => "0010011111000000001000",
			1817 => "0011001110001100000100",
			1818 => "1111111001110010110001",
			1819 => "0000000001110010110001",
			1820 => "0000000001110010110001",
			1821 => "0011110010000100011000",
			1822 => "0000100110101100000100",
			1823 => "0000000001110010110001",
			1824 => "0011001100110000000100",
			1825 => "0000000001110010110001",
			1826 => "0010101100000100001100",
			1827 => "0011101001010100001000",
			1828 => "0001101001100100000100",
			1829 => "0000001001110010110001",
			1830 => "0000000001110010110001",
			1831 => "0000000001110010110001",
			1832 => "0000000001110010110001",
			1833 => "0011111100000000000100",
			1834 => "0000000001110010110001",
			1835 => "0000000001110010110001",
			1836 => "0010110011100000011100",
			1837 => "0011000011011100000100",
			1838 => "0000000001110011111101",
			1839 => "0011111001100000010100",
			1840 => "0000100111011000000100",
			1841 => "0000000001110011111101",
			1842 => "0001001010010000001100",
			1843 => "0011011000011000000100",
			1844 => "0000000001110011111101",
			1845 => "0000101000101000000100",
			1846 => "0000000001110011111101",
			1847 => "0000000001110011111101",
			1848 => "0000000001110011111101",
			1849 => "0000000001110011111101",
			1850 => "0011110011001000000100",
			1851 => "0000000001110011111101",
			1852 => "0011010101110100000100",
			1853 => "0000000001110011111101",
			1854 => "0000000001110011111101",
			1855 => "0000010110101000000100",
			1856 => "0000000001110101000001",
			1857 => "0011111100010000011100",
			1858 => "0010000110001000001000",
			1859 => "0001001110111000000100",
			1860 => "0000000001110101000001",
			1861 => "0000000001110101000001",
			1862 => "0001000100111000001100",
			1863 => "0010111000000000001000",
			1864 => "0000101100111000000100",
			1865 => "0000000001110101000001",
			1866 => "0000000001110101000001",
			1867 => "0000000001110101000001",
			1868 => "0010111010111100000100",
			1869 => "0000000001110101000001",
			1870 => "0000000001110101000001",
			1871 => "0000000001110101000001",
			1872 => "0000100000010000010100",
			1873 => "0000011111001100000100",
			1874 => "1111111001110110101101",
			1875 => "0010110011100000001100",
			1876 => "0000100000010000001000",
			1877 => "0011000011011100000100",
			1878 => "0000000001110110101101",
			1879 => "0000000001110110101101",
			1880 => "0000000001110110101101",
			1881 => "1111111001110110101101",
			1882 => "0001101011001100010000",
			1883 => "0000010110101000000100",
			1884 => "0000000001110110101101",
			1885 => "0000110011001000001000",
			1886 => "0011000110000100000100",
			1887 => "0000000001110110101101",
			1888 => "0000001001110110101101",
			1889 => "0000000001110110101101",
			1890 => "0000111001011100010000",
			1891 => "0010011010011000000100",
			1892 => "0000000001110110101101",
			1893 => "0000101011111000001000",
			1894 => "0011010101110100000100",
			1895 => "0000000001110110101101",
			1896 => "0000000001110110101101",
			1897 => "0000001001110110101101",
			1898 => "1111111001110110101101",
			1899 => "0001110110000100001000",
			1900 => "0011000110000100000100",
			1901 => "0000000001111000001001",
			1902 => "0000000001111000001001",
			1903 => "0000111101000100011000",
			1904 => "0011000100001000010100",
			1905 => "0010011101011100000100",
			1906 => "0000000001111000001001",
			1907 => "0001000000010100000100",
			1908 => "0000000001111000001001",
			1909 => "0000001100101100001000",
			1910 => "0000101000101000000100",
			1911 => "0000000001111000001001",
			1912 => "0000000001111000001001",
			1913 => "0000000001111000001001",
			1914 => "0000000001111000001001",
			1915 => "0010110011100000000100",
			1916 => "0000000001111000001001",
			1917 => "0001101001100100001000",
			1918 => "0010010100111100000100",
			1919 => "0000000001111000001001",
			1920 => "0000000001111000001001",
			1921 => "0000000001111000001001",
			1922 => "0001000011110100000100",
			1923 => "1111111001111001100101",
			1924 => "0000011111001100001100",
			1925 => "0000011101101000000100",
			1926 => "1111111001111001100101",
			1927 => "0001101011001100000100",
			1928 => "0000001001111001100101",
			1929 => "1111111001111001100101",
			1930 => "0011101001010100010000",
			1931 => "0000001110111100000100",
			1932 => "0000001001111001100101",
			1933 => "0000101011101100000100",
			1934 => "0000000001111001100101",
			1935 => "0000100001011100000100",
			1936 => "0000001001111001100101",
			1937 => "0000000001111001100101",
			1938 => "0010001011010100000100",
			1939 => "0000001001111001100101",
			1940 => "0000010000111100000100",
			1941 => "1111111001111001100101",
			1942 => "0000010101011100000100",
			1943 => "0000000001111001100101",
			1944 => "0000000001111001100101",
			1945 => "0001000010100100001000",
			1946 => "0001000011110100000100",
			1947 => "1111111001111011100001",
			1948 => "0000000001111011100001",
			1949 => "0000100110101100011100",
			1950 => "0010001011010100001100",
			1951 => "0000011111001100000100",
			1952 => "0000000001111011100001",
			1953 => "0011111100010100000100",
			1954 => "0000000001111011100001",
			1955 => "0000000001111011100001",
			1956 => "0001101001100100001100",
			1957 => "0010111000000000001000",
			1958 => "0010100110011000000100",
			1959 => "0000000001111011100001",
			1960 => "1111111001111011100001",
			1961 => "0000000001111011100001",
			1962 => "0000000001111011100001",
			1963 => "0011010001011000001100",
			1964 => "0010101100000100001000",
			1965 => "0011001100110000000100",
			1966 => "0000000001111011100001",
			1967 => "0000001001111011100001",
			1968 => "0000000001111011100001",
			1969 => "0000011101011100001000",
			1970 => "0011100100010000000100",
			1971 => "0000000001111011100001",
			1972 => "0000000001111011100001",
			1973 => "0011011110101100000100",
			1974 => "0000000001111011100001",
			1975 => "0000000001111011100001",
			1976 => "0001000010100100000100",
			1977 => "1111111001111100111101",
			1978 => "0011101001010100011100",
			1979 => "0000011111001100011000",
			1980 => "0001000100111000001000",
			1981 => "0011001110001100000100",
			1982 => "0000000001111100111101",
			1983 => "0000000001111100111101",
			1984 => "0010101100000100001100",
			1985 => "0011011010001100001000",
			1986 => "0011110111110000000100",
			1987 => "0000000001111100111101",
			1988 => "0000000001111100111101",
			1989 => "0000000001111100111101",
			1990 => "0000000001111100111101",
			1991 => "0000000001111100111101",
			1992 => "0011001110001100001000",
			1993 => "0011001100110000000100",
			1994 => "0000000001111100111101",
			1995 => "0000000001111100111101",
			1996 => "0011110111011000000100",
			1997 => "0000000001111100111101",
			1998 => "0000000001111100111101",
			1999 => "0000101111010100001100",
			2000 => "0000100111011000000100",
			2001 => "1111111001111111001001",
			2002 => "0000100110111100000100",
			2003 => "0000000001111111001001",
			2004 => "0000000001111111001001",
			2005 => "0011000100001000101100",
			2006 => "0000100110101100011000",
			2007 => "0010001011010100001100",
			2008 => "0011101110101100001000",
			2009 => "0011001100110000000100",
			2010 => "0000000001111111001001",
			2011 => "0000001001111111001001",
			2012 => "0000000001111111001001",
			2013 => "0011001110001100001000",
			2014 => "0000101011111000000100",
			2015 => "1111111001111111001001",
			2016 => "0000000001111111001001",
			2017 => "0000000001111111001001",
			2018 => "0011001100110000001000",
			2019 => "0010101010110000000100",
			2020 => "0000000001111111001001",
			2021 => "0000000001111111001001",
			2022 => "0010100001110000001000",
			2023 => "0000111001011100000100",
			2024 => "0000001001111111001001",
			2025 => "0000000001111111001001",
			2026 => "0000000001111111001001",
			2027 => "0001111110110000001100",
			2028 => "0010111000000000000100",
			2029 => "0000000001111111001001",
			2030 => "0011101001010000000100",
			2031 => "0000000001111111001001",
			2032 => "0000000001111111001001",
			2033 => "1111111001111111001001",
			2034 => "0010011010011000101000",
			2035 => "0000011101011100100100",
			2036 => "0000011111001100011000",
			2037 => "0000101011111000000100",
			2038 => "1111111010000001000101",
			2039 => "0000100110101100001000",
			2040 => "0000010110000000000100",
			2041 => "0000000010000001000101",
			2042 => "0000110010000001000101",
			2043 => "0010111010111100001000",
			2044 => "0011000110000100000100",
			2045 => "1111111010000001000101",
			2046 => "0001100010000001000101",
			2047 => "1111111010000001000101",
			2048 => "0011010101100100001000",
			2049 => "0000000010011000000100",
			2050 => "0000000010000001000101",
			2051 => "0000100010000001000101",
			2052 => "1111111010000001000101",
			2053 => "1111110010000001000101",
			2054 => "0011101110101000010100",
			2055 => "0010010100111100010000",
			2056 => "0011100111110000001000",
			2057 => "0000011101011100000100",
			2058 => "0000001010000001000101",
			2059 => "0000001010000001000101",
			2060 => "0001011011011100000100",
			2061 => "0000001010000001000101",
			2062 => "1111111010000001000101",
			2063 => "0000011010000001000101",
			2064 => "1111111010000001000101",
			2065 => "0000011101101000000100",
			2066 => "1111111010000010111001",
			2067 => "0011000100001000101100",
			2068 => "0011101001010100011100",
			2069 => "0011010010001000001100",
			2070 => "0011111001010000000100",
			2071 => "0000000010000010111001",
			2072 => "0010110001111100000100",
			2073 => "0000000010000010111001",
			2074 => "0000001010000010111001",
			2075 => "0001000010010000001000",
			2076 => "0000001000110000000100",
			2077 => "0000000010000010111001",
			2078 => "0000001010000010111001",
			2079 => "0011110010000000000100",
			2080 => "1111111010000010111001",
			2081 => "0000000010000010111001",
			2082 => "0011001110001100001000",
			2083 => "0010100110011000000100",
			2084 => "0000000010000010111001",
			2085 => "1111111010000010111001",
			2086 => "0011101110101000000100",
			2087 => "0000001010000010111001",
			2088 => "0000000010000010111001",
			2089 => "0001010100010000000100",
			2090 => "0000000010000010111001",
			2091 => "0011000100001000000100",
			2092 => "0000000010000010111001",
			2093 => "1111111010000010111001",
			2094 => "0000101111010100001100",
			2095 => "0000100111011000000100",
			2096 => "1111111010000100110101",
			2097 => "0000100110111100000100",
			2098 => "0000000010000100110101",
			2099 => "0000000010000100110101",
			2100 => "0011001010111100101100",
			2101 => "0011101001010100010100",
			2102 => "0010011110010100000100",
			2103 => "1111111010000100110101",
			2104 => "0010100001010100001100",
			2105 => "0011000100001000001000",
			2106 => "0000000100000000000100",
			2107 => "0000001010000100110101",
			2108 => "0000001010000100110101",
			2109 => "0000000010000100110101",
			2110 => "0000000010000100110101",
			2111 => "0010001011010100001000",
			2112 => "0001001110111000000100",
			2113 => "1111111010000100110101",
			2114 => "0000001010000100110101",
			2115 => "0000100110101100000100",
			2116 => "1111111010000100110101",
			2117 => "0000011001011000000100",
			2118 => "1111111010000100110101",
			2119 => "0010011000010000000100",
			2120 => "0000000010000100110101",
			2121 => "0000000010000100110101",
			2122 => "0001110111001000000100",
			2123 => "0000000010000100110101",
			2124 => "1111111010000100110101",
			2125 => "0000101111010100000100",
			2126 => "1111111010000110101001",
			2127 => "0011000100001000100100",
			2128 => "0000011101101000001100",
			2129 => "0011000110000100000100",
			2130 => "1111111010000110101001",
			2131 => "0001111101111000000100",
			2132 => "0000011010000110101001",
			2133 => "1111111010000110101001",
			2134 => "0011101000011000000100",
			2135 => "0000110010000110101001",
			2136 => "0010000001110100001100",
			2137 => "0011101110101000001000",
			2138 => "0011101110101100000100",
			2139 => "0000001010000110101001",
			2140 => "0000011010000110101001",
			2141 => "1111111010000110101001",
			2142 => "0001101111000000000100",
			2143 => "1111110010000110101001",
			2144 => "1111111010000110101001",
			2145 => "0001110111001000010000",
			2146 => "0010111000000000001000",
			2147 => "0001110111001000000100",
			2148 => "1111111010000110101001",
			2149 => "0000000010000110101001",
			2150 => "0000110111100000000100",
			2151 => "0000001010000110101001",
			2152 => "0000000010000110101001",
			2153 => "1111111010000110101001",
			2154 => "0000101111010100001000",
			2155 => "0000100111011000000100",
			2156 => "1111111010001000010101",
			2157 => "1111111010001000010101",
			2158 => "0011101110101000101100",
			2159 => "0000011101101000001100",
			2160 => "0000010110101000000100",
			2161 => "1111111010001000010101",
			2162 => "0000010110101000000100",
			2163 => "0000100010001000010101",
			2164 => "1111111010001000010101",
			2165 => "0011100001101000001000",
			2166 => "0010001000110000000100",
			2167 => "0000101010001000010101",
			2168 => "0000001010001000010101",
			2169 => "0010000001110100010000",
			2170 => "0000011111001100001000",
			2171 => "0011110010000000000100",
			2172 => "0000010010001000010101",
			2173 => "0000000010001000010101",
			2174 => "0000011101011100000100",
			2175 => "0000000010001000010101",
			2176 => "0000001010001000010101",
			2177 => "0001101001100100000100",
			2178 => "0000000010001000010101",
			2179 => "1111111010001000010101",
			2180 => "1111111010001000010101",
			2181 => "0000101111010100001000",
			2182 => "0000101111010100000100",
			2183 => "1111111010001010001001",
			2184 => "0000000010001010001001",
			2185 => "0011101100101100001000",
			2186 => "0000111011000000000100",
			2187 => "0000000010001010001001",
			2188 => "0001001010001010001001",
			2189 => "0001101011001100001100",
			2190 => "0010111001001000001000",
			2191 => "0000011101101000000100",
			2192 => "0000000010001010001001",
			2193 => "0000001010001010001001",
			2194 => "0000000010001010001001",
			2195 => "0011101110101000011100",
			2196 => "0000011101011100010000",
			2197 => "0000101111100100001000",
			2198 => "0000000011010000000100",
			2199 => "0000000010001010001001",
			2200 => "1111111010001010001001",
			2201 => "0010011010011000000100",
			2202 => "0000000010001010001001",
			2203 => "0000000010001010001001",
			2204 => "0000101011111000001000",
			2205 => "0000111101000100000100",
			2206 => "0000000010001010001001",
			2207 => "0000000010001010001001",
			2208 => "0000001010001010001001",
			2209 => "1111111010001010001001",
			2210 => "0000100110111100001100",
			2211 => "0000100111011000000100",
			2212 => "1111111010001100011101",
			2213 => "0000100110111100000100",
			2214 => "0000000010001100011101",
			2215 => "1111111010001100011101",
			2216 => "0011000100001000110000",
			2217 => "0010011011111100000100",
			2218 => "1111111010001100011101",
			2219 => "0011101001010100010000",
			2220 => "0011101011000000000100",
			2221 => "0000011010001100011101",
			2222 => "0010001010101100001000",
			2223 => "0001010101100100000100",
			2224 => "0000001010001100011101",
			2225 => "0000000010001100011101",
			2226 => "1111111010001100011101",
			2227 => "0010001011010100001100",
			2228 => "0011101110101000001000",
			2229 => "0011001110001100000100",
			2230 => "0000000010001100011101",
			2231 => "0000001010001100011101",
			2232 => "1111111010001100011101",
			2233 => "0000101000100000001000",
			2234 => "0001011010011100000100",
			2235 => "0000000010001100011101",
			2236 => "1111110010001100011101",
			2237 => "0011111111010100000100",
			2238 => "0000000010001100011101",
			2239 => "0000000010001100011101",
			2240 => "0001110111001000001100",
			2241 => "0010111000000000000100",
			2242 => "1111111010001100011101",
			2243 => "0000110111100000000100",
			2244 => "0000001010001100011101",
			2245 => "0000000010001100011101",
			2246 => "1111111010001100011101",
			2247 => "0000101111010100000100",
			2248 => "1111111010001110101011",
			2249 => "0011000100001000110100",
			2250 => "0000011101101000000100",
			2251 => "1111111010001110101011",
			2252 => "0011101001010100011000",
			2253 => "0000011111001100001100",
			2254 => "0010001000101100001000",
			2255 => "0010110111001000000100",
			2256 => "0000011010001110101011",
			2257 => "0000010010001110101011",
			2258 => "0000000010001110101011",
			2259 => "0000011101011100001000",
			2260 => "0011010010001000000100",
			2261 => "0000001010001110101011",
			2262 => "1111111010001110101011",
			2263 => "0000001010001110101011",
			2264 => "0000011001011000001100",
			2265 => "0001001101110100001000",
			2266 => "0001000000010100000100",
			2267 => "1111111010001110101011",
			2268 => "0000000010001110101011",
			2269 => "1111101010001110101011",
			2270 => "0011101110101000001000",
			2271 => "0000100110101100000100",
			2272 => "0000000010001110101011",
			2273 => "0000010010001110101011",
			2274 => "1111111010001110101011",
			2275 => "0001110111001000001100",
			2276 => "0011100111110000001000",
			2277 => "0001010100000100000100",
			2278 => "0000000010001110101011",
			2279 => "0000001010001110101011",
			2280 => "1111111010001110101011",
			2281 => "1111111010001110101011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(726, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(1470, initial_addr_3'length));
	end generate gen_rom_12;

	gen_rom_13: if SELECT_ROM = 13 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0001001110111000000100",
			11 => "0000000000000000110101",
			12 => "0000000000000000110101",
			13 => "0000011011101000000100",
			14 => "0000000000000001001001",
			15 => "0000010000111100000100",
			16 => "0000000000000001001001",
			17 => "0000000000000001001001",
			18 => "0011000110000100001000",
			19 => "0011000000101000000100",
			20 => "0000000000000001011101",
			21 => "0000000000000001011101",
			22 => "0000000000000001011101",
			23 => "0010011101101000000100",
			24 => "0000000000000001110001",
			25 => "0010010100111100000100",
			26 => "0000000000000001110001",
			27 => "0000000000000001110001",
			28 => "0000110111100000001000",
			29 => "0001001101000000000100",
			30 => "0000000000000010000101",
			31 => "0000000000000010000101",
			32 => "0000000000000010000101",
			33 => "0011110110010000001000",
			34 => "0011110010001000000100",
			35 => "0000000000000010100001",
			36 => "0000000000000010100001",
			37 => "0011111011110000000100",
			38 => "0000000000000010100001",
			39 => "0000000000000010100001",
			40 => "0001101011001100001000",
			41 => "0000000010111100000100",
			42 => "0000000000000010111101",
			43 => "0000000000000010111101",
			44 => "0001101000010000000100",
			45 => "0000000000000010111101",
			46 => "0000000000000010111101",
			47 => "0000100100101000000100",
			48 => "0000000000000011011001",
			49 => "0001000001100100001000",
			50 => "0011111011110000000100",
			51 => "0000000000000011011001",
			52 => "0000000000000011011001",
			53 => "0000000000000011011001",
			54 => "0001011011011100001100",
			55 => "0000000010111100000100",
			56 => "0000000000000011110101",
			57 => "0000001010111100000100",
			58 => "0000000000000011110101",
			59 => "0000000000000011110101",
			60 => "0000000000000011110101",
			61 => "0011011011110100001100",
			62 => "0000000010111100000100",
			63 => "0000000000000100010001",
			64 => "0000001010111100000100",
			65 => "0000000000000100010001",
			66 => "0000000000000100010001",
			67 => "0000000000000100010001",
			68 => "0000001110111100000100",
			69 => "0000000000000100101101",
			70 => "0000011100110100000100",
			71 => "0000000000000100101101",
			72 => "0000011101011100000100",
			73 => "0000000000000100101101",
			74 => "0000000000000100101101",
			75 => "0000110010001000001000",
			76 => "0001101001100100000100",
			77 => "0000000000000101010001",
			78 => "0000000000000101010001",
			79 => "0010010100111100001000",
			80 => "0010010001000100000100",
			81 => "0000000000000101010001",
			82 => "0000000000000101010001",
			83 => "0000000000000101010001",
			84 => "0001101011001100001000",
			85 => "0000100100101000000100",
			86 => "0000000000000101111101",
			87 => "0000000000000101111101",
			88 => "0001001100111100001000",
			89 => "0001001000000100000100",
			90 => "0000000000000101111101",
			91 => "0000000000000101111101",
			92 => "0001000100100100000100",
			93 => "0000000000000101111101",
			94 => "0000000000000101111101",
			95 => "0011000011011100001100",
			96 => "0001111001110000000100",
			97 => "0000000000000110101001",
			98 => "0011010100011000000100",
			99 => "0000000000000110101001",
			100 => "0000000000000110101001",
			101 => "0011011001010100001000",
			102 => "0001110110000100000100",
			103 => "0000000000000110101001",
			104 => "0000000000000110101001",
			105 => "0000000000000110101001",
			106 => "0001111100101000010000",
			107 => "0001111001110000000100",
			108 => "0000000000000111001101",
			109 => "0011001100110000001000",
			110 => "0011000000101000000100",
			111 => "0000000000000111001101",
			112 => "0000000000000111001101",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0001011011011100010000",
			116 => "0001001000000100000100",
			117 => "0000000000000111110001",
			118 => "0001001010010000001000",
			119 => "0000100100101000000100",
			120 => "0000000000000111110001",
			121 => "0000000000000111110001",
			122 => "0000000000000111110001",
			123 => "0000000000000111110001",
			124 => "0001011011011100000100",
			125 => "0000000000001000010101",
			126 => "0010010101010000001100",
			127 => "0010010001111000000100",
			128 => "0000000000001000010101",
			129 => "0011010111111100000100",
			130 => "0000000000001000010101",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0000001110111100000100",
			134 => "0000000000001000111001",
			135 => "0000011100110100000100",
			136 => "0000000000001000111001",
			137 => "0000011101011100001000",
			138 => "0010001101010000000100",
			139 => "0000000000001000111001",
			140 => "0000000000001000111001",
			141 => "0000000000001000111001",
			142 => "0000100100101000000100",
			143 => "0000000000001001100101",
			144 => "0011011011110100001000",
			145 => "0000001010111100000100",
			146 => "0000000000001001100101",
			147 => "0000000000001001100101",
			148 => "0001110100011000000100",
			149 => "0000000000001001100101",
			150 => "0001110111010000000100",
			151 => "0000000000001001100101",
			152 => "0000000000001001100101",
			153 => "0000001110111100001100",
			154 => "0000000010111100000100",
			155 => "0000000000001010011001",
			156 => "0001000000100000000100",
			157 => "0000000000001010011001",
			158 => "0000000000001010011001",
			159 => "0010000001110100001100",
			160 => "0001111001110000000100",
			161 => "0000000000001010011001",
			162 => "0001111101010100000100",
			163 => "0000000000001010011001",
			164 => "0000000000001010011001",
			165 => "0000000000001010011001",
			166 => "0000000011111100001100",
			167 => "0010100110011000000100",
			168 => "0000000000001011001101",
			169 => "0010100001010000000100",
			170 => "0000000000001011001101",
			171 => "0000000000001011001101",
			172 => "0011111000101000001100",
			173 => "0010100110011000000100",
			174 => "0000000000001011001101",
			175 => "0000001010111100000100",
			176 => "0000000000001011001101",
			177 => "0000000000001011001101",
			178 => "0000000000001011001101",
			179 => "0010100001010000001100",
			180 => "0010100110011000000100",
			181 => "0000000000001100000001",
			182 => "0011001001110000000100",
			183 => "0000000000001100000001",
			184 => "0000000000001100000001",
			185 => "0010110110100100001100",
			186 => "0011001000111100000100",
			187 => "0000000000001100000001",
			188 => "0001001010010000000100",
			189 => "0000000000001100000001",
			190 => "0000000000001100000001",
			191 => "0000000000001100000001",
			192 => "0000110010001000001000",
			193 => "0001101001100100000100",
			194 => "0000000000001100110101",
			195 => "0000000000001100110101",
			196 => "0001100101010000010000",
			197 => "0000010101011100001100",
			198 => "0010010001000100000100",
			199 => "0000000000001100110101",
			200 => "0001101011001100000100",
			201 => "0000000000001100110101",
			202 => "0000000000001100110101",
			203 => "0000000000001100110101",
			204 => "0000000000001100110101",
			205 => "0001000100001100001100",
			206 => "0001001000000100000100",
			207 => "0000000000001101110001",
			208 => "0001101000010000000100",
			209 => "0000000000001101110001",
			210 => "0000000000001101110001",
			211 => "0001101111000000010000",
			212 => "0000011100110100000100",
			213 => "0000000000001101110001",
			214 => "0000011101011100001000",
			215 => "0001000100111000000100",
			216 => "0000000000001101110001",
			217 => "0000000000001101110001",
			218 => "0000000000001101110001",
			219 => "0000000000001101110001",
			220 => "0001011011011100001100",
			221 => "0001001000000100000100",
			222 => "0000000000001110101101",
			223 => "0001000101001100000100",
			224 => "0000000000001110101101",
			225 => "0000000000001110101101",
			226 => "0011001010111000010000",
			227 => "0000010101011100001100",
			228 => "0011100100010000000100",
			229 => "0000000000001110101101",
			230 => "0010100110011000000100",
			231 => "0000000000001110101101",
			232 => "0000000000001110101101",
			233 => "0000000000001110101101",
			234 => "0000000000001110101101",
			235 => "0001110111001000011100",
			236 => "0010110100011000010000",
			237 => "0001001000000100000100",
			238 => "0000000000001111111001",
			239 => "0001001101000000001000",
			240 => "0000111000000000000100",
			241 => "0000000000001111111001",
			242 => "0000000000001111111001",
			243 => "0000000000001111111001",
			244 => "0011010100010000000100",
			245 => "0000000000001111111001",
			246 => "0001001001000000000100",
			247 => "0000000000001111111001",
			248 => "0000000000001111111001",
			249 => "0000110011000000001000",
			250 => "0011000000001100000100",
			251 => "0000000000001111111001",
			252 => "0000000000001111111001",
			253 => "0000000000001111111001",
			254 => "0011110000010000011100",
			255 => "0011010100010000001000",
			256 => "0011100010001000000100",
			257 => "0000000000010000111101",
			258 => "0000000000010000111101",
			259 => "0010110100011000000100",
			260 => "0000000000010000111101",
			261 => "0011000100001000001100",
			262 => "0000010101011100001000",
			263 => "0011100011001000000100",
			264 => "0000000000010000111101",
			265 => "0000000000010000111101",
			266 => "0000000000010000111101",
			267 => "0000000000010000111101",
			268 => "0000000010011000000100",
			269 => "0000000000010000111101",
			270 => "0000000000010000111101",
			271 => "0000000010111100010100",
			272 => "0000000010011000000100",
			273 => "0000000000010010001001",
			274 => "0001011000000000000100",
			275 => "0000000000010010001001",
			276 => "0010001011010100001000",
			277 => "0001000010100100000100",
			278 => "0000000000010010001001",
			279 => "0000000000010010001001",
			280 => "0000000000010010001001",
			281 => "0011111010010100000100",
			282 => "0000000000010010001001",
			283 => "0001000001100100001100",
			284 => "0000101010001000000100",
			285 => "0000000000010010001001",
			286 => "0011101010000100000100",
			287 => "0000000000010010001001",
			288 => "0000000000010010001001",
			289 => "0000000000010010001001",
			290 => "0011011001010100011000",
			291 => "0000101010001000000100",
			292 => "0000000000010010111101",
			293 => "0000001010111100010000",
			294 => "0000011001011000001100",
			295 => "0000001000111100001000",
			296 => "0000110111100000000100",
			297 => "0000000000010010111101",
			298 => "0000000000010010111101",
			299 => "0000000000010010111101",
			300 => "0000000000010010111101",
			301 => "0000000000010010111101",
			302 => "0000000000010010111101",
			303 => "0000000010111100011000",
			304 => "0010001001101000000100",
			305 => "0000000000010100001001",
			306 => "0010011001111100010000",
			307 => "0011011001110100000100",
			308 => "0000000000010100001001",
			309 => "0010001011010100001000",
			310 => "0001001000000100000100",
			311 => "0000000000010100001001",
			312 => "0000000000010100001001",
			313 => "0000000000010100001001",
			314 => "0000000000010100001001",
			315 => "0010011110010100001100",
			316 => "0001001010010000001000",
			317 => "0011110010110100000100",
			318 => "0000000000010100001001",
			319 => "0000000000010100001001",
			320 => "0000000000010100001001",
			321 => "0000000000010100001001",
			322 => "0010010100110100100000",
			323 => "0000101110010000010100",
			324 => "0000110011100000000100",
			325 => "0000000000010101011101",
			326 => "0010111110001100001100",
			327 => "0010110101101100000100",
			328 => "0000000000010101011101",
			329 => "0000111010011100000100",
			330 => "0000000000010101011101",
			331 => "0000000000010101011101",
			332 => "0000000000010101011101",
			333 => "0001001010010000001000",
			334 => "0011110111110000000100",
			335 => "0000000000010101011101",
			336 => "0000000000010101011101",
			337 => "0000000000010101011101",
			338 => "0000011001011000001000",
			339 => "0010011010011000000100",
			340 => "0000000000010101011101",
			341 => "0000000000010101011101",
			342 => "0000000000010101011101",
			343 => "0011000011011100011000",
			344 => "0010110101101100000100",
			345 => "0000000000010110110001",
			346 => "0010001001101000000100",
			347 => "0000000000010110110001",
			348 => "0000100110010000001100",
			349 => "0001111001110000000100",
			350 => "0000000000010110110001",
			351 => "0011010100011000000100",
			352 => "0000000000010110110001",
			353 => "0000000000010110110001",
			354 => "0000000000010110110001",
			355 => "0011110101110000000100",
			356 => "0000000000010110110001",
			357 => "0000110011000000001100",
			358 => "0000100110101100000100",
			359 => "0000000000010110110001",
			360 => "0001111100101000000100",
			361 => "0000000000010110110001",
			362 => "0000000000010110110001",
			363 => "0000000000010110110001",
			364 => "0011001100110000011100",
			365 => "0011000100000000000100",
			366 => "0000000000010111111101",
			367 => "0000000010111100000100",
			368 => "0000000000010111111101",
			369 => "0011100101101100000100",
			370 => "0000000000010111111101",
			371 => "0001100100110100000100",
			372 => "0000000000010111111101",
			373 => "0000100010010100001000",
			374 => "0000111001011100000100",
			375 => "0000000000010111111101",
			376 => "0000000000010111111101",
			377 => "0000000000010111111101",
			378 => "0000100011000000001000",
			379 => "0000100110101100000100",
			380 => "0000000000010111111101",
			381 => "0000000000010111111101",
			382 => "0000000000010111111101",
			383 => "0011110110010000011100",
			384 => "0001111001110000000100",
			385 => "0000000000011001000001",
			386 => "0011001110001100010100",
			387 => "0000101011101100010000",
			388 => "0001101001100100001100",
			389 => "0001100100110100000100",
			390 => "0000000000011001000001",
			391 => "0011111011011100000100",
			392 => "0000000000011001000001",
			393 => "0000000000011001000001",
			394 => "0000000000011001000001",
			395 => "0000000000011001000001",
			396 => "0000000000011001000001",
			397 => "0011000011011100000100",
			398 => "0000000000011001000001",
			399 => "0000000000011001000001",
			400 => "0010010111101000001000",
			401 => "0000001010111100000100",
			402 => "0000000000011010000101",
			403 => "0000000000011010000101",
			404 => "0001110100011000011000",
			405 => "0011010101110100000100",
			406 => "0000000000011010000101",
			407 => "0010010100111100010000",
			408 => "0000011011101000000100",
			409 => "0000000000011010000101",
			410 => "0011110011001000000100",
			411 => "0000000000011010000101",
			412 => "0010100110011000000100",
			413 => "0000000000011010000101",
			414 => "0000000000011010000101",
			415 => "0000000000011010000101",
			416 => "0000000000011010000101",
			417 => "0010010001000100001000",
			418 => "0001000011111000000100",
			419 => "0000000000011011011001",
			420 => "0000000000011011011001",
			421 => "0000011111001100011000",
			422 => "0001101011001100000100",
			423 => "0000000000011011011001",
			424 => "0000111001011100010000",
			425 => "0011000011011100000100",
			426 => "0000000000011011011001",
			427 => "0000000010111100000100",
			428 => "0000000000011011011001",
			429 => "0010001111000100000100",
			430 => "0000000000011011011001",
			431 => "0000000000011011011001",
			432 => "0000000000011011011001",
			433 => "0011110010000000000100",
			434 => "0000000000011011011001",
			435 => "0001100100111100000100",
			436 => "0000000000011011011001",
			437 => "0000000000011011011001",
			438 => "0011001100110000011100",
			439 => "0011010100011000000100",
			440 => "0000000000011100101101",
			441 => "0010001001101000000100",
			442 => "0000000000011100101101",
			443 => "0011110110010000010000",
			444 => "0001101111000000001100",
			445 => "0000000010111100000100",
			446 => "0000000000011100101101",
			447 => "0011000000101000000100",
			448 => "0000000000011100101101",
			449 => "0000000000011100101101",
			450 => "0000000000011100101101",
			451 => "0000000000011100101101",
			452 => "0000101011111000000100",
			453 => "0000000000011100101101",
			454 => "0000000010111100000100",
			455 => "0000000000011100101101",
			456 => "0000001010111100000100",
			457 => "0000000000011100101101",
			458 => "0000000000011100101101",
			459 => "0011000011011100011100",
			460 => "0011000100000000000100",
			461 => "0000000000011110000001",
			462 => "0010001001101000000100",
			463 => "0000000000011110000001",
			464 => "0000100110010000010000",
			465 => "0010011101101000000100",
			466 => "0000000000011110000001",
			467 => "0011010100011000000100",
			468 => "0000000000011110000001",
			469 => "0001111001110000000100",
			470 => "0000000000011110000001",
			471 => "0000000000011110000001",
			472 => "0000000000011110000001",
			473 => "0011110101110000000100",
			474 => "0000000000011110000001",
			475 => "0000000010111100000100",
			476 => "0000000000011110000001",
			477 => "0001110110000100000100",
			478 => "0000000000011110000001",
			479 => "0000000000011110000001",
			480 => "0010011101101000000100",
			481 => "0000000000011110111101",
			482 => "0000010101011100011000",
			483 => "0010110101101100000100",
			484 => "0000000000011110111101",
			485 => "0010001001101000000100",
			486 => "0000000000011110111101",
			487 => "0001101000010000001100",
			488 => "0001111110110000001000",
			489 => "0000000010011000000100",
			490 => "0000000000011110111101",
			491 => "0000000000011110111101",
			492 => "0000000000011110111101",
			493 => "0000000000011110111101",
			494 => "0000000000011110111101",
			495 => "0011101100101100000100",
			496 => "0000000000011111111001",
			497 => "0011001110001100011000",
			498 => "0010100110011000000100",
			499 => "0000000000011111111001",
			500 => "0010011101101000000100",
			501 => "0000000000011111111001",
			502 => "0011000100000000000100",
			503 => "0000000000011111111001",
			504 => "0010010100111100001000",
			505 => "0011101001011100000100",
			506 => "0000000000011111111001",
			507 => "0000000000011111111001",
			508 => "0000000000011111111001",
			509 => "0000000000011111111001",
			510 => "0001010000011100011000",
			511 => "0000101110010000010000",
			512 => "0000111010111100000100",
			513 => "0000000000100001011101",
			514 => "0000100101001000000100",
			515 => "0000000000100001011101",
			516 => "0011110010110100000100",
			517 => "0000000000100001011101",
			518 => "0000000000100001011101",
			519 => "0000001000111100000100",
			520 => "0000000000100001011101",
			521 => "0000000000100001011101",
			522 => "0000010000111100011000",
			523 => "0011001100110000000100",
			524 => "0000000000100001011101",
			525 => "0000101100001100010000",
			526 => "0000001111000100000100",
			527 => "0000000000100001011101",
			528 => "0010011011111100000100",
			529 => "0000000000100001011101",
			530 => "0011010010001000000100",
			531 => "0000000000100001011101",
			532 => "0000000000100001011101",
			533 => "0000000000100001011101",
			534 => "0000000000100001011101",
			535 => "0000011011101000011100",
			536 => "0011110100101000011000",
			537 => "0011101100101100000100",
			538 => "0000000000100010111001",
			539 => "0001111001110000000100",
			540 => "0000000000100010111001",
			541 => "0011000110000100001100",
			542 => "0010110101101100000100",
			543 => "0000000000100010111001",
			544 => "0011000100000000000100",
			545 => "0000000000100010111001",
			546 => "0000000000100010111001",
			547 => "0000000000100010111001",
			548 => "0000000000100010111001",
			549 => "0000011101011100010000",
			550 => "0000000000110000000100",
			551 => "0000000000100010111001",
			552 => "0001110001101000001000",
			553 => "0010101010110000000100",
			554 => "0000000000100010111001",
			555 => "0000000000100010111001",
			556 => "0000000000100010111001",
			557 => "0000000000100010111001",
			558 => "0000100110101100011100",
			559 => "0010110101101100000100",
			560 => "0000000000100100010101",
			561 => "0011001110001100010100",
			562 => "0000000010111100000100",
			563 => "0000000000100100010101",
			564 => "0010001001101000000100",
			565 => "0000000000100100010101",
			566 => "0011000100000000000100",
			567 => "0000000000100100010101",
			568 => "0001111001110000000100",
			569 => "0000000000100100010101",
			570 => "0000000000100100010101",
			571 => "0000000000100100010101",
			572 => "0000000010111100000100",
			573 => "0000000000100100010101",
			574 => "0011001100110000000100",
			575 => "0000000000100100010101",
			576 => "0001110110000100000100",
			577 => "0000000000100100010101",
			578 => "0000001010111100000100",
			579 => "0000000000100100010101",
			580 => "0000000000100100010101",
			581 => "0001111100101000101100",
			582 => "0000010110101000010100",
			583 => "0001000011101100000100",
			584 => "0000000000100110001001",
			585 => "0011100000001100001100",
			586 => "0001111001110000000100",
			587 => "0000000000100110001001",
			588 => "0000111110001100000100",
			589 => "0000000000100110001001",
			590 => "0000000000100110001001",
			591 => "0000000000100110001001",
			592 => "0001101000010000010100",
			593 => "0001101101011000000100",
			594 => "0000000000100110001001",
			595 => "0011000011011100000100",
			596 => "0000000000100110001001",
			597 => "0000000010111100000100",
			598 => "0000000000100110001001",
			599 => "0010100110011000000100",
			600 => "0000000000100110001001",
			601 => "0000000000100110001001",
			602 => "0000000000100110001001",
			603 => "0000110111100000001100",
			604 => "0010111110110000000100",
			605 => "0000000000100110001001",
			606 => "0000100000010000000100",
			607 => "0000000000100110001001",
			608 => "0000000000100110001001",
			609 => "0000000000100110001001",
			610 => "0001000011010100011000",
			611 => "0011110000110100010000",
			612 => "0011101101111000000100",
			613 => "0000000000101000011101",
			614 => "0010110101101100000100",
			615 => "0000000000101000011101",
			616 => "0010111100101100000100",
			617 => "0000000000101000011101",
			618 => "0000000000101000011101",
			619 => "0001010101110000000100",
			620 => "0000000000101000011101",
			621 => "0000000000101000011101",
			622 => "0010000111000100010100",
			623 => "0010010100111100010000",
			624 => "0010100110011000000100",
			625 => "0000000000101000011101",
			626 => "0000000111111000001000",
			627 => "0000011100110100000100",
			628 => "0000000000101000011101",
			629 => "0000000000101000011101",
			630 => "0000000000101000011101",
			631 => "0000000000101000011101",
			632 => "0001100100111100011000",
			633 => "0011010001011000001100",
			634 => "0001000101001100001000",
			635 => "0000111110110000000100",
			636 => "0000000000101000011101",
			637 => "0000000000101000011101",
			638 => "0000000000101000011101",
			639 => "0001000110110000000100",
			640 => "0000000000101000011101",
			641 => "0000010110101000000100",
			642 => "0000000000101000011101",
			643 => "0000000000101000011101",
			644 => "0011011100100100000100",
			645 => "0000000000101000011101",
			646 => "0000000000101000011101",
			647 => "0011010100011000000100",
			648 => "0000000000101001111001",
			649 => "0001111100101000011000",
			650 => "0000000010111100000100",
			651 => "0000000000101001111001",
			652 => "0000111001011100010000",
			653 => "0010011101101000000100",
			654 => "0000000000101001111001",
			655 => "0010110101101100000100",
			656 => "0000000000101001111001",
			657 => "0011001110001100000100",
			658 => "0000000000101001111001",
			659 => "0000000000101001111001",
			660 => "0000000000101001111001",
			661 => "0000100110101100000100",
			662 => "0000000000101001111001",
			663 => "0000011111001100000100",
			664 => "0000000000101001111001",
			665 => "0000000010111100000100",
			666 => "0000000000101001111001",
			667 => "0000001000111000000100",
			668 => "0000000000101001111001",
			669 => "0000000000101001111001",
			670 => "0011011011000000001000",
			671 => "0001001101000000000100",
			672 => "1111111000101011110101",
			673 => "0000000000101011110101",
			674 => "0000100110010000010100",
			675 => "0001111101100000010000",
			676 => "0011001000111000000100",
			677 => "0000000000101011110101",
			678 => "0010111110001100001000",
			679 => "0000000010111100000100",
			680 => "0000000000101011110101",
			681 => "0000001000101011110101",
			682 => "0000000000101011110101",
			683 => "0000000000101011110101",
			684 => "0000011011101000010000",
			685 => "0001000011111000001000",
			686 => "0011100011100000000100",
			687 => "0000000000101011110101",
			688 => "0000000000101011110101",
			689 => "0001101011001100000100",
			690 => "0000000000101011110101",
			691 => "0000000000101011110101",
			692 => "0010100110011000000100",
			693 => "0000000000101011110101",
			694 => "0000111111101000001100",
			695 => "0010111110110000000100",
			696 => "0000000000101011110101",
			697 => "0000010101011100000100",
			698 => "0000000000101011110101",
			699 => "0000000000101011110101",
			700 => "0000000000101011110101",
			701 => "0011010100011000000100",
			702 => "1111111000101101010001",
			703 => "0011000100001000011100",
			704 => "0010100111000100011000",
			705 => "0000000010011000000100",
			706 => "1111111000101101010001",
			707 => "0000101001011100000100",
			708 => "0000010000101101010001",
			709 => "0001010011100000001000",
			710 => "0000110011100000000100",
			711 => "0000000000101101010001",
			712 => "1111111000101101010001",
			713 => "0001101101011000000100",
			714 => "0000000000101101010001",
			715 => "0000001000101101010001",
			716 => "1111111000101101010001",
			717 => "0000100101000000000100",
			718 => "1111111000101101010001",
			719 => "0011110101000000001000",
			720 => "0001000011101100000100",
			721 => "0000001000101101010001",
			722 => "0000000000101101010001",
			723 => "1111111000101101010001",
			724 => "0001001001000000100100",
			725 => "0001000011010100001100",
			726 => "0000100101000000000100",
			727 => "1111111000101111110101",
			728 => "0000100101000000000100",
			729 => "0000000000101111110101",
			730 => "1111111000101111110101",
			731 => "0010000110001000010100",
			732 => "0010001001101000001100",
			733 => "0001000011110100001000",
			734 => "0001001111100000000100",
			735 => "0000000000101111110101",
			736 => "0000001000101111110101",
			737 => "1111111000101111110101",
			738 => "0010101010110000000100",
			739 => "0000010000101111110101",
			740 => "0000000000101111110101",
			741 => "1111111000101111110101",
			742 => "0000010010001100001100",
			743 => "0000101000101000001000",
			744 => "0000100001011100000100",
			745 => "1111111000101111110101",
			746 => "1111110000101111110101",
			747 => "0000000000101111110101",
			748 => "0000101011110000011000",
			749 => "0000101110110100000100",
			750 => "0000011000101111110101",
			751 => "0011101001010100001100",
			752 => "0000011101011100001000",
			753 => "0001010100011000000100",
			754 => "1111111000101111110101",
			755 => "0000001000101111110101",
			756 => "1111111000101111110101",
			757 => "0000011001011000000100",
			758 => "0000011000101111110101",
			759 => "0000001000101111110101",
			760 => "0010000001110100001000",
			761 => "0010100110011100000100",
			762 => "0000000000101111110101",
			763 => "0000000000101111110101",
			764 => "1111111000101111110101",
			765 => "0011110110010000110100",
			766 => "0001111001110000001000",
			767 => "0010100110001000000100",
			768 => "0000000000110001101001",
			769 => "0000000000110001101001",
			770 => "0001111101100000010100",
			771 => "0000100110010000010000",
			772 => "0011101001110000000100",
			773 => "0000000000110001101001",
			774 => "0010100110011000000100",
			775 => "0000000000110001101001",
			776 => "0011010100011000000100",
			777 => "0000000000110001101001",
			778 => "0000001000110001101001",
			779 => "0000000000110001101001",
			780 => "0001001011001000001000",
			781 => "0000101010001000000100",
			782 => "0000000000110001101001",
			783 => "0000000000110001101001",
			784 => "0011101010111000000100",
			785 => "0000000000110001101001",
			786 => "0001110111001000001000",
			787 => "0010001011010100000100",
			788 => "0000000000110001101001",
			789 => "0000000000110001101001",
			790 => "0000000000110001101001",
			791 => "0011100111111100000100",
			792 => "0000000000110001101001",
			793 => "0000000000110001101001",
			794 => "0001001001000000011000",
			795 => "0001000100001100000100",
			796 => "1111111000110011011101",
			797 => "0010000111000100010000",
			798 => "0001000100001100000100",
			799 => "0000011000110011011101",
			800 => "0000111001011100000100",
			801 => "1111111000110011011101",
			802 => "0001110111010000000100",
			803 => "0000001000110011011101",
			804 => "1111111000110011011101",
			805 => "1111111000110011011101",
			806 => "0000011100110100000100",
			807 => "1111111000110011011101",
			808 => "0001101000010000011100",
			809 => "0000100110010000000100",
			810 => "0000010000110011011101",
			811 => "0001101101011000001000",
			812 => "0011111100100100000100",
			813 => "0000001000110011011101",
			814 => "1111110000110011011101",
			815 => "0011011011000000001000",
			816 => "0000111010111000000100",
			817 => "0000000000110011011101",
			818 => "1111111000110011011101",
			819 => "0010001011010100000100",
			820 => "0000000000110011011101",
			821 => "0000001000110011011101",
			822 => "1111111000110011011101",
			823 => "0000100100101000010000",
			824 => "0011101001110000000100",
			825 => "0000000000110101111001",
			826 => "0001000010111000000100",
			827 => "0000000000110101111001",
			828 => "0010111101100000000100",
			829 => "0000000000110101111001",
			830 => "0000000000110101111001",
			831 => "0000000010111100011000",
			832 => "0010100110011000000100",
			833 => "0000000000110101111001",
			834 => "0000010101011100010000",
			835 => "0010010001000100000100",
			836 => "0000000000110101111001",
			837 => "0010001011010100001000",
			838 => "0001001011110000000100",
			839 => "0000000000110101111001",
			840 => "0000000000110101111001",
			841 => "0000000000110101111001",
			842 => "0000000000110101111001",
			843 => "0001001101110100001100",
			844 => "0010011111000000001000",
			845 => "0000100111111100000100",
			846 => "0000000000110101111001",
			847 => "0000000000110101111001",
			848 => "0000000000110101111001",
			849 => "0001101111000000010000",
			850 => "0011101011000100000100",
			851 => "0000000000110101111001",
			852 => "0010111110110000001000",
			853 => "0001101111000000000100",
			854 => "0000000000110101111001",
			855 => "0000000000110101111001",
			856 => "0000000000110101111001",
			857 => "0011101001100000001000",
			858 => "0000110110100000000100",
			859 => "0000000000110101111001",
			860 => "0000000000110101111001",
			861 => "0000000000110101111001",
			862 => "0001001001000000011100",
			863 => "0001000000010100000100",
			864 => "1111111000110111101101",
			865 => "0010110101101100000100",
			866 => "1111111000110111101101",
			867 => "0010101010110000010000",
			868 => "0000010101011100001100",
			869 => "0010100110011000001000",
			870 => "0001000011110100000100",
			871 => "0000000000110111101101",
			872 => "0000000000110111101101",
			873 => "0000001000110111101101",
			874 => "1111111000110111101101",
			875 => "1111111000110111101101",
			876 => "0000011100110100000100",
			877 => "1111111000110111101101",
			878 => "0001101000010000011000",
			879 => "0001110011100000010100",
			880 => "0010011101101000000100",
			881 => "0000100000110111101101",
			882 => "0001010100011000001000",
			883 => "0000110111001000000100",
			884 => "0000000000110111101101",
			885 => "1111111000110111101101",
			886 => "0010001011010100000100",
			887 => "0000000000110111101101",
			888 => "0000001000110111101101",
			889 => "1111111000110111101101",
			890 => "1111111000110111101101",
			891 => "0001101000010000110000",
			892 => "0011010100011000000100",
			893 => "0000000000111001010001",
			894 => "0000100110010000010100",
			895 => "0001011001110100010000",
			896 => "0010100110011000000100",
			897 => "0000000000111001010001",
			898 => "0011101001110000000100",
			899 => "0000000000111001010001",
			900 => "0000000010111100000100",
			901 => "0000000000111001010001",
			902 => "0000000000111001010001",
			903 => "0000000000111001010001",
			904 => "0001001011001000001000",
			905 => "0011010110100000000100",
			906 => "0000000000111001010001",
			907 => "0000000000111001010001",
			908 => "0000010110101000000100",
			909 => "0000000000111001010001",
			910 => "0010111001110100001000",
			911 => "0010111010111100000100",
			912 => "0000000000111001010001",
			913 => "0000000000111001010001",
			914 => "0000000000111001010001",
			915 => "0000000000111001010001",
			916 => "0001001001000000100100",
			917 => "0001000000010100000100",
			918 => "1111111000111011111101",
			919 => "0000000010111100001100",
			920 => "0000010101011100001000",
			921 => "0010100110011000000100",
			922 => "1111111000111011111101",
			923 => "0000110000111011111101",
			924 => "1111111000111011111101",
			925 => "0010110101101100000100",
			926 => "1111111000111011111101",
			927 => "0001101010011000000100",
			928 => "0000010000111011111101",
			929 => "0010101010110000001000",
			930 => "0000011001011000000100",
			931 => "0000100000111011111101",
			932 => "1111111000111011111101",
			933 => "1111111000111011111101",
			934 => "0010011011101000001000",
			935 => "0000010010001100000100",
			936 => "1111111000111011111101",
			937 => "0000000000111011111101",
			938 => "0001100100111100100000",
			939 => "0011100111110000010000",
			940 => "0010011010011000001100",
			941 => "0000000100010100000100",
			942 => "0000011000111011111101",
			943 => "0011111100010100000100",
			944 => "0000001000111011111101",
			945 => "0000010000111011111101",
			946 => "1111111000111011111101",
			947 => "0001011011011100001000",
			948 => "0011001110001100000100",
			949 => "0000001000111011111101",
			950 => "0000000000111011111101",
			951 => "0001111010111100000100",
			952 => "0010000000111011111101",
			953 => "0000101000111011111101",
			954 => "0010100101000100000100",
			955 => "0000000000111011111101",
			956 => "0011011001110100000100",
			957 => "1111110000111011111101",
			958 => "1111111000111011111101",
			959 => "0010011101101000000100",
			960 => "0000000000111101110001",
			961 => "0011000011011100011000",
			962 => "0010110101101100000100",
			963 => "0000000000111101110001",
			964 => "0000000010111100000100",
			965 => "0000000000111101110001",
			966 => "0001101000010000001100",
			967 => "0011000100000000000100",
			968 => "0000000000111101110001",
			969 => "0001111001110000000100",
			970 => "0000000000111101110001",
			971 => "0000001000111101110001",
			972 => "0000000000111101110001",
			973 => "0000100011110000011100",
			974 => "0010110100011000001100",
			975 => "0001001101000000001000",
			976 => "0011100000001100000100",
			977 => "0000000000111101110001",
			978 => "0000000000111101110001",
			979 => "0000000000111101110001",
			980 => "0000010000111100001100",
			981 => "0000011011101000000100",
			982 => "0000000000111101110001",
			983 => "0001000000010100000100",
			984 => "0000000000111101110001",
			985 => "0000000000111101110001",
			986 => "0000000000111101110001",
			987 => "0000000000111101110001",
			988 => "0011010100011000000100",
			989 => "1111111000111111010101",
			990 => "0010001001101000000100",
			991 => "1111111000111111010101",
			992 => "0000101110010000001000",
			993 => "0010111110001100000100",
			994 => "0000001000111111010101",
			995 => "0000000000111111010101",
			996 => "0001101000010000011000",
			997 => "0010111110001100001000",
			998 => "0000110100011000000100",
			999 => "0000000000111111010101",
			1000 => "1111111000111111010101",
			1001 => "0001101011001100001000",
			1002 => "0001000101100000000100",
			1003 => "0000000000111111010101",
			1004 => "1111111000111111010101",
			1005 => "0000011001011000000100",
			1006 => "0000001000111111010101",
			1007 => "0000000000111111010101",
			1008 => "0010100001010000001000",
			1009 => "0000011110010100000100",
			1010 => "0000000000111111010101",
			1011 => "0000000000111111010101",
			1012 => "1111111000111111010101",
			1013 => "0011010100011000000100",
			1014 => "1111111001000001011001",
			1015 => "0011111101000100010000",
			1016 => "0011111011011100000100",
			1017 => "0000000001000001011001",
			1018 => "0001000010111000000100",
			1019 => "0000000001000001011001",
			1020 => "0011000110000100000100",
			1021 => "0000001001000001011001",
			1022 => "0000000001000001011001",
			1023 => "0010010100110100010100",
			1024 => "0001001101000000001000",
			1025 => "0011000110000100000100",
			1026 => "1111111001000001011001",
			1027 => "0000000001000001011001",
			1028 => "0011000110000100000100",
			1029 => "0000000001000001011001",
			1030 => "0001000100111000000100",
			1031 => "0000000001000001011001",
			1032 => "1111111001000001011001",
			1033 => "0001000011010100000100",
			1034 => "0000000001000001011001",
			1035 => "0010100110011100010000",
			1036 => "0011100100010000001000",
			1037 => "0010011010011000000100",
			1038 => "0000000001000001011001",
			1039 => "0000000001000001011001",
			1040 => "0001111010111100000100",
			1041 => "0000001001000001011001",
			1042 => "0000000001000001011001",
			1043 => "0011011001010100000100",
			1044 => "0000000001000001011001",
			1045 => "0000000001000001011001",
			1046 => "0010100110011000000100",
			1047 => "0000000001000011001101",
			1048 => "0010001011010100010000",
			1049 => "0000010101011100001100",
			1050 => "0011000011011100000100",
			1051 => "0000000001000011001101",
			1052 => "0001000111011100000100",
			1053 => "0000001001000011001101",
			1054 => "0000000001000011001101",
			1055 => "0000000001000011001101",
			1056 => "0001000100001100000100",
			1057 => "0000000001000011001101",
			1058 => "0000101110010000001000",
			1059 => "0000111010111100000100",
			1060 => "0000000001000011001101",
			1061 => "0000001001000011001101",
			1062 => "0000010110101000001100",
			1063 => "0010000010111100001000",
			1064 => "0011110111110000000100",
			1065 => "0000000001000011001101",
			1066 => "0000000001000011001101",
			1067 => "0000000001000011001101",
			1068 => "0001101011001100001000",
			1069 => "0010111010111100000100",
			1070 => "0000000001000011001101",
			1071 => "0000000001000011001101",
			1072 => "0001001101000000000100",
			1073 => "0000000001000011001101",
			1074 => "0000000001000011001101",
			1075 => "0001001001000000101100",
			1076 => "0010110101101100000100",
			1077 => "1111111001000101110001",
			1078 => "0011010110100100010100",
			1079 => "0001011000000000001000",
			1080 => "0000010010001100000100",
			1081 => "0000001001000101110001",
			1082 => "1111111001000101110001",
			1083 => "0000100110010000001000",
			1084 => "0000000010111100000100",
			1085 => "0000000001000101110001",
			1086 => "0000100001000101110001",
			1087 => "0000000001000101110001",
			1088 => "0001000000010100000100",
			1089 => "1111111001000101110001",
			1090 => "0000000010011000001100",
			1091 => "0010100110011000000100",
			1092 => "0000000001000101110001",
			1093 => "0000010111101000000100",
			1094 => "0000001001000101110001",
			1095 => "0000000001000101110001",
			1096 => "1111111001000101110001",
			1097 => "0000011100110100000100",
			1098 => "1111111001000101110001",
			1099 => "0001110111001000011100",
			1100 => "0011110111110000000100",
			1101 => "0000010001000101110001",
			1102 => "0010111110001100001000",
			1103 => "0000000100001000000100",
			1104 => "1111111001000101110001",
			1105 => "0000001001000101110001",
			1106 => "0011001100110000001000",
			1107 => "0000000100010100000100",
			1108 => "0000010001000101110001",
			1109 => "0000001001000101110001",
			1110 => "0001101101011000000100",
			1111 => "1111111001000101110001",
			1112 => "0000001001000101110001",
			1113 => "0011000100001000000100",
			1114 => "0000000001000101110001",
			1115 => "1111111001000101110001",
			1116 => "0010011111001100000100",
			1117 => "1111111001000111110101",
			1118 => "0010100110011100100000",
			1119 => "0000001111000100000100",
			1120 => "1111111001000111110101",
			1121 => "0011001000111000000100",
			1122 => "0000000001000111110101",
			1123 => "0011000011011100001100",
			1124 => "0010100001010000000100",
			1125 => "0000001001000111110101",
			1126 => "0000001010000000000100",
			1127 => "0000000001000111110101",
			1128 => "0000001001000111110101",
			1129 => "0011010010001000000100",
			1130 => "0000000001000111110101",
			1131 => "0010010101010000000100",
			1132 => "0000000001000111110101",
			1133 => "0000000001000111110101",
			1134 => "0000001100101100011000",
			1135 => "0011001110001100010000",
			1136 => "0011001100110000001100",
			1137 => "0001110101101100000100",
			1138 => "0000000001000111110101",
			1139 => "0011111100010000000100",
			1140 => "0000000001000111110101",
			1141 => "0000000001000111110101",
			1142 => "1111111001000111110101",
			1143 => "0011000100001000000100",
			1144 => "0000000001000111110101",
			1145 => "0000000001000111110101",
			1146 => "0000111010110100000100",
			1147 => "0000000001000111110101",
			1148 => "0000000001000111110101",
			1149 => "0010100110011000000100",
			1150 => "0000000001001001110001",
			1151 => "0010001011010100010000",
			1152 => "0000010101011100001100",
			1153 => "0011000011011100000100",
			1154 => "0000000001001001110001",
			1155 => "0001000111011100000100",
			1156 => "0000001001001001110001",
			1157 => "0000000001001001110001",
			1158 => "0000000001001001110001",
			1159 => "0001000100001100000100",
			1160 => "0000000001001001110001",
			1161 => "0000101110010000001000",
			1162 => "0000111010111100000100",
			1163 => "0000000001001001110001",
			1164 => "0000001001001001110001",
			1165 => "0001101011001100010000",
			1166 => "0011100100011000001000",
			1167 => "0011001100110000000100",
			1168 => "0000000001001001110001",
			1169 => "0000000001001001110001",
			1170 => "0010111010111100000100",
			1171 => "0000000001001001110001",
			1172 => "0000000001001001110001",
			1173 => "0001001101000000001000",
			1174 => "0001000011101100000100",
			1175 => "0000000001001001110001",
			1176 => "0000000001001001110001",
			1177 => "0010101111001000000100",
			1178 => "0000000001001001110001",
			1179 => "0000000001001001110001",
			1180 => "0010110101101100000100",
			1181 => "1111111001001011100101",
			1182 => "0001000010111000000100",
			1183 => "1111111001001011100101",
			1184 => "0010000111000100010100",
			1185 => "0000010101011100010000",
			1186 => "0000100011001000000100",
			1187 => "0000001001001011100101",
			1188 => "0001010101100100000100",
			1189 => "0000000001001011100101",
			1190 => "0010100110011000000100",
			1191 => "0000000001001011100101",
			1192 => "0000001001001011100101",
			1193 => "0000000001001011100101",
			1194 => "0011000110000100010000",
			1195 => "0001000001100100000100",
			1196 => "1111111001001011100101",
			1197 => "0000100010010100001000",
			1198 => "0011001100110000000100",
			1199 => "0000001001001011100101",
			1200 => "0000000001001011100101",
			1201 => "0000000001001011100101",
			1202 => "0001101011001100000100",
			1203 => "1111111001001011100101",
			1204 => "0001000110110000000100",
			1205 => "0000000001001011100101",
			1206 => "0011000100001000000100",
			1207 => "0000000001001011100101",
			1208 => "0000000001001011100101",
			1209 => "0011010100011000000100",
			1210 => "1111111001001110000001",
			1211 => "0001101100011000010000",
			1212 => "0011010110100100001100",
			1213 => "0001000010111000000100",
			1214 => "0000000001001110000001",
			1215 => "0011110001011000000100",
			1216 => "0000000001001110000001",
			1217 => "0000001001001110000001",
			1218 => "0000000001001110000001",
			1219 => "0001010000011100010100",
			1220 => "0001001101000000001000",
			1221 => "0011111110101100000100",
			1222 => "0000000001001110000001",
			1223 => "1111111001001110000001",
			1224 => "0011000110000100001000",
			1225 => "0011100000101000000100",
			1226 => "0000000001001110000001",
			1227 => "0000000001001110000001",
			1228 => "0000000001001110000001",
			1229 => "0001110001111100010000",
			1230 => "0000011111001100000100",
			1231 => "0000000001001110000001",
			1232 => "0010001011010100000100",
			1233 => "0000000001001110000001",
			1234 => "0000110110010000000100",
			1235 => "0000000001001110000001",
			1236 => "0000000001001110000001",
			1237 => "0000011001011000001100",
			1238 => "0001101001100100000100",
			1239 => "0000000001001110000001",
			1240 => "0010101100000100000100",
			1241 => "0000000001001110000001",
			1242 => "0000000001001110000001",
			1243 => "0011111110100100001000",
			1244 => "0001101011001100000100",
			1245 => "0000000001001110000001",
			1246 => "0000000001001110000001",
			1247 => "0000000001001110000001",
			1248 => "0001111001110000001000",
			1249 => "0000101000100000000100",
			1250 => "1111111001010000100101",
			1251 => "0000000001010000100101",
			1252 => "0001111001110000001100",
			1253 => "0000100110010000001000",
			1254 => "0011010100011000000100",
			1255 => "0000000001010000100101",
			1256 => "0000001001010000100101",
			1257 => "0000000001010000100101",
			1258 => "0010000111000100010100",
			1259 => "0001000010111000000100",
			1260 => "0000000001010000100101",
			1261 => "0000010101011100001100",
			1262 => "0000011001111000000100",
			1263 => "0000000001010000100101",
			1264 => "0011011011000000000100",
			1265 => "0000000001010000100101",
			1266 => "0000000001010000100101",
			1267 => "0000000001010000100101",
			1268 => "0011110101110000010100",
			1269 => "0001101101011000001100",
			1270 => "0001000100111000000100",
			1271 => "0000000001010000100101",
			1272 => "0001011000000000000100",
			1273 => "0000000001010000100101",
			1274 => "0000000001010000100101",
			1275 => "0000101111010100000100",
			1276 => "0000000001010000100101",
			1277 => "0000000001010000100101",
			1278 => "0000011011101000001000",
			1279 => "0000110100000100000100",
			1280 => "0000000001010000100101",
			1281 => "1111111001010000100101",
			1282 => "0000011111001100001000",
			1283 => "0000101011110000000100",
			1284 => "0000000001010000100101",
			1285 => "0000000001010000100101",
			1286 => "0000011111001100000100",
			1287 => "0000000001010000100101",
			1288 => "0000000001010000100101",
			1289 => "0001001001000000110000",
			1290 => "0010110101101100000100",
			1291 => "1111111001010011100001",
			1292 => "0011010110100100011000",
			1293 => "0011011001110100001000",
			1294 => "0010011011101000000100",
			1295 => "0000001001010011100001",
			1296 => "1111111001010011100001",
			1297 => "0011001000111000000100",
			1298 => "0000000001010011100001",
			1299 => "0010111110001100001000",
			1300 => "0001101011001100000100",
			1301 => "0000011001010011100001",
			1302 => "0000000001010011100001",
			1303 => "0000000001010011100001",
			1304 => "0001000000010100000100",
			1305 => "1111111001010011100001",
			1306 => "0000000010011000001100",
			1307 => "0010100110011000000100",
			1308 => "0000000001010011100001",
			1309 => "0010010100101100000100",
			1310 => "0000001001010011100001",
			1311 => "0000000001010011100001",
			1312 => "1111111001010011100001",
			1313 => "0000011100110100000100",
			1314 => "1111111001010011100001",
			1315 => "0001110111001000100000",
			1316 => "0001101010011000000100",
			1317 => "0000010001010011100001",
			1318 => "0010111110001100001100",
			1319 => "0000111000000000001000",
			1320 => "0011010100011000000100",
			1321 => "0000000001010011100001",
			1322 => "0000001001010011100001",
			1323 => "1111111001010011100001",
			1324 => "0011001100110000001000",
			1325 => "0000000100010100000100",
			1326 => "0000010001010011100001",
			1327 => "0000001001010011100001",
			1328 => "0001101101011000000100",
			1329 => "1111111001010011100001",
			1330 => "0000001001010011100001",
			1331 => "0010100001110000001000",
			1332 => "0001000110110000000100",
			1333 => "1111111001010011100001",
			1334 => "0000000001010011100001",
			1335 => "1111111001010011100001",
			1336 => "0011010100011000000100",
			1337 => "1111111001010110011101",
			1338 => "0000100110010000100100",
			1339 => "0001111101100000010000",
			1340 => "0000000010111100000100",
			1341 => "0000000001010110011101",
			1342 => "0010101010110000001000",
			1343 => "0001111001110000000100",
			1344 => "0000000001010110011101",
			1345 => "0000001001010110011101",
			1346 => "0000000001010110011101",
			1347 => "0001000011010100000100",
			1348 => "0000000001010110011101",
			1349 => "0001010011100000000100",
			1350 => "0000000001010110011101",
			1351 => "0001011001110100001000",
			1352 => "0001111101111000000100",
			1353 => "0000000001010110011101",
			1354 => "0000000001010110011101",
			1355 => "0000000001010110011101",
			1356 => "0011110110010000100000",
			1357 => "0001101011001100001100",
			1358 => "0000101100111000001000",
			1359 => "0011111101000100000100",
			1360 => "0000000001010110011101",
			1361 => "0000000001010110011101",
			1362 => "0000000001010110011101",
			1363 => "0001001101110100001000",
			1364 => "0001000001101100000100",
			1365 => "0000000001010110011101",
			1366 => "0000000001010110011101",
			1367 => "0010111000000000001000",
			1368 => "0010110110000100000100",
			1369 => "0000000001010110011101",
			1370 => "0000001001010110011101",
			1371 => "0000000001010110011101",
			1372 => "0011011110101100001000",
			1373 => "0011111001100000000100",
			1374 => "0000000001010110011101",
			1375 => "1111111001010110011101",
			1376 => "0000010101011100001100",
			1377 => "0000100010110000001000",
			1378 => "0010001001101000000100",
			1379 => "0000000001010110011101",
			1380 => "0000001001010110011101",
			1381 => "0000000001010110011101",
			1382 => "0000000001010110011101",
			1383 => "0011010100011000000100",
			1384 => "1111111001011000111001",
			1385 => "0011000100001000111100",
			1386 => "0011101010111000011100",
			1387 => "0011111011011100000100",
			1388 => "1111111001011000111001",
			1389 => "0001101100011000001000",
			1390 => "0010111100101100000100",
			1391 => "0000010001011000111001",
			1392 => "0000000001011000111001",
			1393 => "0001000001100100001000",
			1394 => "0000111000000000000100",
			1395 => "0000000001011000111001",
			1396 => "0000000001011000111001",
			1397 => "0001111101100000000100",
			1398 => "0000000001011000111001",
			1399 => "0000001001011000111001",
			1400 => "0000010110101000000100",
			1401 => "1111111001011000111001",
			1402 => "0001010000011100010000",
			1403 => "0010011011111100001000",
			1404 => "0011001001110000000100",
			1405 => "0000000001011000111001",
			1406 => "0000001001011000111001",
			1407 => "0011010001011000000100",
			1408 => "1111111001011000111001",
			1409 => "0000000001011000111001",
			1410 => "0010010100111100001000",
			1411 => "0001101000010000000100",
			1412 => "0000001001011000111001",
			1413 => "0000000001011000111001",
			1414 => "0000000001011000111001",
			1415 => "0001101000010000000100",
			1416 => "1111111001011000111001",
			1417 => "0011110101000000001000",
			1418 => "0000011011111100000100",
			1419 => "0000001001011000111001",
			1420 => "0000000001011000111001",
			1421 => "1111111001011000111001",
			1422 => "0001001110111000000100",
			1423 => "1111111001011011110101",
			1424 => "0010000111000100111000",
			1425 => "0010000111000100100000",
			1426 => "0010000110001000011000",
			1427 => "0001000011101100001100",
			1428 => "0011101101101100001000",
			1429 => "0010100110011000000100",
			1430 => "0000000001011011110101",
			1431 => "0000001001011011110101",
			1432 => "0000000001011011110101",
			1433 => "0010001011010100001000",
			1434 => "0001111101010100000100",
			1435 => "0000000001011011110101",
			1436 => "0000000001011011110101",
			1437 => "0000000001011011110101",
			1438 => "0001000000101100000100",
			1439 => "0000000001011011110101",
			1440 => "0000000001011011110101",
			1441 => "0011110101110100001000",
			1442 => "0010111100001000000100",
			1443 => "0000000001011011110101",
			1444 => "0000010001011011110101",
			1445 => "0001000100001100000100",
			1446 => "0000000001011011110101",
			1447 => "0000011101011100001000",
			1448 => "0001010111001000000100",
			1449 => "0000000001011011110101",
			1450 => "0000001001011011110101",
			1451 => "0000000001011011110101",
			1452 => "0001100100111100011100",
			1453 => "0001000001100100000100",
			1454 => "1111111001011011110101",
			1455 => "0011001100110000001000",
			1456 => "0010111110001100000100",
			1457 => "0000000001011011110101",
			1458 => "0000001001011011110101",
			1459 => "0001101001100100001000",
			1460 => "0001000011111000000100",
			1461 => "0000000001011011110101",
			1462 => "1111111001011011110101",
			1463 => "0000011101011100000100",
			1464 => "0000000001011011110101",
			1465 => "0000000001011011110101",
			1466 => "0010011001100100000100",
			1467 => "1111111001011011110101",
			1468 => "0000000001011011110101",
			1469 => "0011010100011000000100",
			1470 => "1111111001011111001011",
			1471 => "0011000011011100011100",
			1472 => "0011100100001000001100",
			1473 => "0001001110111000000100",
			1474 => "0000000001011111001011",
			1475 => "0001101111000000000100",
			1476 => "0000001001011111001011",
			1477 => "0000000001011111001011",
			1478 => "0011000011011100001000",
			1479 => "0001001101000000000100",
			1480 => "1111111001011111001011",
			1481 => "0000000001011111001011",
			1482 => "0000110101110100000100",
			1483 => "0000000001011111001011",
			1484 => "0000001001011111001011",
			1485 => "0001101011001100011100",
			1486 => "0011001100110000001000",
			1487 => "0000001100001000000100",
			1488 => "0000000001011111001011",
			1489 => "0000000001011111001011",
			1490 => "0010110000001100001100",
			1491 => "0010110000001100000100",
			1492 => "0000000001011111001011",
			1493 => "0011010001101000000100",
			1494 => "0000000001011111001011",
			1495 => "1111101001011111001011",
			1496 => "0001111110001100000100",
			1497 => "0000000001011111001011",
			1498 => "1111111001011111001011",
			1499 => "0001101111000000011100",
			1500 => "0001001101110100001100",
			1501 => "0011011001010100000100",
			1502 => "1111111001011111001011",
			1503 => "0011000100001000000100",
			1504 => "0000000001011111001011",
			1505 => "0000000001011111001011",
			1506 => "0000000100010100001000",
			1507 => "0000100110101100000100",
			1508 => "0000001001011111001011",
			1509 => "0000000001011111001011",
			1510 => "0000111101010100000100",
			1511 => "0000000001011111001011",
			1512 => "0000001001011111001011",
			1513 => "0000101000011100001000",
			1514 => "0000110010110100000100",
			1515 => "0000000001011111001011",
			1516 => "1111111001011111001011",
			1517 => "0000111111101000001000",
			1518 => "0010100101000100000100",
			1519 => "0000001001011111001011",
			1520 => "0000000001011111001011",
			1521 => "1111111001011111001011",
			1522 => "0000000001011111001101",
			1523 => "0000000001011111010001",
			1524 => "0000000001011111010101",
			1525 => "0000000001011111011001",
			1526 => "0000000001011111011101",
			1527 => "0000000001011111100001",
			1528 => "0000000001011111100101",
			1529 => "0000000001011111101001",
			1530 => "0000000001011111101101",
			1531 => "0000000001011111110001",
			1532 => "0000100110010000000100",
			1533 => "0000000001011111111101",
			1534 => "0000000001011111111101",
			1535 => "0000011011101000000100",
			1536 => "0000000001100000010001",
			1537 => "0000010000111100000100",
			1538 => "0000000001100000010001",
			1539 => "0000000001100000010001",
			1540 => "0011000110000100001000",
			1541 => "0011000000101000000100",
			1542 => "0000000001100000100101",
			1543 => "0000000001100000100101",
			1544 => "0000000001100000100101",
			1545 => "0001101000010000001000",
			1546 => "0001100100110100000100",
			1547 => "0000000001100000111001",
			1548 => "0000000001100000111001",
			1549 => "0000000001100000111001",
			1550 => "0011101110101100001000",
			1551 => "0001001101000000000100",
			1552 => "0000000001100001001101",
			1553 => "0000000001100001001101",
			1554 => "0000000001100001001101",
			1555 => "0011110110010000001000",
			1556 => "0011110010001000000100",
			1557 => "0000000001100001101001",
			1558 => "0000000001100001101001",
			1559 => "0011111011110000000100",
			1560 => "0000000001100001101001",
			1561 => "0000000001100001101001",
			1562 => "0011110010000000001000",
			1563 => "0011110010001000000100",
			1564 => "0000000001100010000101",
			1565 => "0000000001100010000101",
			1566 => "0011111000110100000100",
			1567 => "0000000001100010000101",
			1568 => "0000000001100010000101",
			1569 => "0000100100101000000100",
			1570 => "0000000001100010100001",
			1571 => "0001001101110100001000",
			1572 => "0011101010000100000100",
			1573 => "0000000001100010100001",
			1574 => "0000000001100010100001",
			1575 => "0000000001100010100001",
			1576 => "0000001000111100001100",
			1577 => "0000000011111100000100",
			1578 => "0000000001100010111101",
			1579 => "0011110101110100000100",
			1580 => "0000000001100010111101",
			1581 => "0000000001100010111101",
			1582 => "0000000001100010111101",
			1583 => "0010000110001000000100",
			1584 => "0000000001100011011001",
			1585 => "0011001000111100000100",
			1586 => "0000000001100011011001",
			1587 => "0000000000111000000100",
			1588 => "0000000001100011011001",
			1589 => "0000000001100011011001",
			1590 => "0011101100101100000100",
			1591 => "0000000001100011110101",
			1592 => "0010100110011000000100",
			1593 => "0000000001100011110101",
			1594 => "0011101101101100000100",
			1595 => "0000000001100011110101",
			1596 => "0000000001100011110101",
			1597 => "0011110010000000001000",
			1598 => "0011110010001000000100",
			1599 => "0000000001100100011001",
			1600 => "0000000001100100011001",
			1601 => "0011111000110100001000",
			1602 => "0011110110010000000100",
			1603 => "0000000001100100011001",
			1604 => "0000000001100100011001",
			1605 => "0000000001100100011001",
			1606 => "0011000011011100001100",
			1607 => "0001111001110000000100",
			1608 => "0000000001100101000101",
			1609 => "0011010100011000000100",
			1610 => "0000000001100101000101",
			1611 => "0000000001100101000101",
			1612 => "0011011001010100001000",
			1613 => "0001110110000100000100",
			1614 => "0000000001100101000101",
			1615 => "0000000001100101000101",
			1616 => "0000000001100101000101",
			1617 => "0001001100111100001100",
			1618 => "0000100100101000000100",
			1619 => "0000000001100101110001",
			1620 => "0000101110100100000100",
			1621 => "0000000001100101110001",
			1622 => "0000000001100101110001",
			1623 => "0011010001011000000100",
			1624 => "0000000001100101110001",
			1625 => "0011011001010000000100",
			1626 => "0000000001100101110001",
			1627 => "0000000001100101110001",
			1628 => "0001111100101000010000",
			1629 => "0001111001110000000100",
			1630 => "0000000001100110010101",
			1631 => "0011001100110000001000",
			1632 => "0011000000101000000100",
			1633 => "0000000001100110010101",
			1634 => "0000000001100110010101",
			1635 => "0000000001100110010101",
			1636 => "0000000001100110010101",
			1637 => "0011001100110000010000",
			1638 => "0000011100110100000100",
			1639 => "0000000001100110111001",
			1640 => "0000011111001100001000",
			1641 => "0011000000101000000100",
			1642 => "0000000001100110111001",
			1643 => "0000000001100110111001",
			1644 => "0000000001100110111001",
			1645 => "0000000001100110111001",
			1646 => "0011101100101100000100",
			1647 => "0000000001100111011101",
			1648 => "0010100110011000000100",
			1649 => "0000000001100111011101",
			1650 => "0011101101101100001000",
			1651 => "0010101100000100000100",
			1652 => "0000000001100111011101",
			1653 => "0000000001100111011101",
			1654 => "0000000001100111011101",
			1655 => "0010011101101000000100",
			1656 => "0000000001101000000001",
			1657 => "0010011101011000001100",
			1658 => "0010110101101100000100",
			1659 => "0000000001101000000001",
			1660 => "0010111011110100000100",
			1661 => "0000000001101000000001",
			1662 => "0000000001101000000001",
			1663 => "0000000001101000000001",
			1664 => "0011001100110000010000",
			1665 => "0001111001110000000100",
			1666 => "0000000001101000110101",
			1667 => "0001111100101000001000",
			1668 => "0011000000101000000100",
			1669 => "0000000001101000110101",
			1670 => "0000000001101000110101",
			1671 => "0000000001101000110101",
			1672 => "0010100001010000000100",
			1673 => "0000000001101000110101",
			1674 => "0010101100000100000100",
			1675 => "0000000001101000110101",
			1676 => "0000000001101000110101",
			1677 => "0000000011111100001100",
			1678 => "0010100110011000000100",
			1679 => "0000000001101001101001",
			1680 => "0010100001010000000100",
			1681 => "0000000001101001101001",
			1682 => "0000000001101001101001",
			1683 => "0001000001100100001100",
			1684 => "0011110101110100000100",
			1685 => "0000000001101001101001",
			1686 => "0011000000001100000100",
			1687 => "0000000001101001101001",
			1688 => "0000000001101001101001",
			1689 => "0000000001101001101001",
			1690 => "0001001100111100001100",
			1691 => "0000100100101000000100",
			1692 => "0000000001101010011101",
			1693 => "0011111011110000000100",
			1694 => "0000000001101010011101",
			1695 => "0000000001101010011101",
			1696 => "0001101101011000000100",
			1697 => "0000000001101010011101",
			1698 => "0001101000010000001000",
			1699 => "0011010101100100000100",
			1700 => "0000000001101010011101",
			1701 => "0000000001101010011101",
			1702 => "0000000001101010011101",
			1703 => "0001000001100100010000",
			1704 => "0010100001010000000100",
			1705 => "0000000001101011011001",
			1706 => "0011110101110100000100",
			1707 => "0000000001101011011001",
			1708 => "0000000010011000000100",
			1709 => "0000000001101011011001",
			1710 => "0000000001101011011001",
			1711 => "0000011111001100001100",
			1712 => "0000010010001100000100",
			1713 => "0000000001101011011001",
			1714 => "0011111000001100000100",
			1715 => "0000000001101011011001",
			1716 => "0000000001101011011001",
			1717 => "0000000001101011011001",
			1718 => "0011100111110000001000",
			1719 => "0001010100010000000100",
			1720 => "0000000001101100001101",
			1721 => "0000000001101100001101",
			1722 => "0000010101011100010000",
			1723 => "0000011011101000000100",
			1724 => "0000000001101100001101",
			1725 => "0001010101100100000100",
			1726 => "0000000001101100001101",
			1727 => "0001010111111100000100",
			1728 => "0000000001101100001101",
			1729 => "0000000001101100001101",
			1730 => "0000000001101100001101",
			1731 => "0001101101011000001000",
			1732 => "0001001110111000000100",
			1733 => "0000000001101101001001",
			1734 => "0000000001101101001001",
			1735 => "0001101001100100010000",
			1736 => "0000010111100100000100",
			1737 => "0000000001101101001001",
			1738 => "0000010000111100001000",
			1739 => "0001001000000100000100",
			1740 => "0000000001101101001001",
			1741 => "0000000001101101001001",
			1742 => "0000000001101101001001",
			1743 => "0001000011111000000100",
			1744 => "0000000001101101001001",
			1745 => "0000000001101101001001",
			1746 => "0010010100110100010000",
			1747 => "0011111110101000000100",
			1748 => "0000000001101110001101",
			1749 => "0001001010010000001000",
			1750 => "0001010100010000000100",
			1751 => "0000000001101110001101",
			1752 => "0000000001101110001101",
			1753 => "0000000001101110001101",
			1754 => "0000010000111100010000",
			1755 => "0010010100111100001100",
			1756 => "0000010000111100001000",
			1757 => "0000011011101000000100",
			1758 => "0000000001101110001101",
			1759 => "0000000001101110001101",
			1760 => "0000000001101110001101",
			1761 => "0000000001101110001101",
			1762 => "0000000001101110001101",
			1763 => "0000110101110100001000",
			1764 => "0000110010001000000100",
			1765 => "0000000001101111001001",
			1766 => "0000000001101111001001",
			1767 => "0000010101011100010100",
			1768 => "0000011011101000000100",
			1769 => "0000000001101111001001",
			1770 => "0011100100010000000100",
			1771 => "0000000001101111001001",
			1772 => "0000111110101100000100",
			1773 => "0000000001101111001001",
			1774 => "0000110010010100000100",
			1775 => "0000000001101111001001",
			1776 => "0000000001101111001001",
			1777 => "0000000001101111001001",
			1778 => "0001000011101100001100",
			1779 => "0001101000010000001000",
			1780 => "0010101010110000000100",
			1781 => "0000000001110000001101",
			1782 => "0000000001110000001101",
			1783 => "0000000001110000001101",
			1784 => "0001101000010000010100",
			1785 => "0001110100011000010000",
			1786 => "0001101101011000000100",
			1787 => "0000000001110000001101",
			1788 => "0010011001011000000100",
			1789 => "0000000001110000001101",
			1790 => "0010100110011000000100",
			1791 => "0000000001110000001101",
			1792 => "0000000001110000001101",
			1793 => "0000000001110000001101",
			1794 => "0000000001110000001101",
			1795 => "0000000010111100010100",
			1796 => "0000000010011000000100",
			1797 => "0000000001110001100001",
			1798 => "0001011000000000000100",
			1799 => "0000000001110001100001",
			1800 => "0000010101011100001000",
			1801 => "0010001011010100000100",
			1802 => "0000000001110001100001",
			1803 => "0000000001110001100001",
			1804 => "0000000001110001100001",
			1805 => "0011111010010100001000",
			1806 => "0011101001110000000100",
			1807 => "0000000001110001100001",
			1808 => "0000000001110001100001",
			1809 => "0001000001100100001100",
			1810 => "0000101010001000000100",
			1811 => "0000000001110001100001",
			1812 => "0011101010000100000100",
			1813 => "0000000001110001100001",
			1814 => "0000000001110001100001",
			1815 => "0000000001110001100001",
			1816 => "0011101100101100000100",
			1817 => "0000000001110010010101",
			1818 => "0010100110011000000100",
			1819 => "0000000001110010010101",
			1820 => "0001110110100100010000",
			1821 => "0010011101101000000100",
			1822 => "0000000001110010010101",
			1823 => "0000010101011100001000",
			1824 => "0001111001110000000100",
			1825 => "0000000001110010010101",
			1826 => "0000000001110010010101",
			1827 => "0000000001110010010101",
			1828 => "0000000001110010010101",
			1829 => "0011001100110000011000",
			1830 => "0011010100011000000100",
			1831 => "0000000001110011100001",
			1832 => "0010001001101000000100",
			1833 => "0000000001110011100001",
			1834 => "0000100110111000001100",
			1835 => "0000000010111100000100",
			1836 => "0000000001110011100001",
			1837 => "0001111001110000000100",
			1838 => "0000000001110011100001",
			1839 => "0000000001110011100001",
			1840 => "0000000001110011100001",
			1841 => "0000101011111000000100",
			1842 => "0000000001110011100001",
			1843 => "0000000010111100000100",
			1844 => "0000000001110011100001",
			1845 => "0000001010111100000100",
			1846 => "0000000001110011100001",
			1847 => "0000000001110011100001",
			1848 => "0000000010111100010100",
			1849 => "0000000010011000000100",
			1850 => "0000000001110100111101",
			1851 => "0001011000000000000100",
			1852 => "0000000001110100111101",
			1853 => "0010001011010100001000",
			1854 => "0001000010100100000100",
			1855 => "0000000001110100111101",
			1856 => "0000000001110100111101",
			1857 => "0000000001110100111101",
			1858 => "0011111010010100001100",
			1859 => "0011101001110000000100",
			1860 => "0000000001110100111101",
			1861 => "0000111010111100000100",
			1862 => "0000000001110100111101",
			1863 => "0000000001110100111101",
			1864 => "0000001010111100001100",
			1865 => "0011101001100000001000",
			1866 => "0000101010001000000100",
			1867 => "0000000001110100111101",
			1868 => "0000000001110100111101",
			1869 => "0000000001110100111101",
			1870 => "0000000001110100111101",
			1871 => "0010010001000100001000",
			1872 => "0001000011111000000100",
			1873 => "0000000001110110001001",
			1874 => "0000000001110110001001",
			1875 => "0000011111001100011000",
			1876 => "0001101011001100000100",
			1877 => "0000000001110110001001",
			1878 => "0000111001011100010000",
			1879 => "0000000010111100000100",
			1880 => "0000000001110110001001",
			1881 => "0010111110001100000100",
			1882 => "0000000001110110001001",
			1883 => "0001101000010000000100",
			1884 => "0000000001110110001001",
			1885 => "0000000001110110001001",
			1886 => "0000000001110110001001",
			1887 => "0011110010000000000100",
			1888 => "0000000001110110001001",
			1889 => "0000000001110110001001",
			1890 => "0001000011101100001100",
			1891 => "0001101000010000001000",
			1892 => "0010101010110000000100",
			1893 => "0000000001110111010101",
			1894 => "0000000001110111010101",
			1895 => "0000000001110111010101",
			1896 => "0001101000010000011000",
			1897 => "0001110100011000010100",
			1898 => "0001101101011000000100",
			1899 => "0000000001110111010101",
			1900 => "0000011001111000000100",
			1901 => "0000000001110111010101",
			1902 => "0010100110011000000100",
			1903 => "0000000001110111010101",
			1904 => "0001111101100000000100",
			1905 => "0000000001110111010101",
			1906 => "0000000001110111010101",
			1907 => "0000000001110111010101",
			1908 => "0000000001110111010101",
			1909 => "0011110110010000011100",
			1910 => "0011000000101000000100",
			1911 => "0000000001111000011001",
			1912 => "0010101001000100000100",
			1913 => "0000000001111000011001",
			1914 => "0011111011011100000100",
			1915 => "0000000001111000011001",
			1916 => "0000101011101100001100",
			1917 => "0010100001110000001000",
			1918 => "0011001110001100000100",
			1919 => "0000000001111000011001",
			1920 => "0000000001111000011001",
			1921 => "0000000001111000011001",
			1922 => "0000000001111000011001",
			1923 => "0011000011011100000100",
			1924 => "0000000001111000011001",
			1925 => "0000000001111000011001",
			1926 => "0001000011010100011000",
			1927 => "0000100100101000010000",
			1928 => "0010110101101100000100",
			1929 => "0000000001111010001101",
			1930 => "0010110110000100001000",
			1931 => "0001100100110100000100",
			1932 => "0000000001111010001101",
			1933 => "0000000001111010001101",
			1934 => "0000000001111010001101",
			1935 => "0001110111010000000100",
			1936 => "0000000001111010001101",
			1937 => "0000000001111010001101",
			1938 => "0010100101000100010000",
			1939 => "0000010101011100001100",
			1940 => "0010100110011000000100",
			1941 => "0000000001111010001101",
			1942 => "0011010100011000000100",
			1943 => "0000000001111010001101",
			1944 => "0000000001111010001101",
			1945 => "0000000001111010001101",
			1946 => "0011110001000000000100",
			1947 => "0000000001111010001101",
			1948 => "0000101011101100000100",
			1949 => "0000000001111010001101",
			1950 => "0000111111011100000100",
			1951 => "0000000001111010001101",
			1952 => "0011011011110100000100",
			1953 => "0000000001111010001101",
			1954 => "0000000001111010001101",
			1955 => "0001101011001100010000",
			1956 => "0010011001100100001100",
			1957 => "0011111010010100000100",
			1958 => "0000000001111011100001",
			1959 => "0010101100000100000100",
			1960 => "0000000001111011100001",
			1961 => "0000000001111011100001",
			1962 => "0000000001111011100001",
			1963 => "0010011101011000011000",
			1964 => "0010010001000100000100",
			1965 => "0000000001111011100001",
			1966 => "0000111001011100010000",
			1967 => "0011000011011100000100",
			1968 => "0000000001111011100001",
			1969 => "0001001000000100000100",
			1970 => "0000000001111011100001",
			1971 => "0010101100000100000100",
			1972 => "0000000001111011100001",
			1973 => "0000000001111011100001",
			1974 => "0000000001111011100001",
			1975 => "0000000001111011100001",
			1976 => "0011110000010000100100",
			1977 => "0000110101110100001100",
			1978 => "0001001101000000001000",
			1979 => "0011111010010100000100",
			1980 => "0000000001111100110101",
			1981 => "0000000001111100110101",
			1982 => "0000000001111100110101",
			1983 => "0000010111100100000100",
			1984 => "0000000001111100110101",
			1985 => "0011000100001000010000",
			1986 => "0001101011001100000100",
			1987 => "0000000001111100110101",
			1988 => "0011000011011100000100",
			1989 => "0000000001111100110101",
			1990 => "0001001000000100000100",
			1991 => "0000000001111100110101",
			1992 => "0000000001111100110101",
			1993 => "0000000001111100110101",
			1994 => "0000000010011000000100",
			1995 => "0000000001111100110101",
			1996 => "0000000001111100110101",
			1997 => "0011010100011000000100",
			1998 => "0000000001111101110001",
			1999 => "0001111100101000011000",
			2000 => "0000000010111100000100",
			2001 => "0000000001111101110001",
			2002 => "0000111001011100010000",
			2003 => "0010000111000100001100",
			2004 => "0011001110001100001000",
			2005 => "0001111001110000000100",
			2006 => "0000000001111101110001",
			2007 => "0000000001111101110001",
			2008 => "0000000001111101110001",
			2009 => "0000000001111101110001",
			2010 => "0000000001111101110001",
			2011 => "0000000001111101110001",
			2012 => "0000010110101000000100",
			2013 => "0000000001111110101101",
			2014 => "0000010101011100011000",
			2015 => "0010101001000100000100",
			2016 => "0000000001111110101101",
			2017 => "0001111001110000000100",
			2018 => "0000000001111110101101",
			2019 => "0011011001110100000100",
			2020 => "0000000001111110101101",
			2021 => "0001100101010000001000",
			2022 => "0011001000111000000100",
			2023 => "0000000001111110101101",
			2024 => "0000000001111110101101",
			2025 => "0000000001111110101101",
			2026 => "0000000001111110101101",
			2027 => "0011101100101100000100",
			2028 => "0000000001111111101001",
			2029 => "0001111100101000011000",
			2030 => "0010001001101000000100",
			2031 => "0000000001111111101001",
			2032 => "0010011101101000000100",
			2033 => "0000000001111111101001",
			2034 => "0001111001110000000100",
			2035 => "0000000001111111101001",
			2036 => "0001101000010000001000",
			2037 => "0001001000000100000100",
			2038 => "0000000001111111101001",
			2039 => "0000000001111111101001",
			2040 => "0000000001111111101001",
			2041 => "0000000001111111101001",
			2042 => "0000010110101000010100",
			2043 => "0011111010010100001100",
			2044 => "0011101001110000000100",
			2045 => "0000000010000001011101",
			2046 => "0001001110111000000100",
			2047 => "0000000010000001011101",
			2048 => "0000000010000001011101",
			2049 => "0010000010111100000100",
			2050 => "0000000010000001011101",
			2051 => "0000000010000001011101",
			2052 => "0000011111001100011000",
			2053 => "0000000010111100000100",
			2054 => "0000000010000001011101",
			2055 => "0001111001110000000100",
			2056 => "0000000010000001011101",
			2057 => "0000111001011100001100",
			2058 => "0001011000000000000100",
			2059 => "0000000010000001011101",
			2060 => "0011001000111000000100",
			2061 => "0000000010000001011101",
			2062 => "0000000010000001011101",
			2063 => "0000000010000001011101",
			2064 => "0000100110101100000100",
			2065 => "0000000010000001011101",
			2066 => "0001111101111000000100",
			2067 => "0000000010000001011101",
			2068 => "0001110111010000000100",
			2069 => "0000000010000001011101",
			2070 => "0000000010000001011101",
			2071 => "0000100110101100011100",
			2072 => "0010011101101000000100",
			2073 => "0000000010000010111001",
			2074 => "0000000010111100000100",
			2075 => "0000000010000010111001",
			2076 => "0010110101101100000100",
			2077 => "0000000010000010111001",
			2078 => "0001101001100100001100",
			2079 => "0010001001101000000100",
			2080 => "0000000010000010111001",
			2081 => "0001111001110000000100",
			2082 => "0000000010000010111001",
			2083 => "0000000010000010111001",
			2084 => "0000000010000010111001",
			2085 => "0011001100110000000100",
			2086 => "0000000010000010111001",
			2087 => "0011101010000100001100",
			2088 => "0000000010111100000100",
			2089 => "0000000010000010111001",
			2090 => "0000001010111100000100",
			2091 => "0000000010000010111001",
			2092 => "0000000010000010111001",
			2093 => "0000000010000010111001",
			2094 => "0001111100101000100100",
			2095 => "0011010100011000000100",
			2096 => "0000000010000100010101",
			2097 => "0001101000010000011100",
			2098 => "0001000011010100010000",
			2099 => "0010001011010100001100",
			2100 => "0001111101100000001000",
			2101 => "0010001001101000000100",
			2102 => "0000000010000100010101",
			2103 => "0000000010000100010101",
			2104 => "0000000010000100010101",
			2105 => "0000000010000100010101",
			2106 => "0000011100110100000100",
			2107 => "0000000010000100010101",
			2108 => "0010001011010100000100",
			2109 => "0000000010000100010101",
			2110 => "0000000010000100010101",
			2111 => "0000000010000100010101",
			2112 => "0011011001010100001000",
			2113 => "0000100000010000000100",
			2114 => "0000000010000100010101",
			2115 => "0000000010000100010101",
			2116 => "0000000010000100010101",
			2117 => "0011010100011000000100",
			2118 => "1111111010000101111001",
			2119 => "0001111100101000100100",
			2120 => "0010000111000100010000",
			2121 => "0000000010111100000100",
			2122 => "0000000010000101111001",
			2123 => "0001111001110000000100",
			2124 => "0000000010000101111001",
			2125 => "0001101000010000000100",
			2126 => "0000001010000101111001",
			2127 => "0000000010000101111001",
			2128 => "0001001101000000001000",
			2129 => "0010110000001100000100",
			2130 => "0000000010000101111001",
			2131 => "0000000010000101111001",
			2132 => "0001101101011000000100",
			2133 => "0000000010000101111001",
			2134 => "0000000001001000000100",
			2135 => "0000000010000101111001",
			2136 => "0000000010000101111001",
			2137 => "0000101000100000001000",
			2138 => "0010100110011000000100",
			2139 => "0000000010000101111001",
			2140 => "0000000010000101111001",
			2141 => "0000000010000101111001",
			2142 => "0001111001110000001000",
			2143 => "0000101000100000000100",
			2144 => "1111111010000111011101",
			2145 => "0000000010000111011101",
			2146 => "0011000100001000011100",
			2147 => "0010100111000100011000",
			2148 => "0000000010011000000100",
			2149 => "1111111010000111011101",
			2150 => "0000100100101000000100",
			2151 => "0000010010000111011101",
			2152 => "0010111100101100001000",
			2153 => "0001000010010000000100",
			2154 => "1111111010000111011101",
			2155 => "0000000010000111011101",
			2156 => "0001101000010000000100",
			2157 => "0000000010000111011101",
			2158 => "1111111010000111011101",
			2159 => "1111111010000111011101",
			2160 => "0000100101000000000100",
			2161 => "1111111010000111011101",
			2162 => "0000111111101000001000",
			2163 => "0000111101101100000100",
			2164 => "0000000010000111011101",
			2165 => "0000001010000111011101",
			2166 => "1111111010000111011101",
			2167 => "0000000010111100011000",
			2168 => "0010001001101000000100",
			2169 => "0000000010001001100001",
			2170 => "0011001000111000000100",
			2171 => "0000000010001001100001",
			2172 => "0000010101011100001100",
			2173 => "0010001011010100001000",
			2174 => "0001001000000100000100",
			2175 => "0000000010001001100001",
			2176 => "0000001010001001100001",
			2177 => "0000000010001001100001",
			2178 => "0000000010001001100001",
			2179 => "0001101100011000010000",
			2180 => "0000110100011000000100",
			2181 => "0000000010001001100001",
			2182 => "0000010010001100000100",
			2183 => "0000000010001001100001",
			2184 => "0001000011001100000100",
			2185 => "0000000010001001100001",
			2186 => "0000000010001001100001",
			2187 => "0001001011001000000100",
			2188 => "0000000010001001100001",
			2189 => "0001101111000000010000",
			2190 => "0011101001010100001100",
			2191 => "0000011111001100001000",
			2192 => "0010011001011000000100",
			2193 => "0000000010001001100001",
			2194 => "0000000010001001100001",
			2195 => "0000000010001001100001",
			2196 => "0000000010001001100001",
			2197 => "0001000101001100000100",
			2198 => "0000000010001001100001",
			2199 => "0000000010001001100001",
			2200 => "0011110110010000110100",
			2201 => "0001111001110000001000",
			2202 => "0010100110001000000100",
			2203 => "0000000010001011011101",
			2204 => "0000000010001011011101",
			2205 => "0001111101100000010100",
			2206 => "0000100110010000010000",
			2207 => "0011101001110000000100",
			2208 => "0000000010001011011101",
			2209 => "0000000010111100000100",
			2210 => "0000000010001011011101",
			2211 => "0010000111000100000100",
			2212 => "0000001010001011011101",
			2213 => "0000000010001011011101",
			2214 => "0000000010001011011101",
			2215 => "0010001010101100001100",
			2216 => "0011110011001000001000",
			2217 => "0000111010111000000100",
			2218 => "0000000010001011011101",
			2219 => "0000000010001011011101",
			2220 => "0000000010001011011101",
			2221 => "0001101101011000000100",
			2222 => "0000000010001011011101",
			2223 => "0000000101100100000100",
			2224 => "0000000010001011011101",
			2225 => "0000000010001011011101",
			2226 => "0010110110100100000100",
			2227 => "0000000010001011011101",
			2228 => "0011000100001000000100",
			2229 => "0000000010001011011101",
			2230 => "0000000010001011011101",
			2231 => "0001001110111000000100",
			2232 => "0000000010001101000001",
			2233 => "0010000111000100011000",
			2234 => "0000010101011100010100",
			2235 => "0000011100110100000100",
			2236 => "0000000010001101000001",
			2237 => "0010101100011100001100",
			2238 => "0010100110011000000100",
			2239 => "0000000010001101000001",
			2240 => "0011010100011000000100",
			2241 => "0000000010001101000001",
			2242 => "0000000010001101000001",
			2243 => "0000000010001101000001",
			2244 => "0000000010001101000001",
			2245 => "0001100100111100010100",
			2246 => "0001000110110000001000",
			2247 => "0000011101011100000100",
			2248 => "0000000010001101000001",
			2249 => "0000000010001101000001",
			2250 => "0001101011001100000100",
			2251 => "0000000010001101000001",
			2252 => "0000010010001100000100",
			2253 => "0000000010001101000001",
			2254 => "0000000010001101000001",
			2255 => "0000000010001101000001",
			2256 => "0001001001000000100100",
			2257 => "0001000011010100001100",
			2258 => "0000100101000000000100",
			2259 => "1111111010001111000101",
			2260 => "0000100101000000000100",
			2261 => "0000000010001111000101",
			2262 => "1111111010001111000101",
			2263 => "0010000110001000010100",
			2264 => "0010100110011000001100",
			2265 => "0001000011110100001000",
			2266 => "0001101101011000000100",
			2267 => "0000000010001111000101",
			2268 => "0000001010001111000101",
			2269 => "1111111010001111000101",
			2270 => "0011001000011000000100",
			2271 => "0000010010001111000101",
			2272 => "0000000010001111000101",
			2273 => "1111111010001111000101",
			2274 => "0000111110001100000100",
			2275 => "1111111010001111000101",
			2276 => "0001101000010000011000",
			2277 => "0011000100001000010100",
			2278 => "0001010100011000000100",
			2279 => "1111111010001111000101",
			2280 => "0000101011111000001000",
			2281 => "0010100110011000000100",
			2282 => "0000000010001111000101",
			2283 => "0000001010001111000101",
			2284 => "0001001100111100000100",
			2285 => "1111111010001111000101",
			2286 => "0000001010001111000101",
			2287 => "1111111010001111000101",
			2288 => "1111111010001111000101",
			2289 => "0001000001100100111000",
			2290 => "0001000011101100011100",
			2291 => "0001001110111000000100",
			2292 => "1100000010010001110001",
			2293 => "0010001011010100001100",
			2294 => "0000110010010100001000",
			2295 => "0010100110011000000100",
			2296 => "1100000010010001110001",
			2297 => "1110001010010001110001",
			2298 => "1100000010010001110001",
			2299 => "0010110101101100000100",
			2300 => "1100000010010001110001",
			2301 => "0011010011100000000100",
			2302 => "1100010010010001110001",
			2303 => "1100000010010001110001",
			2304 => "0001011011011100001100",
			2305 => "0001010011100000000100",
			2306 => "1100000010010001110001",
			2307 => "0000110111110000000100",
			2308 => "1100110010010001110001",
			2309 => "1100000010010001110001",
			2310 => "0010100001010000000100",
			2311 => "1110000010010001110001",
			2312 => "0010000110001000001000",
			2313 => "0000011001011000000100",
			2314 => "1101001010010001110001",
			2315 => "1100000010010001110001",
			2316 => "1100000010010001110001",
			2317 => "0000010010001100000100",
			2318 => "1100000010010001110001",
			2319 => "0011111100010100001100",
			2320 => "0001001011100100001000",
			2321 => "0011011011011100000100",
			2322 => "1100000010010001110001",
			2323 => "1111110010010001110001",
			2324 => "0001000010010001110001",
			2325 => "0011000100001000001100",
			2326 => "0001000110110000001000",
			2327 => "0010110011100000000100",
			2328 => "1100000010010001110001",
			2329 => "1100110010010001110001",
			2330 => "1111010010010001110001",
			2331 => "1100000010010001110001",
			2332 => "0011010100011000000100",
			2333 => "0000000010010011100101",
			2334 => "0000101110010000001100",
			2335 => "0000000010111100000100",
			2336 => "0000000010010011100101",
			2337 => "0011000011011100000100",
			2338 => "0000000010010011100101",
			2339 => "0000000010010011100101",
			2340 => "0000011011101000001100",
			2341 => "0011100000001100000100",
			2342 => "0000000010010011100101",
			2343 => "0000001010111100000100",
			2344 => "0000000010010011100101",
			2345 => "0000000010010011100101",
			2346 => "0000011111001100001100",
			2347 => "0010101100011100000100",
			2348 => "0000000010010011100101",
			2349 => "0011111111100100000100",
			2350 => "0000000010010011100101",
			2351 => "0000000010010011100101",
			2352 => "0000100110101100001100",
			2353 => "0001010101100100000100",
			2354 => "0000000010010011100101",
			2355 => "0011101110101000000100",
			2356 => "0000000010010011100101",
			2357 => "0000000010010011100101",
			2358 => "0000101000011100000100",
			2359 => "0000000010010011100101",
			2360 => "0000000010010011100101",
			2361 => "0001000000010100000100",
			2362 => "1111111010010101110001",
			2363 => "0010000111000100101000",
			2364 => "0000001110111100011000",
			2365 => "0000101011111000001100",
			2366 => "0010100110011000000100",
			2367 => "0000000010010101110001",
			2368 => "0011001001110000000100",
			2369 => "0000000010010101110001",
			2370 => "0000000010010101110001",
			2371 => "0011101011111000000100",
			2372 => "0000000010010101110001",
			2373 => "0000100011110000000100",
			2374 => "0000000010010101110001",
			2375 => "0000000010010101110001",
			2376 => "0010001111001000000100",
			2377 => "0000000010010101110001",
			2378 => "0000000111111000001000",
			2379 => "0000111010111100000100",
			2380 => "0000000010010101110001",
			2381 => "0000001010010101110001",
			2382 => "0000000010010101110001",
			2383 => "0011111001100000010100",
			2384 => "0010011001011000001000",
			2385 => "0000101011101100000100",
			2386 => "0000000010010101110001",
			2387 => "0000000010010101110001",
			2388 => "0010011010011000001000",
			2389 => "0010111010111100000100",
			2390 => "0000000010010101110001",
			2391 => "0000001010010101110001",
			2392 => "0000000010010101110001",
			2393 => "0000011011101000000100",
			2394 => "1111111010010101110001",
			2395 => "0000000010010101110001",
			2396 => "0001000000010100000100",
			2397 => "1111111010010111110101",
			2398 => "0010000111000100100100",
			2399 => "0000001110111100010100",
			2400 => "0001101011001100001000",
			2401 => "0001101101011000000100",
			2402 => "0000000010010111110101",
			2403 => "0000000010010111110101",
			2404 => "0011001110001100000100",
			2405 => "0000000010010111110101",
			2406 => "0011001001110100000100",
			2407 => "0000000010010111110101",
			2408 => "0000000010010111110101",
			2409 => "0010001111001000000100",
			2410 => "0000000010010111110101",
			2411 => "0000000111111000001000",
			2412 => "0000111010111100000100",
			2413 => "0000000010010111110101",
			2414 => "0000001010010111110101",
			2415 => "0000000010010111110101",
			2416 => "0001100100111100011000",
			2417 => "0001011001110100001000",
			2418 => "0000001110001100000100",
			2419 => "0000000010010111110101",
			2420 => "0000000010010111110101",
			2421 => "0001101011001100000100",
			2422 => "0000000010010111110101",
			2423 => "0010011010011000001000",
			2424 => "0001000010010000000100",
			2425 => "0000000010010111110101",
			2426 => "0000001010010111110101",
			2427 => "0000000010010111110101",
			2428 => "1111111010010111110101",
			2429 => "0001000011010100001100",
			2430 => "0000100101000000000100",
			2431 => "1111111010011010001001",
			2432 => "0011110101000000000100",
			2433 => "0000001010011010001001",
			2434 => "1111111010011010001001",
			2435 => "0000011001111000011000",
			2436 => "0010000111000100001000",
			2437 => "0010001111001000000100",
			2438 => "0000000010011010001001",
			2439 => "0000011010011010001001",
			2440 => "0000101000101000001100",
			2441 => "0000010010001100000100",
			2442 => "1111111010011010001001",
			2443 => "0000010010001100000100",
			2444 => "0000000010011010001001",
			2445 => "1111111010011010001001",
			2446 => "0000000010011010001001",
			2447 => "0000100011110000100100",
			2448 => "0000111010011100001000",
			2449 => "0001010011100000000100",
			2450 => "0000000010011010001001",
			2451 => "0000001010011010001001",
			2452 => "0001101011001100001100",
			2453 => "0011001100110000000100",
			2454 => "0000000010011010001001",
			2455 => "0000100000010000000100",
			2456 => "0000000010011010001001",
			2457 => "1111111010011010001001",
			2458 => "0001000000101100001000",
			2459 => "0010111000000000000100",
			2460 => "1111111010011010001001",
			2461 => "0000001010011010001001",
			2462 => "0000011101011100000100",
			2463 => "0000001010011010001001",
			2464 => "1111111010011010001001",
			2465 => "1111111010011010001001",
			2466 => "0001001001000000011100",
			2467 => "0001000100001100000100",
			2468 => "1111111010011100000101",
			2469 => "0000001110111100010100",
			2470 => "0000100100101000000100",
			2471 => "0000011010011100000101",
			2472 => "0010101010110000001100",
			2473 => "0000101111100100000100",
			2474 => "1111111010011100000101",
			2475 => "0001010110010000000100",
			2476 => "0000001010011100000101",
			2477 => "0000000010011100000101",
			2478 => "1111111010011100000101",
			2479 => "1111111010011100000101",
			2480 => "0000011100110100000100",
			2481 => "1111111010011100000101",
			2482 => "0001101000010000011100",
			2483 => "0011000000101000000100",
			2484 => "0000101010011100000101",
			2485 => "0000011001111000001000",
			2486 => "0011100101101100000100",
			2487 => "0000001010011100000101",
			2488 => "1111111010011100000101",
			2489 => "0000101011111000001000",
			2490 => "0001101001100100000100",
			2491 => "0000001010011100000101",
			2492 => "0000000010011100000101",
			2493 => "0000011101011100000100",
			2494 => "0000001010011100000101",
			2495 => "1111111010011100000101",
			2496 => "1111111010011100000101",
			2497 => "0010011101101000000100",
			2498 => "0000000010011101111001",
			2499 => "0011000011011100011000",
			2500 => "0011011011000000000100",
			2501 => "0000000010011101111001",
			2502 => "0011001000111000000100",
			2503 => "0000000010011101111001",
			2504 => "0010001001101000000100",
			2505 => "0000000010011101111001",
			2506 => "0001101000010000001000",
			2507 => "0001111001110000000100",
			2508 => "0000000010011101111001",
			2509 => "0000000010011101111001",
			2510 => "0000000010011101111001",
			2511 => "0000100011110000011100",
			2512 => "0010110100011000001100",
			2513 => "0001001101000000001000",
			2514 => "0011100000001100000100",
			2515 => "0000000010011101111001",
			2516 => "0000000010011101111001",
			2517 => "0000000010011101111001",
			2518 => "0010100110011000000100",
			2519 => "0000000010011101111001",
			2520 => "0000011011101000000100",
			2521 => "0000000010011101111001",
			2522 => "0000010101011100000100",
			2523 => "0000000010011101111001",
			2524 => "0000000010011101111001",
			2525 => "0000000010011101111001",
			2526 => "0000011001111000011000",
			2527 => "0011010100011000000100",
			2528 => "1111111010011111111101",
			2529 => "0001010111001000000100",
			2530 => "0000100010011111111101",
			2531 => "0001110110000100001100",
			2532 => "0011010011100000000100",
			2533 => "0000000010011111111101",
			2534 => "0011011011000000000100",
			2535 => "0000000010011111111101",
			2536 => "0000000010011111111101",
			2537 => "1111111010011111111101",
			2538 => "0010100110011000000100",
			2539 => "1111111010011111111101",
			2540 => "0001100101010000100100",
			2541 => "0001010011100000001000",
			2542 => "0011100101101100000100",
			2543 => "0000000010011111111101",
			2544 => "1111111010011111111101",
			2545 => "0000100110010000001100",
			2546 => "0011100001101000001000",
			2547 => "0000000000111000000100",
			2548 => "0000000010011111111101",
			2549 => "0000001010011111111101",
			2550 => "0000011010011111111101",
			2551 => "0001101011001100001000",
			2552 => "0000011101101000000100",
			2553 => "0000001010011111111101",
			2554 => "1111111010011111111101",
			2555 => "0000101000001100000100",
			2556 => "1111111010011111111101",
			2557 => "0000001010011111111101",
			2558 => "1111111010011111111101",
			2559 => "0001111001110000001000",
			2560 => "0010100110001000000100",
			2561 => "1111111010100010010001",
			2562 => "0000000010100010010001",
			2563 => "0000100111111100010000",
			2564 => "0000101001010000000100",
			2565 => "0000000010100010010001",
			2566 => "0001000010111000000100",
			2567 => "0000000010100010010001",
			2568 => "0001111110001100000100",
			2569 => "0000001010100010010001",
			2570 => "0000000010100010010001",
			2571 => "0001001011001000001100",
			2572 => "0000101110100100000100",
			2573 => "1111111010100010010001",
			2574 => "0000111111101000000100",
			2575 => "0000000010100010010001",
			2576 => "0000000010100010010001",
			2577 => "0000001100001000010000",
			2578 => "0000111001011100001100",
			2579 => "0001111010111100001000",
			2580 => "0011001101111000000100",
			2581 => "0000001010100010010001",
			2582 => "0000000010100010010001",
			2583 => "0000000010100010010001",
			2584 => "0000000010100010010001",
			2585 => "0001001101000000001000",
			2586 => "0010010100110100000100",
			2587 => "0000000010100010010001",
			2588 => "0000000010100010010001",
			2589 => "0011101110110000001000",
			2590 => "0011000110000100000100",
			2591 => "0000000010100010010001",
			2592 => "0000000010100010010001",
			2593 => "0000111100010000000100",
			2594 => "0000000010100010010001",
			2595 => "0000000010100010010001",
			2596 => "0001000000010100000100",
			2597 => "1111111010100100011101",
			2598 => "0010000111000100101000",
			2599 => "0000001110111100011000",
			2600 => "0001101011001100001000",
			2601 => "0010110000001100000100",
			2602 => "0000000010100100011101",
			2603 => "0000000010100100011101",
			2604 => "0010110011100000000100",
			2605 => "0000000010100100011101",
			2606 => "0010101010110000001000",
			2607 => "0011101101101100000100",
			2608 => "0000000010100100011101",
			2609 => "0000000010100100011101",
			2610 => "0000000010100100011101",
			2611 => "0010001111001000000100",
			2612 => "0000000010100100011101",
			2613 => "0000000111111000001000",
			2614 => "0000111010111100000100",
			2615 => "0000000010100100011101",
			2616 => "0000001010100100011101",
			2617 => "0000000010100100011101",
			2618 => "0001100100111100011000",
			2619 => "0001011001110100001000",
			2620 => "0000001110001100000100",
			2621 => "0000000010100100011101",
			2622 => "0000000010100100011101",
			2623 => "0001101011001100000100",
			2624 => "0000000010100100011101",
			2625 => "0010101100011100000100",
			2626 => "0000000010100100011101",
			2627 => "0001000001100100000100",
			2628 => "0000000010100100011101",
			2629 => "0000001010100100011101",
			2630 => "1111111010100100011101",
			2631 => "0001000011010100011100",
			2632 => "0001101011001100000100",
			2633 => "1111111010100111011001",
			2634 => "0001101011001100001100",
			2635 => "0010010001000100000100",
			2636 => "0000000010100111011001",
			2637 => "0011010000110100000100",
			2638 => "0000011010100111011001",
			2639 => "0000000010100111011001",
			2640 => "0010011101011000001000",
			2641 => "0000011111001100000100",
			2642 => "1111111010100111011001",
			2643 => "0000001010100111011001",
			2644 => "1111111010100111011001",
			2645 => "0000011001111000011100",
			2646 => "0000000111111000001000",
			2647 => "0000000111111000000100",
			2648 => "0000000010100111011001",
			2649 => "0000010010100111011001",
			2650 => "0010011101101000000100",
			2651 => "1111111010100111011001",
			2652 => "0000010010001100001100",
			2653 => "0000010010001100001000",
			2654 => "0010011101101000000100",
			2655 => "0000000010100111011001",
			2656 => "0000000010100111011001",
			2657 => "0000000010100111011001",
			2658 => "1111111010100111011001",
			2659 => "0001100101010000100100",
			2660 => "0000111010011100001000",
			2661 => "0001010011100000000100",
			2662 => "0000000010100111011001",
			2663 => "0000001010100111011001",
			2664 => "0001101011001100001100",
			2665 => "0011001100110000000100",
			2666 => "0000000010100111011001",
			2667 => "0011001110001100000100",
			2668 => "1111111010100111011001",
			2669 => "0000000010100111011001",
			2670 => "0000010111100100001000",
			2671 => "0001000000000000000100",
			2672 => "1111111010100111011001",
			2673 => "0000000010100111011001",
			2674 => "0000011101011100000100",
			2675 => "0000001010100111011001",
			2676 => "0000000010100111011001",
			2677 => "1111111010100111011001",
			2678 => "0010110101101100000100",
			2679 => "1111111010101001100101",
			2680 => "0011111010010100001100",
			2681 => "0011110010001000000100",
			2682 => "0000000010101001100101",
			2683 => "0001001110111000000100",
			2684 => "0000000010101001100101",
			2685 => "0000001010101001100101",
			2686 => "0010010100110100011000",
			2687 => "0001001010010000010000",
			2688 => "0011111110101100000100",
			2689 => "0000000010101001100101",
			2690 => "0010011110010100000100",
			2691 => "1111111010101001100101",
			2692 => "0010010100110100000100",
			2693 => "0000000010101001100101",
			2694 => "0000000010101001100101",
			2695 => "0001011011011100000100",
			2696 => "0000000010101001100101",
			2697 => "0000000010101001100101",
			2698 => "0000011001011000010000",
			2699 => "0001101011001100000100",
			2700 => "0000000010101001100101",
			2701 => "0000001011000100001000",
			2702 => "0001010101100100000100",
			2703 => "0000000010101001100101",
			2704 => "0000001010101001100101",
			2705 => "0000000010101001100101",
			2706 => "0000010101011100001100",
			2707 => "0011011001010100000100",
			2708 => "0000000010101001100101",
			2709 => "0001000011010100000100",
			2710 => "0000000010101001100101",
			2711 => "0000000010101001100101",
			2712 => "0000000010101001100101",
			2713 => "0000011001111000000100",
			2714 => "1111111010101100000001",
			2715 => "0011001100110000100000",
			2716 => "0011001000111000001000",
			2717 => "0001001101000000000100",
			2718 => "1111111010101100000001",
			2719 => "0000000010101100000001",
			2720 => "0011000011011100010000",
			2721 => "0000000010111100000100",
			2722 => "0000000010101100000001",
			2723 => "0010100001010000000100",
			2724 => "0000001010101100000001",
			2725 => "0010101100011100000100",
			2726 => "0000000010101100000001",
			2727 => "0000001010101100000001",
			2728 => "0001000010010000000100",
			2729 => "0000000010101100000001",
			2730 => "0000001010101100000001",
			2731 => "0001010000011100010000",
			2732 => "0010001111000100001100",
			2733 => "0011000110000100001000",
			2734 => "0000101111100100000100",
			2735 => "0000000010101100000001",
			2736 => "1111111010101100000001",
			2737 => "0000000010101100000001",
			2738 => "0000000010101100000001",
			2739 => "0001000000010100000100",
			2740 => "1111111010101100000001",
			2741 => "0010101100011100001100",
			2742 => "0000010101011100001000",
			2743 => "0010110011100000000100",
			2744 => "0000000010101100000001",
			2745 => "0000001010101100000001",
			2746 => "0000000010101100000001",
			2747 => "0000000100010100000100",
			2748 => "0000000010101100000001",
			2749 => "0011000100001000000100",
			2750 => "0000000010101100000001",
			2751 => "0000000010101100000001",
			2752 => "0011010100011000000100",
			2753 => "1111111010101110100101",
			2754 => "0011000011011100011100",
			2755 => "0011100100001000001100",
			2756 => "0001001110111000000100",
			2757 => "0000000010101110100101",
			2758 => "0000111001110100000100",
			2759 => "0000001010101110100101",
			2760 => "0000000010101110100101",
			2761 => "0011000011011100001000",
			2762 => "0001001101000000000100",
			2763 => "1111111010101110100101",
			2764 => "0000000010101110100101",
			2765 => "0010010001000100000100",
			2766 => "0000000010101110100101",
			2767 => "0000001010101110100101",
			2768 => "0010110000001100010000",
			2769 => "0010110000001100001000",
			2770 => "0000000011011100000100",
			2771 => "0000000010101110100101",
			2772 => "0000000010101110100101",
			2773 => "0000010110101000000100",
			2774 => "0000000010101110100101",
			2775 => "1111000010101110100101",
			2776 => "0011001010111000100000",
			2777 => "0000011011101000010000",
			2778 => "0010001101010000001000",
			2779 => "0000101011101100000100",
			2780 => "0000000010101110100101",
			2781 => "1111111010101110100101",
			2782 => "0000011001111000000100",
			2783 => "0000000010101110100101",
			2784 => "0000001010101110100101",
			2785 => "0010100110011000001000",
			2786 => "0000101111100100000100",
			2787 => "0000000010101110100101",
			2788 => "0000000010101110100101",
			2789 => "0000100110101100000100",
			2790 => "0000001010101110100101",
			2791 => "0000000010101110100101",
			2792 => "1111111010101110100101",
			2793 => "0001001110111000000100",
			2794 => "1111111010110001010001",
			2795 => "0010000111000100111000",
			2796 => "0010000111000100100000",
			2797 => "0010000110001000011000",
			2798 => "0001000011101100001100",
			2799 => "0011101101101100001000",
			2800 => "0010100110011000000100",
			2801 => "0000000010110001010001",
			2802 => "0000001010110001010001",
			2803 => "0000000010110001010001",
			2804 => "0000101011111000001000",
			2805 => "0011110011001000000100",
			2806 => "0000000010110001010001",
			2807 => "0000000010110001010001",
			2808 => "0000000010110001010001",
			2809 => "0001000000101100000100",
			2810 => "0000000010110001010001",
			2811 => "0000000010110001010001",
			2812 => "0011110101110100001000",
			2813 => "0001000011010100000100",
			2814 => "0000000010110001010001",
			2815 => "0000011010110001010001",
			2816 => "0000011101011100001100",
			2817 => "0001000100001100000100",
			2818 => "0000000010110001010001",
			2819 => "0001010111001000000100",
			2820 => "0000000010110001010001",
			2821 => "0000001010110001010001",
			2822 => "0000000010110001010001",
			2823 => "0001001010010000010000",
			2824 => "0010010100110100000100",
			2825 => "1111111010110001010001",
			2826 => "0000011101011100001000",
			2827 => "0011111110000000000100",
			2828 => "0000000010110001010001",
			2829 => "0000000010110001010001",
			2830 => "0000000010110001010001",
			2831 => "0010011101101000000100",
			2832 => "0000000010110001010001",
			2833 => "0000101110000000000100",
			2834 => "0000000010110001010001",
			2835 => "0000000010110001010001",
			2836 => "0011010100011000000100",
			2837 => "1111111010110011111101",
			2838 => "0011110110010000111100",
			2839 => "0001111101100000011000",
			2840 => "0001101011001100010000",
			2841 => "0000000010111100000100",
			2842 => "0000000010110011111101",
			2843 => "0010101010110000001000",
			2844 => "0001111001110000000100",
			2845 => "0000000010110011111101",
			2846 => "0000001010110011111101",
			2847 => "0000000010110011111101",
			2848 => "0000000100001000000100",
			2849 => "0000000010110011111101",
			2850 => "0000000010110011111101",
			2851 => "0001101011001100010100",
			2852 => "0011001100110000001100",
			2853 => "0000000000111000000100",
			2854 => "0000000010110011111101",
			2855 => "0001010011100000000100",
			2856 => "0000000010110011111101",
			2857 => "0000000010110011111101",
			2858 => "0001101011001100000100",
			2859 => "1111111010110011111101",
			2860 => "0000000010110011111101",
			2861 => "0001001101110100000100",
			2862 => "0000000010110011111101",
			2863 => "0010111000000000001000",
			2864 => "0010000110001000000100",
			2865 => "0000000010110011111101",
			2866 => "0000001010110011111101",
			2867 => "0000000010110011111101",
			2868 => "0001010100010000001000",
			2869 => "0011111001100000000100",
			2870 => "0000000010110011111101",
			2871 => "1111111010110011111101",
			2872 => "0011001010111000001100",
			2873 => "0001000011010100000100",
			2874 => "0000000010110011111101",
			2875 => "0011011110101100000100",
			2876 => "0000000010110011111101",
			2877 => "0000000010110011111101",
			2878 => "0000000010110011111101",
			2879 => "0001111001110000001000",
			2880 => "0010000000111000000100",
			2881 => "0000000010110110011001",
			2882 => "0000000010110110011001",
			2883 => "0001111101100000010100",
			2884 => "0000100110010000010000",
			2885 => "0011101001110000000100",
			2886 => "0000000010110110011001",
			2887 => "0010001001101000000100",
			2888 => "0000000010110110011001",
			2889 => "0011010100011000000100",
			2890 => "0000000010110110011001",
			2891 => "0000001010110110011001",
			2892 => "0000000010110110011001",
			2893 => "0001000000010100000100",
			2894 => "0000000010110110011001",
			2895 => "0000000011111100010000",
			2896 => "0011001110001100000100",
			2897 => "0000000010110110011001",
			2898 => "0000010101011100001000",
			2899 => "0001011011011100000100",
			2900 => "0000000010110110011001",
			2901 => "0000000010110110011001",
			2902 => "0000000010110110011001",
			2903 => "0001101011001100010000",
			2904 => "0011000110000100001000",
			2905 => "0001000001100100000100",
			2906 => "0000000010110110011001",
			2907 => "0000000010110110011001",
			2908 => "0001101011001100000100",
			2909 => "0000000010110110011001",
			2910 => "0000000010110110011001",
			2911 => "0001001101000000001000",
			2912 => "0000111000001100000100",
			2913 => "0000000010110110011001",
			2914 => "0000000010110110011001",
			2915 => "0010001010000000000100",
			2916 => "0000000010110110011001",
			2917 => "0000000010110110011001",
			2918 => "0011010100011000000100",
			2919 => "1111111010111001000101",
			2920 => "0011001100110000101100",
			2921 => "0011001001110000010100",
			2922 => "0011100100001000001100",
			2923 => "0001000111011100000100",
			2924 => "0000000010111001000101",
			2925 => "0001101001100100000100",
			2926 => "0000001010111001000101",
			2927 => "0000000010111001000101",
			2928 => "0001001101000000000100",
			2929 => "1111111010111001000101",
			2930 => "0000000010111001000101",
			2931 => "0000000010111100000100",
			2932 => "0000000010111001000101",
			2933 => "0010100001010000000100",
			2934 => "0000001010111001000101",
			2935 => "0000000111111000001000",
			2936 => "0000001010000000000100",
			2937 => "0000000010111001000101",
			2938 => "0000000010111001000101",
			2939 => "0000011001111000000100",
			2940 => "0000000010111001000101",
			2941 => "0000001010111001000101",
			2942 => "0001101101011000001000",
			2943 => "0011001100110000000100",
			2944 => "0000000010111001000101",
			2945 => "1111111010111001000101",
			2946 => "0000010101011100011100",
			2947 => "0000000000111000001100",
			2948 => "0001010101100100000100",
			2949 => "0000000010111001000101",
			2950 => "0010100110011000000100",
			2951 => "0000000010111001000101",
			2952 => "0000001010111001000101",
			2953 => "0011110111011000001000",
			2954 => "0000001000111100000100",
			2955 => "0000000010111001000101",
			2956 => "0000001010111001000101",
			2957 => "0000011101011100000100",
			2958 => "1111111010111001000101",
			2959 => "0000000010111001000101",
			2960 => "1111111010111001000101",
			2961 => "0011010100011000000100",
			2962 => "1111111010111011010001",
			2963 => "0010001001101000000100",
			2964 => "1111111010111011010001",
			2965 => "0010100001010000011000",
			2966 => "0011001001110000000100",
			2967 => "0000000010111011010001",
			2968 => "0000101011111000001000",
			2969 => "0010001001101000000100",
			2970 => "0000000010111011010001",
			2971 => "0000001010111011010001",
			2972 => "0000110111100000000100",
			2973 => "0000000010111011010001",
			2974 => "0000111111101000000100",
			2975 => "0000001010111011010001",
			2976 => "0000000010111011010001",
			2977 => "0011101101010100010100",
			2978 => "0011000110000100001100",
			2979 => "0001000111011100000100",
			2980 => "0000000010111011010001",
			2981 => "0000011100110100000100",
			2982 => "0000000010111011010001",
			2983 => "0000001010111011010001",
			2984 => "0000011001111000000100",
			2985 => "1111111010111011010001",
			2986 => "0000000010111011010001",
			2987 => "0011011010001100001000",
			2988 => "0001001010101000000100",
			2989 => "1111111010111011010001",
			2990 => "0000000010111011010001",
			2991 => "0011001010111000001000",
			2992 => "0011000000001100000100",
			2993 => "0000000010111011010001",
			2994 => "0000000010111011010001",
			2995 => "1111111010111011010001",
			2996 => "0011010100011000000100",
			2997 => "1111111010111101111101",
			2998 => "0010000111000100110000",
			2999 => "0000000010011000001000",
			3000 => "0001000000010100000100",
			3001 => "0000000010111101111101",
			3002 => "0000000010111101111101",
			3003 => "0000000010111100010000",
			3004 => "0010100001010000001100",
			3005 => "0001011000000000000100",
			3006 => "0000000010111101111101",
			3007 => "0000010101011100000100",
			3008 => "0000001010111101111101",
			3009 => "0000000010111101111101",
			3010 => "0000000010111101111101",
			3011 => "0000001110111100010000",
			3012 => "0010100001010000001000",
			3013 => "0011001110001100000100",
			3014 => "0000000010111101111101",
			3015 => "0000000010111101111101",
			3016 => "0011000000001100000100",
			3017 => "0000000010111101111101",
			3018 => "0000000010111101111101",
			3019 => "0010011101011000000100",
			3020 => "0000001010111101111101",
			3021 => "0000000010111101111101",
			3022 => "0001100100111100100000",
			3023 => "0000011111001100011000",
			3024 => "0010011001011000001100",
			3025 => "0000111110110000000100",
			3026 => "0000000010111101111101",
			3027 => "0000001010111100000100",
			3028 => "0000000010111101111101",
			3029 => "0000000010111101111101",
			3030 => "0001000110110000000100",
			3031 => "0000000010111101111101",
			3032 => "0001101011001100000100",
			3033 => "0000000010111101111101",
			3034 => "0000001010111101111101",
			3035 => "0001101001100100000100",
			3036 => "0000000010111101111101",
			3037 => "0000000010111101111101",
			3038 => "1111111010111101111101",
			3039 => "0010110101101100000100",
			3040 => "1111111011000000001011",
			3041 => "0001000010111000000100",
			3042 => "1111111011000000001011",
			3043 => "0010000111000100011000",
			3044 => "0000010101011100010100",
			3045 => "0000100011001000000100",
			3046 => "0000001011000000001011",
			3047 => "0011010101110100001000",
			3048 => "0000001110111100000100",
			3049 => "1111111011000000001011",
			3050 => "0000000011000000001011",
			3051 => "0011100111110000000100",
			3052 => "0000000011000000001011",
			3053 => "0000001011000000001011",
			3054 => "0000000011000000001011",
			3055 => "0011000110000100010000",
			3056 => "0001000001100100000100",
			3057 => "1111111011000000001011",
			3058 => "0000100010010100001000",
			3059 => "0011001100110000000100",
			3060 => "0000001011000000001011",
			3061 => "0000000011000000001011",
			3062 => "0000000011000000001011",
			3063 => "0011010100000100001100",
			3064 => "0001011010011100001000",
			3065 => "0010111010111100000100",
			3066 => "1111111011000000001011",
			3067 => "0000000011000000001011",
			3068 => "0000000011000000001011",
			3069 => "0011000100001000001000",
			3070 => "0000000100010100000100",
			3071 => "0000000011000000001011",
			3072 => "0000001011000000001011",
			3073 => "0000000011000000001011",
			3074 => "0000000011000000001101",
			3075 => "0000000011000000010001",
			3076 => "0000000011000000010101",
			3077 => "0000000011000000011001",
			3078 => "0000000011000000011101",
			3079 => "0000000011000000100001",
			3080 => "0000000011000000100101",
			3081 => "0000000011000000101001",
			3082 => "0000000011000000101101",
			3083 => "0001001110111000000100",
			3084 => "0000000011000000111001",
			3085 => "0000000011000000111001",
			3086 => "0001101011001100000100",
			3087 => "0000000011000001001101",
			3088 => "0001101000010000000100",
			3089 => "0000000011000001001101",
			3090 => "0000000011000001001101",
			3091 => "0000011011101000000100",
			3092 => "0000000011000001100001",
			3093 => "0000010000111100000100",
			3094 => "0000000011000001100001",
			3095 => "0000000011000001100001",
			3096 => "0000110101110100001000",
			3097 => "0001101001100100000100",
			3098 => "0000000011000001110101",
			3099 => "0000000011000001110101",
			3100 => "0000000011000001110101",
			3101 => "0011101110101100001000",
			3102 => "0001001101000000000100",
			3103 => "0000000011000010001001",
			3104 => "0000000011000010001001",
			3105 => "0000000011000010001001",
			3106 => "0011101100101100000100",
			3107 => "0000000011000010011101",
			3108 => "0011101101101100000100",
			3109 => "0000000011000010011101",
			3110 => "0000000011000010011101",
			3111 => "0011110110010000001000",
			3112 => "0011110010001000000100",
			3113 => "0000000011000010111001",
			3114 => "0000000011000010111001",
			3115 => "0011111011110000000100",
			3116 => "0000000011000010111001",
			3117 => "0000000011000010111001",
			3118 => "0000100100101000000100",
			3119 => "0000000011000011010101",
			3120 => "0011101010000100001000",
			3121 => "0000000100010100000100",
			3122 => "0000000011000011010101",
			3123 => "0000000011000011010101",
			3124 => "0000000011000011010101",
			3125 => "0000100100101000000100",
			3126 => "0000000011000011110001",
			3127 => "0001000011011000001000",
			3128 => "0011111011110000000100",
			3129 => "0000000011000011110001",
			3130 => "0000000011000011110001",
			3131 => "0000000011000011110001",
			3132 => "0000011101011100001100",
			3133 => "0000011100110100000100",
			3134 => "0000000011000100001101",
			3135 => "0000011111001100000100",
			3136 => "0000000011000100001101",
			3137 => "0000000011000100001101",
			3138 => "0000000011000100001101",
			3139 => "0000110010001000000100",
			3140 => "0000000011000100101001",
			3141 => "0010010100111100001000",
			3142 => "0010010001000100000100",
			3143 => "0000000011000100101001",
			3144 => "0000000011000100101001",
			3145 => "0000000011000100101001",
			3146 => "0011001100110000001000",
			3147 => "0011010110100100000100",
			3148 => "0000000011000101001101",
			3149 => "0000000011000101001101",
			3150 => "0011111011110000001000",
			3151 => "0001110110000100000100",
			3152 => "0000000011000101001101",
			3153 => "0000000011000101001101",
			3154 => "0000000011000101001101",
			3155 => "0011110010000000001000",
			3156 => "0011110010001000000100",
			3157 => "0000000011000101110001",
			3158 => "0000000011000101110001",
			3159 => "0011111000110100001000",
			3160 => "0011110110010000000100",
			3161 => "0000000011000101110001",
			3162 => "0000000011000101110001",
			3163 => "0000000011000101110001",
			3164 => "0011000011011100001100",
			3165 => "0001111001110000000100",
			3166 => "0000000011000110011101",
			3167 => "0010111100110000000100",
			3168 => "0000000011000110011101",
			3169 => "0000000011000110011101",
			3170 => "0000110011000000001000",
			3171 => "0001110110000100000100",
			3172 => "0000000011000110011101",
			3173 => "0000000011000110011101",
			3174 => "0000000011000110011101",
			3175 => "0001001100111100001100",
			3176 => "0000100100101000000100",
			3177 => "0000000011000111001001",
			3178 => "0000101110100100000100",
			3179 => "0000000011000111001001",
			3180 => "0000000011000111001001",
			3181 => "0011010001011000000100",
			3182 => "0000000011000111001001",
			3183 => "0011011001010000000100",
			3184 => "0000000011000111001001",
			3185 => "0000000011000111001001",
			3186 => "0000100100101000000100",
			3187 => "0000000011000111101101",
			3188 => "0001000010010000001100",
			3189 => "0011111011110000001000",
			3190 => "0011110101110100000100",
			3191 => "0000000011000111101101",
			3192 => "0000000011000111101101",
			3193 => "0000000011000111101101",
			3194 => "0000000011000111101101",
			3195 => "0011001100110000010000",
			3196 => "0000011100110100000100",
			3197 => "0000000011001000010001",
			3198 => "0000011111001100001000",
			3199 => "0011000000101000000100",
			3200 => "0000000011001000010001",
			3201 => "0000000011001000010001",
			3202 => "0000000011001000010001",
			3203 => "0000000011001000010001",
			3204 => "0001011011011100010000",
			3205 => "0001001010010000001100",
			3206 => "0000101010001000000100",
			3207 => "0000000011001000110101",
			3208 => "0011110101110100000100",
			3209 => "0000000011001000110101",
			3210 => "0000000011001000110101",
			3211 => "0000000011001000110101",
			3212 => "0000000011001000110101",
			3213 => "0000001110111100001000",
			3214 => "0000000010111100000100",
			3215 => "0000000011001001100001",
			3216 => "0000000011001001100001",
			3217 => "0010000001110100001100",
			3218 => "0001111001110000000100",
			3219 => "0000000011001001100001",
			3220 => "0001111101010100000100",
			3221 => "0000000011001001100001",
			3222 => "0000000011001001100001",
			3223 => "0000000011001001100001",
			3224 => "0000001110111100001100",
			3225 => "0000000010111100000100",
			3226 => "0000000011001010010101",
			3227 => "0001000000100000000100",
			3228 => "0000000011001010010101",
			3229 => "0000000011001010010101",
			3230 => "0010000001110100001100",
			3231 => "0001111001110000000100",
			3232 => "0000000011001010010101",
			3233 => "0001111101010100000100",
			3234 => "0000000011001010010101",
			3235 => "0000000011001010010101",
			3236 => "0000000011001010010101",
			3237 => "0000000011111100001100",
			3238 => "0010100110011000000100",
			3239 => "0000000011001011001001",
			3240 => "0010100001010000000100",
			3241 => "0000000011001011001001",
			3242 => "0000000011001011001001",
			3243 => "0010100110011000000100",
			3244 => "0000000011001011001001",
			3245 => "0000001010111100001000",
			3246 => "0011000000001100000100",
			3247 => "0000000011001011001001",
			3248 => "0000000011001011001001",
			3249 => "0000000011001011001001",
			3250 => "0001011011011100010000",
			3251 => "0001001010010000001100",
			3252 => "0000101010001000000100",
			3253 => "0000000011001011111101",
			3254 => "0011110101110100000100",
			3255 => "0000000011001011111101",
			3256 => "0000000011001011111101",
			3257 => "0000000011001011111101",
			3258 => "0011001010111000001000",
			3259 => "0011001110001100000100",
			3260 => "0000000011001011111101",
			3261 => "0000000011001011111101",
			3262 => "0000000011001011111101",
			3263 => "0001000001100100010000",
			3264 => "0010100001010000000100",
			3265 => "0000000011001100111001",
			3266 => "0011110101110100000100",
			3267 => "0000000011001100111001",
			3268 => "0000000010011000000100",
			3269 => "0000000011001100111001",
			3270 => "0000000011001100111001",
			3271 => "0000011111001100001100",
			3272 => "0000010010001100000100",
			3273 => "0000000011001100111001",
			3274 => "0011111000001100000100",
			3275 => "0000000011001100111001",
			3276 => "0000000011001100111001",
			3277 => "0000000011001100111001",
			3278 => "0000011101011100010100",
			3279 => "0000011100110100000100",
			3280 => "0000000011001101100101",
			3281 => "0000000010111100000100",
			3282 => "0000000011001101100101",
			3283 => "0010100001110000001000",
			3284 => "0010101001000100000100",
			3285 => "0000000011001101100101",
			3286 => "0000000011001101100101",
			3287 => "0000000011001101100101",
			3288 => "0000000011001101100101",
			3289 => "0001101101011000001000",
			3290 => "0001001110111000000100",
			3291 => "0000000011001110100001",
			3292 => "0000000011001110100001",
			3293 => "0001101001100100010000",
			3294 => "0000010111100100000100",
			3295 => "0000000011001110100001",
			3296 => "0000010000111100001000",
			3297 => "0001001000000100000100",
			3298 => "0000000011001110100001",
			3299 => "0000000011001110100001",
			3300 => "0000000011001110100001",
			3301 => "0001000011111000000100",
			3302 => "0000000011001110100001",
			3303 => "0000000011001110100001",
			3304 => "0010010100110100011100",
			3305 => "0000101110010000001100",
			3306 => "0000110011100000000100",
			3307 => "0000000011001111101101",
			3308 => "0011100011100000000100",
			3309 => "0000000011001111101101",
			3310 => "0000000011001111101101",
			3311 => "0001001010010000001100",
			3312 => "0011110111110000000100",
			3313 => "0000000011001111101101",
			3314 => "0001010100010000000100",
			3315 => "0000000011001111101101",
			3316 => "0000000011001111101101",
			3317 => "0000000011001111101101",
			3318 => "0000011001011000001000",
			3319 => "0010011010011000000100",
			3320 => "0000000011001111101101",
			3321 => "0000000011001111101101",
			3322 => "0000000011001111101101",
			3323 => "0011001100110000011000",
			3324 => "0011000100000000000100",
			3325 => "0000000011010000110001",
			3326 => "0001001000000100000100",
			3327 => "0000000011010000110001",
			3328 => "0000110100011000000100",
			3329 => "0000000011010000110001",
			3330 => "0000100010010100001000",
			3331 => "0000111001011100000100",
			3332 => "0000000011010000110001",
			3333 => "0000000011010000110001",
			3334 => "0000000011010000110001",
			3335 => "0000100011000000001000",
			3336 => "0000100110101100000100",
			3337 => "0000000011010000110001",
			3338 => "0000000011010000110001",
			3339 => "0000000011010000110001",
			3340 => "0010010001000100001100",
			3341 => "0011111010010100000100",
			3342 => "0000000011010001111101",
			3343 => "0010000010011000000100",
			3344 => "0000000011010001111101",
			3345 => "0000000011010001111101",
			3346 => "0001101000010000010100",
			3347 => "0010100110011000000100",
			3348 => "0000000011010001111101",
			3349 => "0001101011001100000100",
			3350 => "0000000011010001111101",
			3351 => "0010011101011000001000",
			3352 => "0011000011011100000100",
			3353 => "0000000011010001111101",
			3354 => "0000000011010001111101",
			3355 => "0000000011010001111101",
			3356 => "0010100001010000000100",
			3357 => "0000000011010001111101",
			3358 => "0000000011010001111101",
			3359 => "0010011101101000000100",
			3360 => "0000000011010010110001",
			3361 => "0001001110111000000100",
			3362 => "0000000011010010110001",
			3363 => "0010010101010000010000",
			3364 => "0001000100111000001100",
			3365 => "0000110010010100001000",
			3366 => "0010110101101100000100",
			3367 => "0000000011010010110001",
			3368 => "0000000011010010110001",
			3369 => "0000000011010010110001",
			3370 => "0000000011010010110001",
			3371 => "0000000011010010110001",
			3372 => "0000000010111100011000",
			3373 => "0010001001101000000100",
			3374 => "0000000011010011111101",
			3375 => "0000010101011100010000",
			3376 => "0011011001110100000100",
			3377 => "0000000011010011111101",
			3378 => "0010001011010100001000",
			3379 => "0001001000000100000100",
			3380 => "0000000011010011111101",
			3381 => "0000000011010011111101",
			3382 => "0000000011010011111101",
			3383 => "0000000011010011111101",
			3384 => "0000011011101000001100",
			3385 => "0001001010010000001000",
			3386 => "0011110010110100000100",
			3387 => "0000000011010011111101",
			3388 => "0000000011010011111101",
			3389 => "0000000011010011111101",
			3390 => "0000000011010011111101",
			3391 => "0001000011101100001100",
			3392 => "0000100010011100000100",
			3393 => "0000000011010101010001",
			3394 => "0001110111010000000100",
			3395 => "0000000011010101010001",
			3396 => "0000000011010101010001",
			3397 => "0010000010101000010100",
			3398 => "0000010000111100010000",
			3399 => "0000001011000100001100",
			3400 => "0000011100110100000100",
			3401 => "0000000011010101010001",
			3402 => "0010001001101000000100",
			3403 => "0000000011010101010001",
			3404 => "0000000011010101010001",
			3405 => "0000000011010101010001",
			3406 => "0000000011010101010001",
			3407 => "0001001101000000000100",
			3408 => "0000000011010101010001",
			3409 => "0001001111110000000100",
			3410 => "0000000011010101010001",
			3411 => "0000000011010101010001",
			3412 => "0001000011101100001100",
			3413 => "0000100010011100000100",
			3414 => "0000000011010110100101",
			3415 => "0001101000010000000100",
			3416 => "0000000011010110100101",
			3417 => "0000000011010110100101",
			3418 => "0001100100111100011100",
			3419 => "0011010101100100010000",
			3420 => "0011111111010000001000",
			3421 => "0000111110001100000100",
			3422 => "0000000011010110100101",
			3423 => "0000000011010110100101",
			3424 => "0011101101010100000100",
			3425 => "0000000011010110100101",
			3426 => "0000000011010110100101",
			3427 => "0011000100001000001000",
			3428 => "0010001001101000000100",
			3429 => "0000000011010110100101",
			3430 => "0000000011010110100101",
			3431 => "0000000011010110100101",
			3432 => "0000000011010110100101",
			3433 => "0010000111000100011100",
			3434 => "0010110101101100000100",
			3435 => "0000000011010111110001",
			3436 => "0010001001101000000100",
			3437 => "0000000011010111110001",
			3438 => "0000010101011100010000",
			3439 => "0010101100011100001100",
			3440 => "0011000100000000000100",
			3441 => "0000000011010111110001",
			3442 => "0001001000000100000100",
			3443 => "0000000011010111110001",
			3444 => "0000000011010111110001",
			3445 => "0000000011010111110001",
			3446 => "0000000011010111110001",
			3447 => "0001001010010000001000",
			3448 => "0010111000011000000100",
			3449 => "0000000011010111110001",
			3450 => "0000000011010111110001",
			3451 => "0000000011010111110001",
			3452 => "0001111100101000011100",
			3453 => "0010110101101100000100",
			3454 => "0000000011011000111101",
			3455 => "0000011111001100010100",
			3456 => "0000000010111100000100",
			3457 => "0000000011011000111101",
			3458 => "0000010010001100000100",
			3459 => "0000000011011000111101",
			3460 => "0000100010010100001000",
			3461 => "0011000100000000000100",
			3462 => "0000000011011000111101",
			3463 => "0000000011011000111101",
			3464 => "0000000011011000111101",
			3465 => "0000000011011000111101",
			3466 => "0000000010111100000100",
			3467 => "0000000011011000111101",
			3468 => "0000101000100000000100",
			3469 => "0000000011011000111101",
			3470 => "0000000011011000111101",
			3471 => "0011110110010000011100",
			3472 => "0001111001110000000100",
			3473 => "0000000011011010000001",
			3474 => "0010001001101000000100",
			3475 => "0000000011011010000001",
			3476 => "0011001100110000010000",
			3477 => "0001111101111000001100",
			3478 => "0010001010000000001000",
			3479 => "0011000000101000000100",
			3480 => "0000000011011010000001",
			3481 => "0000000011011010000001",
			3482 => "0000000011011010000001",
			3483 => "0000000011011010000001",
			3484 => "0000000011011010000001",
			3485 => "0011000011011100000100",
			3486 => "0000000011011010000001",
			3487 => "0000000011011010000001",
			3488 => "0001111100101000011100",
			3489 => "0011010100011000000100",
			3490 => "0000000011011011010101",
			3491 => "0001101000010000010100",
			3492 => "0000000010111100000100",
			3493 => "0000000011011011010101",
			3494 => "0000011100110100000100",
			3495 => "0000000011011011010101",
			3496 => "0010001001101000000100",
			3497 => "0000000011011011010101",
			3498 => "0001111001110000000100",
			3499 => "0000000011011011010101",
			3500 => "0000000011011011010101",
			3501 => "0000000011011011010101",
			3502 => "0011011001010100001100",
			3503 => "0010111110110000000100",
			3504 => "0000000011011011010101",
			3505 => "0000100000010000000100",
			3506 => "0000000011011011010101",
			3507 => "0000000011011011010101",
			3508 => "0000000011011011010101",
			3509 => "0010011010011000100100",
			3510 => "0000101110010000011000",
			3511 => "0000110011100000000100",
			3512 => "0000000011011100101001",
			3513 => "0011100011100000010000",
			3514 => "0010110101101100000100",
			3515 => "0000000011011100101001",
			3516 => "0010111110001100001000",
			3517 => "0011001001110000000100",
			3518 => "0000000011011100101001",
			3519 => "0000000011011100101001",
			3520 => "0000000011011100101001",
			3521 => "0000000011011100101001",
			3522 => "0001001010010000001000",
			3523 => "0011101000111000000100",
			3524 => "0000000011011100101001",
			3525 => "0000000011011100101001",
			3526 => "0000000011011100101001",
			3527 => "0000011001011000000100",
			3528 => "0000000011011100101001",
			3529 => "0000000011011100101001",
			3530 => "0000100110101100011100",
			3531 => "0010011101101000000100",
			3532 => "0000000011011101111101",
			3533 => "0000000010111100000100",
			3534 => "0000000011011101111101",
			3535 => "0010110101101100000100",
			3536 => "0000000011011101111101",
			3537 => "0001101001100100001100",
			3538 => "0001111001110000000100",
			3539 => "0000000011011101111101",
			3540 => "0011010100011000000100",
			3541 => "0000000011011101111101",
			3542 => "0000000011011101111101",
			3543 => "0000000011011101111101",
			3544 => "0011111011110000001100",
			3545 => "0001001010010000001000",
			3546 => "0000000010111100000100",
			3547 => "0000000011011101111101",
			3548 => "0000000011011101111101",
			3549 => "0000000011011101111101",
			3550 => "0000000011011101111101",
			3551 => "0001110001111100011100",
			3552 => "0011010100011000000100",
			3553 => "0000000011011110111001",
			3554 => "0010100110011100010100",
			3555 => "0000000010111100000100",
			3556 => "0000000011011110111001",
			3557 => "0001111001110000000100",
			3558 => "0000000011011110111001",
			3559 => "0011110000010000001000",
			3560 => "0010001001101000000100",
			3561 => "0000000011011110111001",
			3562 => "0000000011011110111001",
			3563 => "0000000011011110111001",
			3564 => "0000000011011110111001",
			3565 => "0000000011011110111001",
			3566 => "0000010110101000000100",
			3567 => "0000000011011111110101",
			3568 => "0000010101011100011000",
			3569 => "0010101001000100000100",
			3570 => "0000000011011111110101",
			3571 => "0001111001110000000100",
			3572 => "0000000011011111110101",
			3573 => "0011011001110100000100",
			3574 => "0000000011011111110101",
			3575 => "0010111011110100001000",
			3576 => "0001011000000000000100",
			3577 => "0000000011011111110101",
			3578 => "0000000011011111110101",
			3579 => "0000000011011111110101",
			3580 => "0000000011011111110101",
			3581 => "0011101100101100000100",
			3582 => "0000000011100000110001",
			3583 => "0011110000010000011000",
			3584 => "0000011101011100010100",
			3585 => "0010101001000100000100",
			3586 => "0000000011100000110001",
			3587 => "0010011101101000000100",
			3588 => "0000000011100000110001",
			3589 => "0010011101011000001000",
			3590 => "0001101000010000000100",
			3591 => "0000000011100000110001",
			3592 => "0000000011100000110001",
			3593 => "0000000011100000110001",
			3594 => "0000000011100000110001",
			3595 => "0000000011100000110001",
			3596 => "0001001110111000000100",
			3597 => "0000000011100010001101",
			3598 => "0010000111000100010000",
			3599 => "0001111001110000000100",
			3600 => "0000000011100010001101",
			3601 => "0000100011110000001000",
			3602 => "0010001001101000000100",
			3603 => "0000000011100010001101",
			3604 => "0000000011100010001101",
			3605 => "0000000011100010001101",
			3606 => "0001100100111100010100",
			3607 => "0001000110110000001000",
			3608 => "0000101100111000000100",
			3609 => "0000000011100010001101",
			3610 => "0000000011100010001101",
			3611 => "0001101011001100000100",
			3612 => "0000000011100010001101",
			3613 => "0000000110100100000100",
			3614 => "0000000011100010001101",
			3615 => "0000000011100010001101",
			3616 => "0011011100100100000100",
			3617 => "0000000011100010001101",
			3618 => "0000000011100010001101",
			3619 => "0000100110101100011100",
			3620 => "0010011101101000000100",
			3621 => "0000000011100011101001",
			3622 => "0000000010111100000100",
			3623 => "0000000011100011101001",
			3624 => "0010110101101100000100",
			3625 => "0000000011100011101001",
			3626 => "0001101001100100001100",
			3627 => "0010001001101000000100",
			3628 => "0000000011100011101001",
			3629 => "0001111001110000000100",
			3630 => "0000000011100011101001",
			3631 => "0000000011100011101001",
			3632 => "0000000011100011101001",
			3633 => "0011001100110000000100",
			3634 => "0000000011100011101001",
			3635 => "0011111011110000001100",
			3636 => "0000000010111100000100",
			3637 => "0000000011100011101001",
			3638 => "0000001010111100000100",
			3639 => "0000000011100011101001",
			3640 => "0000000011100011101001",
			3641 => "0000000011100011101001",
			3642 => "0000000010111100011000",
			3643 => "0010001001101000000100",
			3644 => "0000000011100101011101",
			3645 => "0011001000111000000100",
			3646 => "0000000011100101011101",
			3647 => "0000010101011100001100",
			3648 => "0010001011010100001000",
			3649 => "0001001000000100000100",
			3650 => "0000000011100101011101",
			3651 => "0000001011100101011101",
			3652 => "0000000011100101011101",
			3653 => "0000000011100101011101",
			3654 => "0000100100101000001000",
			3655 => "0000111010111000000100",
			3656 => "0000000011100101011101",
			3657 => "0000000011100101011101",
			3658 => "0001001011001000000100",
			3659 => "1111111011100101011101",
			3660 => "0000100110101100001100",
			3661 => "0001011001001000000100",
			3662 => "0000000011100101011101",
			3663 => "0011101101100000000100",
			3664 => "0000000011100101011101",
			3665 => "0000000011100101011101",
			3666 => "0000001010111100001000",
			3667 => "0001011011011100000100",
			3668 => "0000000011100101011101",
			3669 => "0000000011100101011101",
			3670 => "0000000011100101011101",
			3671 => "0000000010111100011000",
			3672 => "0010001001101000000100",
			3673 => "0000000011100111010001",
			3674 => "0011001000111000000100",
			3675 => "0000000011100111010001",
			3676 => "0000010101011100001100",
			3677 => "0010001011010100001000",
			3678 => "0001001000000100000100",
			3679 => "0000000011100111010001",
			3680 => "0000001011100111010001",
			3681 => "0000000011100111010001",
			3682 => "0000000011100111010001",
			3683 => "0000100100101000001000",
			3684 => "0000111010111000000100",
			3685 => "0000000011100111010001",
			3686 => "0000000011100111010001",
			3687 => "0001001011001000000100",
			3688 => "0000000011100111010001",
			3689 => "0000100110101100001000",
			3690 => "0000010110101000000100",
			3691 => "0000000011100111010001",
			3692 => "0000000011100111010001",
			3693 => "0000001010111100001100",
			3694 => "0001011011011100001000",
			3695 => "0011111110101000000100",
			3696 => "0000000011100111010001",
			3697 => "0000000011100111010001",
			3698 => "0000000011100111010001",
			3699 => "0000000011100111010001",
			3700 => "0000100100101000010000",
			3701 => "0001111001110000000100",
			3702 => "0000000011101001010101",
			3703 => "0011101001110000000100",
			3704 => "0000000011101001010101",
			3705 => "0010001001101000000100",
			3706 => "0000000011101001010101",
			3707 => "0000000011101001010101",
			3708 => "0000000010111100011000",
			3709 => "0010100110011000000100",
			3710 => "0000000011101001010101",
			3711 => "0000010101011100010000",
			3712 => "0000110101110100000100",
			3713 => "0000000011101001010101",
			3714 => "0010001011010100001000",
			3715 => "0001001000000100000100",
			3716 => "0000000011101001010101",
			3717 => "0000000011101001010101",
			3718 => "0000000011101001010101",
			3719 => "0000000011101001010101",
			3720 => "0001001101000000001100",
			3721 => "0010110100011000001000",
			3722 => "0000100111111100000100",
			3723 => "0000000011101001010101",
			3724 => "0000000011101001010101",
			3725 => "0000000011101001010101",
			3726 => "0010100111000100001100",
			3727 => "0010111001110100001000",
			3728 => "0001101010011000000100",
			3729 => "0000000011101001010101",
			3730 => "0000000011101001010101",
			3731 => "0000000011101001010101",
			3732 => "0000000011101001010101",
			3733 => "0001001110111000000100",
			3734 => "0000000011101010111001",
			3735 => "0010000111000100011000",
			3736 => "0000010101011100010100",
			3737 => "0000011100110100000100",
			3738 => "0000000011101010111001",
			3739 => "0010101100011100001100",
			3740 => "0010100110011000000100",
			3741 => "0000000011101010111001",
			3742 => "0011010100011000000100",
			3743 => "0000000011101010111001",
			3744 => "0000000011101010111001",
			3745 => "0000000011101010111001",
			3746 => "0000000011101010111001",
			3747 => "0001100100111100010000",
			3748 => "0001101011001100000100",
			3749 => "0000000011101010111001",
			3750 => "0001000110110000000100",
			3751 => "0000000011101010111001",
			3752 => "0000010010001100000100",
			3753 => "0000000011101010111001",
			3754 => "0000000011101010111001",
			3755 => "0011011100100100000100",
			3756 => "0000000011101010111001",
			3757 => "0000000011101010111001",
			3758 => "0011110110010000110100",
			3759 => "0001111001110000001000",
			3760 => "0010100110001000000100",
			3761 => "0000000011101100111101",
			3762 => "0000000011101100111101",
			3763 => "0001111101100000010100",
			3764 => "0000100110010000010000",
			3765 => "0010100110011000000100",
			3766 => "0000000011101100111101",
			3767 => "0011010100011000000100",
			3768 => "0000000011101100111101",
			3769 => "0001101011001100000100",
			3770 => "0000000011101100111101",
			3771 => "0000000011101100111101",
			3772 => "0000000011101100111101",
			3773 => "0001001011001000001000",
			3774 => "0000101010001000000100",
			3775 => "0000000011101100111101",
			3776 => "0000000011101100111101",
			3777 => "0000011001111000000100",
			3778 => "0000000011101100111101",
			3779 => "0001101101011000000100",
			3780 => "0000000011101100111101",
			3781 => "0001110111001000000100",
			3782 => "0000000011101100111101",
			3783 => "0000000011101100111101",
			3784 => "0010011010011000001000",
			3785 => "0011111001100000000100",
			3786 => "0000000011101100111101",
			3787 => "0000000011101100111101",
			3788 => "0000011001011000000100",
			3789 => "0000000011101100111101",
			3790 => "0000000011101100111101",
			3791 => "0000011011101000011100",
			3792 => "0011110100101000011000",
			3793 => "0011010100011000000100",
			3794 => "0000000011101110101001",
			3795 => "0011000110000100010000",
			3796 => "0010100110011000000100",
			3797 => "0000000011101110101001",
			3798 => "0001101111000000001000",
			3799 => "0000111110001100000100",
			3800 => "0000000011101110101001",
			3801 => "0000000011101110101001",
			3802 => "0000000011101110101001",
			3803 => "0000000011101110101001",
			3804 => "0000000011101110101001",
			3805 => "0010100110011000000100",
			3806 => "0000000011101110101001",
			3807 => "0000010101011100010100",
			3808 => "0011011011011100000100",
			3809 => "0000000011101110101001",
			3810 => "0000100011110000001100",
			3811 => "0001100101010000001000",
			3812 => "0001000000010100000100",
			3813 => "0000000011101110101001",
			3814 => "0000000011101110101001",
			3815 => "0000000011101110101001",
			3816 => "0000000011101110101001",
			3817 => "0000000011101110101001",
			3818 => "0001010100011000001000",
			3819 => "0001001101000000000100",
			3820 => "1111111011110000011101",
			3821 => "0000000011110000011101",
			3822 => "0011000011011100010000",
			3823 => "0011001000111000000100",
			3824 => "0000000011110000011101",
			3825 => "0011110000010000001000",
			3826 => "0010001001101000000100",
			3827 => "0000000011110000011101",
			3828 => "0000001011110000011101",
			3829 => "0000000011110000011101",
			3830 => "0010100110011000000100",
			3831 => "0000000011110000011101",
			3832 => "0001111101111000010000",
			3833 => "0010101100000100001100",
			3834 => "0001101101011000000100",
			3835 => "0000000011110000011101",
			3836 => "0010010001111000000100",
			3837 => "0000000011110000011101",
			3838 => "0000000011110000011101",
			3839 => "0000000011110000011101",
			3840 => "0000111111101000001100",
			3841 => "0001101101011000000100",
			3842 => "0000000011110000011101",
			3843 => "0010010001000100000100",
			3844 => "0000000011110000011101",
			3845 => "0000000011110000011101",
			3846 => "0000000011110000011101",
			3847 => "0011010100011000000100",
			3848 => "1111111011110010000001",
			3849 => "0011000100001000100000",
			3850 => "0001101000010000011100",
			3851 => "0000000010011000000100",
			3852 => "1111111011110010000001",
			3853 => "0000101110010000001000",
			3854 => "0010111110001100000100",
			3855 => "0000010011110010000001",
			3856 => "0000000011110010000001",
			3857 => "0010111110001100001000",
			3858 => "0000110011100000000100",
			3859 => "0000000011110010000001",
			3860 => "1111111011110010000001",
			3861 => "0011001100110000000100",
			3862 => "0000001011110010000001",
			3863 => "0000000011110010000001",
			3864 => "1111111011110010000001",
			3865 => "0000100101000000000100",
			3866 => "1111111011110010000001",
			3867 => "0011110101000000001000",
			3868 => "0000000010111100000100",
			3869 => "0000001011110010000001",
			3870 => "0000000011110010000001",
			3871 => "1111111011110010000001",
			3872 => "0011010100011000000100",
			3873 => "1111111011110011111101",
			3874 => "0001111100101000101100",
			3875 => "0010000111000100010100",
			3876 => "0000000010111100000100",
			3877 => "0000000011110011111101",
			3878 => "0001111001110000000100",
			3879 => "0000000011110011111101",
			3880 => "0011001110001100001000",
			3881 => "0011101110010000000100",
			3882 => "0000001011110011111101",
			3883 => "0000000011110011111101",
			3884 => "0000000011110011111101",
			3885 => "0001001101000000001100",
			3886 => "0011000011011100001000",
			3887 => "0001101101011000000100",
			3888 => "0000000011110011111101",
			3889 => "0000000011110011111101",
			3890 => "0000000011110011111101",
			3891 => "0001101101011000000100",
			3892 => "0000000011110011111101",
			3893 => "0000000001001000000100",
			3894 => "0000000011110011111101",
			3895 => "0000000011110011111101",
			3896 => "0000101000100000001000",
			3897 => "0011001110001100000100",
			3898 => "0000000011110011111101",
			3899 => "0000000011110011111101",
			3900 => "0011101010111000000100",
			3901 => "0000000011110011111101",
			3902 => "0000000011110011111101",
			3903 => "0001010100011000001000",
			3904 => "0001001101000000000100",
			3905 => "1111111011110110001001",
			3906 => "0000000011110110001001",
			3907 => "0000100110010000010000",
			3908 => "0010111110001100001100",
			3909 => "0011000011011100001000",
			3910 => "0000000010111100000100",
			3911 => "0000000011110110001001",
			3912 => "0000001011110110001001",
			3913 => "0000000011110110001001",
			3914 => "0000000011110110001001",
			3915 => "0001111101111000010000",
			3916 => "0000001100101100001100",
			3917 => "0011111101000100000100",
			3918 => "0000000011110110001001",
			3919 => "0010010001111000000100",
			3920 => "0000000011110110001001",
			3921 => "0000000011110110001001",
			3922 => "0000000011110110001001",
			3923 => "0001001100111100010000",
			3924 => "0000101110100100001000",
			3925 => "0000101011111000000100",
			3926 => "0000000011110110001001",
			3927 => "0000000011110110001001",
			3928 => "0000111111101000000100",
			3929 => "0000000011110110001001",
			3930 => "0000000011110110001001",
			3931 => "0001110111001000001100",
			3932 => "0001101101011000000100",
			3933 => "0000000011110110001001",
			3934 => "0010000110001000000100",
			3935 => "0000000011110110001001",
			3936 => "0000000011110110001001",
			3937 => "0000000011110110001001",
			3938 => "0001101101011000011100",
			3939 => "0010011011101000001000",
			3940 => "0011110101110000000100",
			3941 => "1111111011111000111101",
			3942 => "1111110011111000111101",
			3943 => "0011110010110100001100",
			3944 => "0010001001101000000100",
			3945 => "1111111011111000111101",
			3946 => "0001010011100000000100",
			3947 => "1111111011111000111101",
			3948 => "0000011011111000111101",
			3949 => "0000111110110000000100",
			3950 => "0000000011111000111101",
			3951 => "1111111011111000111101",
			3952 => "0011000100001000110000",
			3953 => "0000100000010000010100",
			3954 => "0010111110001100000100",
			3955 => "1111111011111000111101",
			3956 => "0001111001110000000100",
			3957 => "0000100011111000111101",
			3958 => "0000001100110000000100",
			3959 => "1111111011111000111101",
			3960 => "0011100110001000000100",
			3961 => "0000000011111000111101",
			3962 => "0000001011111000111101",
			3963 => "0001101000010000011000",
			3964 => "0011111010000100010000",
			3965 => "0011110110010000001000",
			3966 => "0011100100010000000100",
			3967 => "0000001011111000111101",
			3968 => "0000010011111000111101",
			3969 => "0010010100111100000100",
			3970 => "0000000011111000111101",
			3971 => "1111111011111000111101",
			3972 => "0000000010111100000100",
			3973 => "0000000011111000111101",
			3974 => "0000010011111000111101",
			3975 => "1111111011111000111101",
			3976 => "0011101101101100001100",
			3977 => "0000110011000000000100",
			3978 => "1111111011111000111101",
			3979 => "0000111111101000000100",
			3980 => "0000001011111000111101",
			3981 => "1111111011111000111101",
			3982 => "1111111011111000111101",
			3983 => "0011010100011000000100",
			3984 => "1111111011111011000001",
			3985 => "0001111100101000110000",
			3986 => "0010000111000100011000",
			3987 => "0000000010111100000100",
			3988 => "0000000011111011000001",
			3989 => "0001111001110000000100",
			3990 => "0000000011111011000001",
			3991 => "0001111101100000001000",
			3992 => "0001101011001100000100",
			3993 => "0000001011111011000001",
			3994 => "0000000011111011000001",
			3995 => "0000110010110100000100",
			3996 => "0000000011111011000001",
			3997 => "0000000011111011000001",
			3998 => "0000010110101000001100",
			3999 => "0011111110101000000100",
			4000 => "0000000011111011000001",
			4001 => "0000001100101100000100",
			4002 => "0000000011111011000001",
			4003 => "0000000011111011000001",
			4004 => "0000000100000000000100",
			4005 => "0000000011111011000001",
			4006 => "0010100110001000000100",
			4007 => "0000000011111011000001",
			4008 => "0000000011111011000001",
			4009 => "0000101000100000001000",
			4010 => "0011001110001100000100",
			4011 => "0000000011111011000001",
			4012 => "0000000011111011000001",
			4013 => "0010111110110000000100",
			4014 => "0000000011111011000001",
			4015 => "0000000011111011000001",
			4016 => "0010011101101000000100",
			4017 => "0000000011111100111101",
			4018 => "0000100110010000011000",
			4019 => "0010110101101100000100",
			4020 => "0000000011111100111101",
			4021 => "0011001100110000010000",
			4022 => "0010001001101000000100",
			4023 => "0000000011111100111101",
			4024 => "0001111001110000000100",
			4025 => "0000000011111100111101",
			4026 => "0001101011001100000100",
			4027 => "0000001011111100111101",
			4028 => "0000000011111100111101",
			4029 => "0000000011111100111101",
			4030 => "0000011011101000001000",
			4031 => "0011101010001100000100",
			4032 => "0000000011111100111101",
			4033 => "0000000011111100111101",
			4034 => "0011011011011100001000",
			4035 => "0001101111000000000100",
			4036 => "0000000011111100111101",
			4037 => "0000000011111100111101",
			4038 => "0011000100001000001100",
			4039 => "0010001011010100000100",
			4040 => "0000000011111100111101",
			4041 => "0000010000111100000100",
			4042 => "0000000011111100111101",
			4043 => "0000000011111100111101",
			4044 => "0001101000010000000100",
			4045 => "0000000011111100111101",
			4046 => "0000000011111100111101",
			4047 => "0001001001000000100100",
			4048 => "0001001110111000000100",
			4049 => "1111111011111111110001",
			4050 => "0010000110001000010100",
			4051 => "0000000011010000001100",
			4052 => "0000010101011100001000",
			4053 => "0001111101010100000100",
			4054 => "1111111011111111110001",
			4055 => "0000001011111111110001",
			4056 => "1111111011111111110001",
			4057 => "0011101011000100000100",
			4058 => "0000000011111111110001",
			4059 => "0000011011111111110001",
			4060 => "0010110101101100000100",
			4061 => "1111111011111111110001",
			4062 => "0001011010111000000100",
			4063 => "0000001011111111110001",
			4064 => "1111111011111111110001",
			4065 => "0010011011101000010000",
			4066 => "0011110101001000001100",
			4067 => "0010011101101000000100",
			4068 => "1111111011111111110001",
			4069 => "0011100110000100000100",
			4070 => "0000001011111111110001",
			4071 => "0000000011111111110001",
			4072 => "1111111011111111110001",
			4073 => "0001110011100000100100",
			4074 => "0000001100001000010100",
			4075 => "0010001011010100001000",
			4076 => "0001111101010100000100",
			4077 => "1111111011111111110001",
			4078 => "0000010011111111110001",
			4079 => "0010000010101000001000",
			4080 => "0000101011111000000100",
			4081 => "0000011011111111110001",
			4082 => "0000001011111111110001",
			4083 => "0000000011111111110001",
			4084 => "0000001000111100000100",
			4085 => "0000000011111111110001",
			4086 => "0001001011100100000100",
			4087 => "1111111011111111110001",
			4088 => "0010100001110000000100",
			4089 => "0000000011111111110001",
			4090 => "0000001011111111110001",
			4091 => "1111111011111111110001",
			4092 => "0011010100011000000100",
			4093 => "1111111100000001110101",
			4094 => "0011110010110100010000",
			4095 => "0011111011011100000100",
			4096 => "0000000100000001110101",
			4097 => "0001000010111000000100",
			4098 => "0000000100000001110101",
			4099 => "0011000110000100000100",
			4100 => "0000001100000001110101",
			4101 => "0000000100000001110101",
			4102 => "0000011011101000001100",
			4103 => "0001001010010000000100",
			4104 => "1111111100000001110101",
			4105 => "0001011011011100000100",
			4106 => "0000000100000001110101",
			4107 => "0000000100000001110101",
			4108 => "0001111100101000001100",
			4109 => "0010111010111000000100",
			4110 => "0000000100000001110101",
			4111 => "0010001011010100000100",
			4112 => "0000000100000001110101",
			4113 => "0000001100000001110101",
			4114 => "0001010101100100001100",
			4115 => "0000101100111000001000",
			4116 => "0011001110001100000100",
			4117 => "1111111100000001110101",
			4118 => "0000000100000001110101",
			4119 => "0000000100000001110101",
			4120 => "0011001010111000001000",
			4121 => "0010100001010000000100",
			4122 => "0000000100000001110101",
			4123 => "0000000100000001110101",
			4124 => "0000000100000001110101",
			4125 => "0001111001110000001000",
			4126 => "0010100110001000000100",
			4127 => "1111111100000100001001",
			4128 => "0000000100000100001001",
			4129 => "0000100111111100010000",
			4130 => "0000101001010000000100",
			4131 => "0000000100000100001001",
			4132 => "0001000010111000000100",
			4133 => "0000000100000100001001",
			4134 => "0001111110001100000100",
			4135 => "0000001100000100001001",
			4136 => "0000000100000100001001",
			4137 => "0001001011001000001100",
			4138 => "0000101110100100000100",
			4139 => "0000000100000100001001",
			4140 => "0000111111101000000100",
			4141 => "0000000100000100001001",
			4142 => "0000000100000100001001",
			4143 => "0000001100001000010000",
			4144 => "0000111001011100001100",
			4145 => "0001111010111100001000",
			4146 => "0011001101111000000100",
			4147 => "0000000100000100001001",
			4148 => "0000000100000100001001",
			4149 => "0000000100000100001001",
			4150 => "0000000100000100001001",
			4151 => "0001001101000000001000",
			4152 => "0010010100110100000100",
			4153 => "0000000100000100001001",
			4154 => "0000000100000100001001",
			4155 => "0011101110110000001000",
			4156 => "0011000110000100000100",
			4157 => "0000000100000100001001",
			4158 => "0000000100000100001001",
			4159 => "0000111100010000000100",
			4160 => "0000000100000100001001",
			4161 => "0000000100000100001001",
			4162 => "0001001001000000100000",
			4163 => "0001001110111000000100",
			4164 => "1111111100000110111101",
			4165 => "0010000110001000010000",
			4166 => "0000110010010100001100",
			4167 => "0010001011010100001000",
			4168 => "0011000000001100000100",
			4169 => "1111111100000110111101",
			4170 => "0000001100000110111101",
			4171 => "0000100100000110111101",
			4172 => "1111111100000110111101",
			4173 => "0011010100011000000100",
			4174 => "1111111100000110111101",
			4175 => "0000111001001000000100",
			4176 => "0000010100000110111101",
			4177 => "1111111100000110111101",
			4178 => "0010011011101000010000",
			4179 => "0011110101001000001100",
			4180 => "0010011101101000000100",
			4181 => "1111111100000110111101",
			4182 => "0011100110000100000100",
			4183 => "0000001100000110111101",
			4184 => "0000000100000110111101",
			4185 => "1111110100000110111101",
			4186 => "0001101000010000101000",
			4187 => "0001000001001100010100",
			4188 => "0000111000011000000100",
			4189 => "0000111100000110111101",
			4190 => "0000111101000100001000",
			4191 => "0000011101011100000100",
			4192 => "0000010100000110111101",
			4193 => "1111111100000110111101",
			4194 => "0001011011011100000100",
			4195 => "0010010100000110111101",
			4196 => "0000011100000110111101",
			4197 => "0001101101011000001000",
			4198 => "0000101011111000000100",
			4199 => "0000001100000110111101",
			4200 => "1111111100000110111101",
			4201 => "0011111100010100001000",
			4202 => "0010100001110000000100",
			4203 => "0000001100000110111101",
			4204 => "0000001100000110111101",
			4205 => "0000001100000110111101",
			4206 => "1111111100000110111101",
			4207 => "0001001001000000110000",
			4208 => "0010110101101100000100",
			4209 => "1111111100001001011001",
			4210 => "0011010110100100011000",
			4211 => "0011011001110100001000",
			4212 => "0010011011101000000100",
			4213 => "0000001100001001011001",
			4214 => "1111111100001001011001",
			4215 => "0000000010111100000100",
			4216 => "0000000100001001011001",
			4217 => "0000000011111100000100",
			4218 => "0001100100001001011001",
			4219 => "0001111101100000000100",
			4220 => "0000000100001001011001",
			4221 => "0000010100001001011001",
			4222 => "0001000000010100000100",
			4223 => "1111111100001001011001",
			4224 => "0000000010011000001100",
			4225 => "0000011011111100001000",
			4226 => "0010001100000100000100",
			4227 => "0000000100001001011001",
			4228 => "0000001100001001011001",
			4229 => "0000000100001001011001",
			4230 => "1111111100001001011001",
			4231 => "0000011100110100000100",
			4232 => "1111111100001001011001",
			4233 => "0001111110110000011000",
			4234 => "0001101000010000010100",
			4235 => "0001111001110000001000",
			4236 => "0011000100000000000100",
			4237 => "1111111100001001011001",
			4238 => "0000000100001001011001",
			4239 => "0000101110110100000100",
			4240 => "0000010100001001011001",
			4241 => "0001101101011000000100",
			4242 => "0000000100001001011001",
			4243 => "0000001100001001011001",
			4244 => "1111111100001001011001",
			4245 => "1111111100001001011001",
			4246 => "0001001001000000011100",
			4247 => "0001001110111000000100",
			4248 => "1111111100001100000101",
			4249 => "0010110101101100000100",
			4250 => "1111111100001100000101",
			4251 => "0000101100010100000100",
			4252 => "0000100100001100000101",
			4253 => "0010101010110000001100",
			4254 => "0000101111100100000100",
			4255 => "1111111100001100000101",
			4256 => "0000110010010100000100",
			4257 => "0000010100001100000101",
			4258 => "1111111100001100000101",
			4259 => "1111111100001100000101",
			4260 => "0010011011101000010000",
			4261 => "0011110101001000001100",
			4262 => "0010011101101000000100",
			4263 => "1111111100001100000101",
			4264 => "0000100111011000000100",
			4265 => "0000000100001100000101",
			4266 => "0000001100001100000101",
			4267 => "1111110100001100000101",
			4268 => "0001101000010000101000",
			4269 => "0000001100001000011000",
			4270 => "0000000011010000001000",
			4271 => "0011110110010000000100",
			4272 => "1111111100001100000101",
			4273 => "0000001100001100000101",
			4274 => "0000110110100000001000",
			4275 => "0011101001001000000100",
			4276 => "0000100100001100000101",
			4277 => "0000001100001100000101",
			4278 => "0001010110110100000100",
			4279 => "0001000100001100000101",
			4280 => "0000001100001100000101",
			4281 => "0001101101011000000100",
			4282 => "0000000100001100000101",
			4283 => "0001001101000000000100",
			4284 => "0000000100001100000101",
			4285 => "0011111100010100000100",
			4286 => "0000001100001100000101",
			4287 => "0000001100001100000101",
			4288 => "1111111100001100000101",
			4289 => "0001111001110000001000",
			4290 => "0000101000100000000100",
			4291 => "1111111100001110100001",
			4292 => "0000000100001110100001",
			4293 => "0001111001110000001100",
			4294 => "0000100110010000001000",
			4295 => "0011010100011000000100",
			4296 => "0000000100001110100001",
			4297 => "0000001100001110100001",
			4298 => "0000000100001110100001",
			4299 => "0010000111000100010100",
			4300 => "0001000010111000000100",
			4301 => "1111111100001110100001",
			4302 => "0000010101011100001100",
			4303 => "0000011001111000000100",
			4304 => "0000000100001110100001",
			4305 => "0011001000111000000100",
			4306 => "0000000100001110100001",
			4307 => "0000000100001110100001",
			4308 => "0000000100001110100001",
			4309 => "0011110101110000011000",
			4310 => "0011101100101100001100",
			4311 => "0000101111100100001000",
			4312 => "0011001000111000000100",
			4313 => "0000000100001110100001",
			4314 => "0000000100001110100001",
			4315 => "0000000100001110100001",
			4316 => "0001000001100100000100",
			4317 => "0000000100001110100001",
			4318 => "0011001000111000000100",
			4319 => "0000000100001110100001",
			4320 => "0000000100001110100001",
			4321 => "0000101000100000000100",
			4322 => "0000000100001110100001",
			4323 => "0011011011110100000100",
			4324 => "1111111100001110100001",
			4325 => "0000111001011100000100",
			4326 => "0000000100001110100001",
			4327 => "0000000100001110100001",
			4328 => "0011010100011000000100",
			4329 => "1111111100010000111101",
			4330 => "0011001110001100011100",
			4331 => "0000000010111100000100",
			4332 => "1111111100010000111101",
			4333 => "0000000010111100001000",
			4334 => "0010001011010100000100",
			4335 => "0000011100010000111101",
			4336 => "0000000100010000111101",
			4337 => "0001000100001100000100",
			4338 => "1111111100010000111101",
			4339 => "0001010111001000000100",
			4340 => "0000010100010000111101",
			4341 => "0001001011001000000100",
			4342 => "0000000100010000111101",
			4343 => "0000001100010000111101",
			4344 => "0011000100001000011100",
			4345 => "0011011110101100010100",
			4346 => "0011011011110100001100",
			4347 => "0001111100101000001000",
			4348 => "0001111100101000000100",
			4349 => "0000000100010000111101",
			4350 => "0000000100010000111101",
			4351 => "1111111100010000111101",
			4352 => "0000011001011000000100",
			4353 => "0000000100010000111101",
			4354 => "1111111100010000111101",
			4355 => "0001001010110100000100",
			4356 => "0000000100010000111101",
			4357 => "0000001100010000111101",
			4358 => "0000100101000000000100",
			4359 => "1111111100010000111101",
			4360 => "0011001010111000000100",
			4361 => "0000001100010000111101",
			4362 => "0000100101000000001000",
			4363 => "0011001001110100000100",
			4364 => "0000000100010000111101",
			4365 => "0000000100010000111101",
			4366 => "1111111100010000111101",
			4367 => "0011010100011000000100",
			4368 => "1111111100010011100001",
			4369 => "0000100110010000011000",
			4370 => "0001011001001000010000",
			4371 => "0010000111000100001100",
			4372 => "0000000010111100000100",
			4373 => "0000000100010011100001",
			4374 => "0011000011011100000100",
			4375 => "0000001100010011100001",
			4376 => "0000000100010011100001",
			4377 => "0000000100010011100001",
			4378 => "0010100110011100000100",
			4379 => "0000000100010011100001",
			4380 => "0000000100010011100001",
			4381 => "0000011101101000011000",
			4382 => "0011100100000100010100",
			4383 => "0001011001110100001000",
			4384 => "0011100110000100000100",
			4385 => "0000000100010011100001",
			4386 => "0000000100010011100001",
			4387 => "0001101101011000000100",
			4388 => "0000000100010011100001",
			4389 => "0000000101110100000100",
			4390 => "0000000100010011100001",
			4391 => "0000000100010011100001",
			4392 => "1111111100010011100001",
			4393 => "0000011001011000010000",
			4394 => "0000101100001100001100",
			4395 => "0001101011001100000100",
			4396 => "0000000100010011100001",
			4397 => "0000011011101000000100",
			4398 => "0000000100010011100001",
			4399 => "0000000100010011100001",
			4400 => "0000000100010011100001",
			4401 => "0000100110001100000100",
			4402 => "0000000100010011100001",
			4403 => "0010100001010000001000",
			4404 => "0010011001111100000100",
			4405 => "0000000100010011100001",
			4406 => "0000000100010011100001",
			4407 => "0000000100010011100001",
			4408 => "0000101000001100101000",
			4409 => "0000010010001100000100",
			4410 => "1111111100010110110101",
			4411 => "0010100101000100011100",
			4412 => "0011110000110100011000",
			4413 => "0010101010110000010000",
			4414 => "0011110000110100001000",
			4415 => "0010100110011000000100",
			4416 => "1111111100010110110101",
			4417 => "0000000100010110110101",
			4418 => "0010101001000100000100",
			4419 => "0000000100010110110101",
			4420 => "0000011100010110110101",
			4421 => "0000111110110000000100",
			4422 => "1111111100010110110101",
			4423 => "0000110100010110110101",
			4424 => "1111111100010110110101",
			4425 => "0010111100101100000100",
			4426 => "1111111100010110110101",
			4427 => "0000001100010110110101",
			4428 => "0011000100001000110100",
			4429 => "0001100100111100101000",
			4430 => "0011010100010000010100",
			4431 => "0010011011101000001000",
			4432 => "0000101000001100000100",
			4433 => "0000000100010110110101",
			4434 => "1111111100010110110101",
			4435 => "0010101010110000000100",
			4436 => "1111111100010110110101",
			4437 => "0001101101011000000100",
			4438 => "0000000100010110110101",
			4439 => "0000001100010110110101",
			4440 => "0010011000010000010000",
			4441 => "0011100111110000001000",
			4442 => "0010011101011000000100",
			4443 => "0000010100010110110101",
			4444 => "0000000100010110110101",
			4445 => "0010001011010100000100",
			4446 => "0000010100010110110101",
			4447 => "0000100100010110110101",
			4448 => "1111111100010110110101",
			4449 => "0001011110101100001000",
			4450 => "0010001101010000000100",
			4451 => "1111111100010110110101",
			4452 => "1111110100010110110101",
			4453 => "0000001100010110110101",
			4454 => "0011101101101100001100",
			4455 => "0000100101000000000100",
			4456 => "1111111100010110110101",
			4457 => "0010000001110100000100",
			4458 => "0000011100010110110101",
			4459 => "0000000100010110110101",
			4460 => "1111111100010110110101",
			4461 => "0011010100011000000100",
			4462 => "1111111100011001101001",
			4463 => "0011000011011100011100",
			4464 => "0011100100001000001100",
			4465 => "0001001110111000000100",
			4466 => "0000000100011001101001",
			4467 => "0001101111000000000100",
			4468 => "0000001100011001101001",
			4469 => "0000000100011001101001",
			4470 => "0011000011011100001000",
			4471 => "0001001101000000000100",
			4472 => "1111111100011001101001",
			4473 => "0000000100011001101001",
			4474 => "0010010001000100000100",
			4475 => "0000000100011001101001",
			4476 => "0000001100011001101001",
			4477 => "0001101011001100001100",
			4478 => "0011001100110000001000",
			4479 => "0011101010111100000100",
			4480 => "0000000100011001101001",
			4481 => "0000000100011001101001",
			4482 => "1111111100011001101001",
			4483 => "0001101111000000011100",
			4484 => "0001001101110100001100",
			4485 => "0011011001010100000100",
			4486 => "0000000100011001101001",
			4487 => "0000010000111100000100",
			4488 => "0000000100011001101001",
			4489 => "0000000100011001101001",
			4490 => "0000011101011100001000",
			4491 => "0010011111001100000100",
			4492 => "0000000100011001101001",
			4493 => "0000001100011001101001",
			4494 => "0000101111100100000100",
			4495 => "0000000100011001101001",
			4496 => "0000000100011001101001",
			4497 => "0000101000011100001000",
			4498 => "0000110010110100000100",
			4499 => "0000000100011001101001",
			4500 => "1111111100011001101001",
			4501 => "0000111111101000001000",
			4502 => "0010100101000100000100",
			4503 => "0000001100011001101001",
			4504 => "0000000100011001101001",
			4505 => "1111111100011001101001",
			4506 => "0011010100011000000100",
			4507 => "1111111100011100010101",
			4508 => "0011001100110000101100",
			4509 => "0011001001110000011000",
			4510 => "0011100100001000010000",
			4511 => "0001000111011100000100",
			4512 => "0000000100011100010101",
			4513 => "0001101001100100001000",
			4514 => "0011011000011000000100",
			4515 => "0000001100011100010101",
			4516 => "0000000100011100010101",
			4517 => "0000000100011100010101",
			4518 => "0001001101000000000100",
			4519 => "1111111100011100010101",
			4520 => "0000000100011100010101",
			4521 => "0011110110010000010000",
			4522 => "0010001001101000000100",
			4523 => "0000000100011100010101",
			4524 => "0000011001111000000100",
			4525 => "0000000100011100010101",
			4526 => "0010100001010000000100",
			4527 => "0000001100011100010101",
			4528 => "0000001100011100010101",
			4529 => "0000000100011100010101",
			4530 => "0001101101011000001000",
			4531 => "0011001100110000000100",
			4532 => "0000000100011100010101",
			4533 => "1111111100011100010101",
			4534 => "0000010101011100011100",
			4535 => "0010101010110000001100",
			4536 => "0011010101110100000100",
			4537 => "0000000100011100010101",
			4538 => "0010100110011000000100",
			4539 => "0000000100011100010101",
			4540 => "0000001100011100010101",
			4541 => "0011110111011000001000",
			4542 => "0010100101000100000100",
			4543 => "0000000100011100010101",
			4544 => "0000001100011100010101",
			4545 => "0010011001100100000100",
			4546 => "1111111100011100010101",
			4547 => "0000000100011100010101",
			4548 => "1111111100011100010101",
			4549 => "0011010100011000000100",
			4550 => "1111111100011110100001",
			4551 => "0000100010011100001100",
			4552 => "0010110110000100001000",
			4553 => "0001001111100100000100",
			4554 => "0000000100011110100001",
			4555 => "0000001100011110100001",
			4556 => "0000000100011110100001",
			4557 => "0001000011010100000100",
			4558 => "1111111100011110100001",
			4559 => "0010100110011100011100",
			4560 => "0011001110001100001100",
			4561 => "0011001000111000000100",
			4562 => "0000000100011110100001",
			4563 => "0010100110011000000100",
			4564 => "0000000100011110100001",
			4565 => "0000001100011110100001",
			4566 => "0011110111011000001000",
			4567 => "0011111100010100000100",
			4568 => "0000000100011110100001",
			4569 => "0000000100011110100001",
			4570 => "0000010101011100000100",
			4571 => "0000000100011110100001",
			4572 => "0000000100011110100001",
			4573 => "0001100100111100010000",
			4574 => "0001101001100100001000",
			4575 => "0011001100110000000100",
			4576 => "0000000100011110100001",
			4577 => "0000000100011110100001",
			4578 => "0001000110110000000100",
			4579 => "0000000100011110100001",
			4580 => "0000000100011110100001",
			4581 => "0000011101011100000100",
			4582 => "1111111100011110100001",
			4583 => "0000000100011110100001",
			4584 => "0010110101101100000100",
			4585 => "1111111100100000101101",
			4586 => "0001000010111000000100",
			4587 => "1111111100100000101101",
			4588 => "0010000111000100011000",
			4589 => "0000010101011100010100",
			4590 => "0011000011011100000100",
			4591 => "0000001100100000101101",
			4592 => "0011001110001100001000",
			4593 => "0011010101110100000100",
			4594 => "0000000100100000101101",
			4595 => "0000000100100000101101",
			4596 => "0011010101110100000100",
			4597 => "0000000100100000101101",
			4598 => "0000001100100000101101",
			4599 => "0000000100100000101101",
			4600 => "0001101011001100010100",
			4601 => "0011001100110000001100",
			4602 => "0001000001100100000100",
			4603 => "0000000100100000101101",
			4604 => "0000010010001100000100",
			4605 => "0000000100100000101101",
			4606 => "0000000100100000101101",
			4607 => "0011100100011000000100",
			4608 => "1111111100100000101101",
			4609 => "0000000100100000101101",
			4610 => "0001101111000000001100",
			4611 => "0001000010010000000100",
			4612 => "0000000100100000101101",
			4613 => "0000011111001100000100",
			4614 => "0000001100100000101101",
			4615 => "0000000100100000101101",
			4616 => "0011111100010100000100",
			4617 => "0000000100100000101101",
			4618 => "1111111100100000101101",
			4619 => "0000011001111000000100",
			4620 => "1111111100100011011011",
			4621 => "0010100110011100100100",
			4622 => "0000001111000100000100",
			4623 => "1111111100100011011011",
			4624 => "0011001000111000000100",
			4625 => "0000000100100011011011",
			4626 => "0010100001010000001100",
			4627 => "0000010000111100001000",
			4628 => "0010101001000100000100",
			4629 => "0000000100100011011011",
			4630 => "0000001100100011011011",
			4631 => "0000000100100011011011",
			4632 => "0001001100111100001000",
			4633 => "0011000000001100000100",
			4634 => "0000000100100011011011",
			4635 => "0000000100100011011011",
			4636 => "0011100100010000000100",
			4637 => "0000000100100011011011",
			4638 => "0000001100100011011011",
			4639 => "0000001100101100101000",
			4640 => "0011001110001100011100",
			4641 => "0011001100110000010000",
			4642 => "0001011001110100001000",
			4643 => "0001101011001100000100",
			4644 => "0000000100100011011011",
			4645 => "0000000100100011011011",
			4646 => "0001101000010000000100",
			4647 => "0000000100100011011011",
			4648 => "0000000100100011011011",
			4649 => "0000101111100100000100",
			4650 => "0000000100100011011011",
			4651 => "0000100011000000000100",
			4652 => "1111111100100011011011",
			4653 => "0000000100100011011011",
			4654 => "0011000100001000001000",
			4655 => "0010010111101000000100",
			4656 => "0000000100100011011011",
			4657 => "0000000100100011011011",
			4658 => "0000000100100011011011",
			4659 => "0000101100001100000100",
			4660 => "0000001100100011011011",
			4661 => "0000000100100011011011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1522, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(3074, initial_addr_3'length));
	end generate gen_rom_13;

	gen_rom_14: if SELECT_ROM = 14 generate
		bank <= (
			0 => "0001111101111001011000",
			1 => "0001001011100101010100",
			2 => "0001100001000100010100",
			3 => "0000110000111000001000",
			4 => "0011111000000000000100",
			5 => "0000001000000011010101",
			6 => "0000000000000011010101",
			7 => "0000110111111000001000",
			8 => "0011101010101100000100",
			9 => "1111111000000011010101",
			10 => "0000000000000011010101",
			11 => "1111111000000011010101",
			12 => "0001111100001000100000",
			13 => "0000111101100000010000",
			14 => "0001110111111000001000",
			15 => "0000100010000000000100",
			16 => "0000001000000011010101",
			17 => "1111111000000011010101",
			18 => "0010100111110100000100",
			19 => "0000001000000011010101",
			20 => "0000000000000011010101",
			21 => "0000101001010000001000",
			22 => "0001000010111000000100",
			23 => "0000001000000011010101",
			24 => "0000010000000011010101",
			25 => "0010100110011000000100",
			26 => "0000000000000011010101",
			27 => "0000001000000011010101",
			28 => "0011101101111000010000",
			29 => "0000101100010100001000",
			30 => "0001100001111000000100",
			31 => "1111111000000011010101",
			32 => "0000000000000011010101",
			33 => "0001111000111000000100",
			34 => "0000000000000011010101",
			35 => "0000001000000011010101",
			36 => "0001111000111000001000",
			37 => "0011100100000100000100",
			38 => "0000001000000011010101",
			39 => "1111111000000011010101",
			40 => "0001101111000000000100",
			41 => "0000000000000011010101",
			42 => "1111111000000011010101",
			43 => "1111111000000011010101",
			44 => "0010100111110100010000",
			45 => "0011111000101000001100",
			46 => "0001111100101000001000",
			47 => "0010000000001000000100",
			48 => "1111111000000011010101",
			49 => "0000001000000011010101",
			50 => "1111111000000011010101",
			51 => "0000010000000011010101",
			52 => "1111111000000011010101",
			53 => "0000001100001010001000",
			54 => "0001011000111100011100",
			55 => "0000000111111000001100",
			56 => "0010011100110100001000",
			57 => "0001011100001000000100",
			58 => "0000000000001001011001",
			59 => "0000000000001001011001",
			60 => "0000001000001001011001",
			61 => "0001001111100000000100",
			62 => "1111111000001001011001",
			63 => "0010111010000000000100",
			64 => "0000000000001001011001",
			65 => "0010100001010000000100",
			66 => "0000000000001001011001",
			67 => "0000001000001001011001",
			68 => "0000011110100000110000",
			69 => "0010011001111000100000",
			70 => "0000101001010000010000",
			71 => "0001101101111100001000",
			72 => "0011111011011100000100",
			73 => "0000000000001001011001",
			74 => "0000010000001001011001",
			75 => "0000010110000000000100",
			76 => "0000000000001001011001",
			77 => "0000001000001001011001",
			78 => "0000100101110000001000",
			79 => "0000000000111000000100",
			80 => "0000001000001001011001",
			81 => "1111111000001001011001",
			82 => "0000010110000000000100",
			83 => "0000000000001001011001",
			84 => "0000000000001001011001",
			85 => "0001010011011100001000",
			86 => "0011101110111100000100",
			87 => "1111111000001001011001",
			88 => "0000000000001001011001",
			89 => "0010101010110000000100",
			90 => "1111111000001001011001",
			91 => "0000000000001001011001",
			92 => "0011011100101100011100",
			93 => "0000110101101100001100",
			94 => "0010111100001000001000",
			95 => "0010110000101000000100",
			96 => "0000000000001001011001",
			97 => "0000000000001001011001",
			98 => "1111111000001001011001",
			99 => "0000101100010100001000",
			100 => "0000000000111000000100",
			101 => "0000000000001001011001",
			102 => "0000001000001001011001",
			103 => "0010010110101000000100",
			104 => "0000000000001001011001",
			105 => "1111111000001001011001",
			106 => "0000011100110100010000",
			107 => "0010110100000000001000",
			108 => "0011011101111000000100",
			109 => "0000000000001001011001",
			110 => "1111111000001001011001",
			111 => "0000011110100000000100",
			112 => "0000001000001001011001",
			113 => "0000000000001001011001",
			114 => "0010010111100100001000",
			115 => "0000111101111000000100",
			116 => "0000000000001001011001",
			117 => "0000001000001001011001",
			118 => "0000011100110100000100",
			119 => "0000000000001001011001",
			120 => "0000000000001001011001",
			121 => "0000100010000000100100",
			122 => "0011100000101000100000",
			123 => "0000110100000000010100",
			124 => "0011110110110100010000",
			125 => "0010100110011100001000",
			126 => "0011100011111100000100",
			127 => "1111111000001001011001",
			128 => "0000000000001001011001",
			129 => "0000001000111100000100",
			130 => "0000000000001001011001",
			131 => "0000000000001001011001",
			132 => "0000001000001001011001",
			133 => "0010100001010100000100",
			134 => "1111111000001001011001",
			135 => "0011111011011100000100",
			136 => "0000000000001001011001",
			137 => "0000000000001001011001",
			138 => "0000001000001001011001",
			139 => "0000010010001100010000",
			140 => "0010001000110000000100",
			141 => "1111111000001001011001",
			142 => "0000011110100000001000",
			143 => "0011110101110100000100",
			144 => "0000000000001001011001",
			145 => "0000001000001001011001",
			146 => "1111111000001001011001",
			147 => "0010111100110000000100",
			148 => "0000001000001001011001",
			149 => "1111111000001001011001",
			150 => "0010011001111001010000",
			151 => "0011000100010100101100",
			152 => "0011000100010100101000",
			153 => "0000100010000000100000",
			154 => "0001000001101100010000",
			155 => "0011101111000100001000",
			156 => "0010110100010100000100",
			157 => "0000000000001110111101",
			158 => "1111111000001110111101",
			159 => "0011000000110000000100",
			160 => "0000000000001110111101",
			161 => "0000000000001110111101",
			162 => "0010100001010100001000",
			163 => "0011011000111000000100",
			164 => "0000010000001110111101",
			165 => "0000000000001110111101",
			166 => "0010110111111000000100",
			167 => "0000000000001110111101",
			168 => "0000001000001110111101",
			169 => "0001000100001100000100",
			170 => "0000000000001110111101",
			171 => "1111111000001110111101",
			172 => "1111111000001110111101",
			173 => "0000010110000000001100",
			174 => "0011100000111000001000",
			175 => "0000010000011000000100",
			176 => "0000000000001110111101",
			177 => "1111111000001110111101",
			178 => "0000000000001110111101",
			179 => "0011000000101000010100",
			180 => "0011101110111100010000",
			181 => "0011011100110000001000",
			182 => "0010010010001100000100",
			183 => "0000001000001110111101",
			184 => "0000000000001110111101",
			185 => "0010111011000100000100",
			186 => "0000000000001110111101",
			187 => "0000000000001110111101",
			188 => "0000001000001110111101",
			189 => "1111111000001110111101",
			190 => "0000011110100000110000",
			191 => "0011000000110000000100",
			192 => "0000001000001110111101",
			193 => "0000101001011100010100",
			194 => "0001001011100000010000",
			195 => "0011100100010100001000",
			196 => "0001110111111000000100",
			197 => "0000001000001110111101",
			198 => "0000000000001110111101",
			199 => "0000011110100000000100",
			200 => "0000000000001110111101",
			201 => "0000001000001110111101",
			202 => "0000001000001110111101",
			203 => "0010011001111000001100",
			204 => "0010011001111000001000",
			205 => "0011111011110100000100",
			206 => "1111111000001110111101",
			207 => "0000000000001110111101",
			208 => "0000000000001110111101",
			209 => "0001100100110100000100",
			210 => "1111111000001110111101",
			211 => "0000001011000100000100",
			212 => "0000000000001110111101",
			213 => "1111111000001110111101",
			214 => "0001110111111000000100",
			215 => "0000001000001110111101",
			216 => "0011001010000000010100",
			217 => "0011010110000100001100",
			218 => "0000011110100000001000",
			219 => "0011100100010100000100",
			220 => "1111111000001110111101",
			221 => "0000000000001110111101",
			222 => "0000001000001110111101",
			223 => "0001001110111000000100",
			224 => "1111111000001110111101",
			225 => "0000000000001110111101",
			226 => "0011001110111100001100",
			227 => "0000101111010000000100",
			228 => "0000000000001110111101",
			229 => "0001110100010100000100",
			230 => "0000001000001110111101",
			231 => "0000000000001110111101",
			232 => "0011011100110000001000",
			233 => "0001001110111000000100",
			234 => "1111111000001110111101",
			235 => "0000000000001110111101",
			236 => "0011001000111000000100",
			237 => "0000000000001110111101",
			238 => "0000000000001110111101",
			239 => "0011000100000010010100",
			240 => "0001111001110001100100",
			241 => "0001111000111000111100",
			242 => "0011000100000000100000",
			243 => "0000100100101000010000",
			244 => "0000100100101000001000",
			245 => "0000010010001100000100",
			246 => "0000000000010101110001",
			247 => "0000000000010101110001",
			248 => "0010101010110000000100",
			249 => "0000001000010101110001",
			250 => "0000000000010101110001",
			251 => "0010101010110000001000",
			252 => "0011101101100000000100",
			253 => "0000000000010101110001",
			254 => "0000000000010101110001",
			255 => "0011000100010100000100",
			256 => "0000000000010101110001",
			257 => "0000000000010101110001",
			258 => "0010101100011100010000",
			259 => "0010110100000000001000",
			260 => "0000101001010000000100",
			261 => "0000000000010101110001",
			262 => "0000001000010101110001",
			263 => "0011110110100000000100",
			264 => "1111111000010101110001",
			265 => "0000000000010101110001",
			266 => "0010101100011100000100",
			267 => "0000001000010101110001",
			268 => "0001101101011000000100",
			269 => "0000000000010101110001",
			270 => "0000001000010101110001",
			271 => "0000000111111000100000",
			272 => "0010000110001000010000",
			273 => "0011111100100100001000",
			274 => "0011000000101000000100",
			275 => "0000000000010101110001",
			276 => "0000001000010101110001",
			277 => "0010100001010000000100",
			278 => "1111111000010101110001",
			279 => "0000001000010101110001",
			280 => "0010101010110000001000",
			281 => "0011011010111000000100",
			282 => "0000001000010101110001",
			283 => "0000001000010101110001",
			284 => "0000110001101000000100",
			285 => "0000000000010101110001",
			286 => "0000001000010101110001",
			287 => "0011010111001000000100",
			288 => "1111111000010101110001",
			289 => "0000000000010101110001",
			290 => "0000100010000100011100",
			291 => "0000010110101000010000",
			292 => "0000100101110000000100",
			293 => "0000000000010101110001",
			294 => "0001111101100000000100",
			295 => "1111111000010101110001",
			296 => "0011101110110000000100",
			297 => "0000000000010101110001",
			298 => "1111111000010101110001",
			299 => "0011011001001000000100",
			300 => "0000001000010101110001",
			301 => "0001111101100000000100",
			302 => "1111111000010101110001",
			303 => "0000000000010101110001",
			304 => "0000000000111000001000",
			305 => "0010111110001100000100",
			306 => "1111111000010101110001",
			307 => "0000000000010101110001",
			308 => "0001101011001100000100",
			309 => "0000001000010101110001",
			310 => "0001111101100000000100",
			311 => "1111111000010101110001",
			312 => "0000000000010101110001",
			313 => "0011000100000000011000",
			314 => "0000100011001000001000",
			315 => "0000101111010000000100",
			316 => "0000000000010101110001",
			317 => "0000001000010101110001",
			318 => "0000101100010100000100",
			319 => "0000000000010101110001",
			320 => "0011011010111100000100",
			321 => "0000000000010101110001",
			322 => "0000011001111000000100",
			323 => "0000001000010101110001",
			324 => "0000000000010101110001",
			325 => "0000000100010100101000",
			326 => "0010000010101000100000",
			327 => "0011001000111100010000",
			328 => "0011001000111100001000",
			329 => "0011101010111000000100",
			330 => "0000000000010101110001",
			331 => "0000001000010101110001",
			332 => "0001101010011000000100",
			333 => "0000000000010101110001",
			334 => "1111111000010101110001",
			335 => "0000010010001100001000",
			336 => "0001101010011000000100",
			337 => "0000000000010101110001",
			338 => "1111111000010101110001",
			339 => "0001101010011000000100",
			340 => "0000000000010101110001",
			341 => "0000000000010101110001",
			342 => "0000100111010100000100",
			343 => "0000010000010101110001",
			344 => "0000000000010101110001",
			345 => "0010111001110000000100",
			346 => "0000000000010101110001",
			347 => "1111111000010101110001",
			348 => "0001110101101101111000",
			349 => "0000010000011000001000",
			350 => "0001100100110100000100",
			351 => "1111111000011011010101",
			352 => "0000000000011011010101",
			353 => "0001001110111000111100",
			354 => "0001101101111100100000",
			355 => "0000100101110000010000",
			356 => "0000000000110000001000",
			357 => "0001101101111100000100",
			358 => "0000000000011011010101",
			359 => "0000001000011011010101",
			360 => "0001000101010100000100",
			361 => "1111111000011011010101",
			362 => "0000000000011011010101",
			363 => "0000001111000100001000",
			364 => "0001001011110000000100",
			365 => "0000000000011011010101",
			366 => "1111111000011011010101",
			367 => "0000111101111000000100",
			368 => "0000000000011011010101",
			369 => "0000001000011011010101",
			370 => "0011000100000000001100",
			371 => "0000010110101000001000",
			372 => "0001000011001100000100",
			373 => "0000001000011011010101",
			374 => "0000001000011011010101",
			375 => "1111111000011011010101",
			376 => "0011000100000000001000",
			377 => "0001000011001100000100",
			378 => "1111111000011011010101",
			379 => "1111111000011011010101",
			380 => "0001101001100100000100",
			381 => "0000000000011011010101",
			382 => "1111111000011011010101",
			383 => "0011000100010100010100",
			384 => "0010100110011000000100",
			385 => "1111111000011011010101",
			386 => "0010011001111000001000",
			387 => "0000111100001000000100",
			388 => "0000000000011011010101",
			389 => "0000010000011011010101",
			390 => "0000111001110000000100",
			391 => "0000000000011011010101",
			392 => "0000001000011011010101",
			393 => "0001101100011000010000",
			394 => "0000101001011100001000",
			395 => "0001110100010100000100",
			396 => "1111111000011011010101",
			397 => "0000000000011011010101",
			398 => "0010010111100100000100",
			399 => "0000000000011011010101",
			400 => "1111111000011011010101",
			401 => "0001000010100100001000",
			402 => "0010010110101000000100",
			403 => "0000001000011011010101",
			404 => "0000000000011011010101",
			405 => "0011000100010100000100",
			406 => "0000000000011011010101",
			407 => "0000000000011011010101",
			408 => "0011000110000100100100",
			409 => "0011010111010000010000",
			410 => "0011101001001000000100",
			411 => "1111111000011011010101",
			412 => "0011100100000100001000",
			413 => "0000001101010000000100",
			414 => "1111111000011011010101",
			415 => "0000001000011011010101",
			416 => "1111111000011011010101",
			417 => "0001001001001100010000",
			418 => "0000001001101000000100",
			419 => "1111111000011011010101",
			420 => "0001101111000000000100",
			421 => "0000010000011011010101",
			422 => "0010101100011100000100",
			423 => "1111111000011011010101",
			424 => "0000000000011011010101",
			425 => "1111111000011011010101",
			426 => "0011001010111100010100",
			427 => "0001110110100100010000",
			428 => "0001111101111000001100",
			429 => "0001111110001100000100",
			430 => "1111111000011011010101",
			431 => "0011000110000100000100",
			432 => "0000000000011011010101",
			433 => "0000000000011011010101",
			434 => "1111111000011011010101",
			435 => "0000010000011011010101",
			436 => "1111111000011011010101",
			437 => "0011101000000010010000",
			438 => "0010011111001101011100",
			439 => "0000011001111000110000",
			440 => "0010011011101000100000",
			441 => "0001101100011000010000",
			442 => "0000101100010100001000",
			443 => "0011000000101000000100",
			444 => "0000000000100010101001",
			445 => "0000000000100010101001",
			446 => "0010011101101000000100",
			447 => "0000000000100010101001",
			448 => "1111111000100010101001",
			449 => "0011000100000000001000",
			450 => "0000110101101100000100",
			451 => "0000000000100010101001",
			452 => "0000000000100010101001",
			453 => "0000110100011000000100",
			454 => "0000000000100010101001",
			455 => "0000000000100010101001",
			456 => "0001000011010100001100",
			457 => "0001010111001000001000",
			458 => "0000001110111100000100",
			459 => "0000000000100010101001",
			460 => "1111111000100010101001",
			461 => "1111111000100010101001",
			462 => "0000001000100010101001",
			463 => "0001000011110000010100",
			464 => "0001100001111000001000",
			465 => "0010011011101000000100",
			466 => "0000000000100010101001",
			467 => "0000010000100010101001",
			468 => "0000111110110000001000",
			469 => "0001111000111000000100",
			470 => "0000001000100010101001",
			471 => "0000000000100010101001",
			472 => "0000001000100010101001",
			473 => "0000111000000000001100",
			474 => "0010011011101000000100",
			475 => "0000001000100010101001",
			476 => "0000000000110000000100",
			477 => "0000000000100010101001",
			478 => "1111111000100010101001",
			479 => "0001000100001100001000",
			480 => "0000011001111000000100",
			481 => "0000001000100010101001",
			482 => "0000000000100010101001",
			483 => "0000000000100010101001",
			484 => "0000000000110000011100",
			485 => "0000011001111000000100",
			486 => "1111111000100010101001",
			487 => "0001001000001000001100",
			488 => "0000010110101000001000",
			489 => "0000111001001000000100",
			490 => "0000000000100010101001",
			491 => "0000000000100010101001",
			492 => "1111111000100010101001",
			493 => "0001000010111000000100",
			494 => "0000001000100010101001",
			495 => "0000100110010000000100",
			496 => "1111111000100010101001",
			497 => "0000001000100010101001",
			498 => "0010011001011000010000",
			499 => "0001101001100100000100",
			500 => "1111111000100010101001",
			501 => "0001010100011000000100",
			502 => "1111111000100010101001",
			503 => "0000011001111000000100",
			504 => "0000001000100010101001",
			505 => "0000000000100010101001",
			506 => "0010110000001100000100",
			507 => "0000001000100010101001",
			508 => "0000000000100010101001",
			509 => "0001101001100101000100",
			510 => "0011001000111100100100",
			511 => "0011000000101000001000",
			512 => "0001000011110000000100",
			513 => "0000001000100010101001",
			514 => "1111111000100010101001",
			515 => "0010000110001000010000",
			516 => "0010001001101000001000",
			517 => "0000100111111100000100",
			518 => "0000000000100010101001",
			519 => "0000001000100010101001",
			520 => "0010001011010100000100",
			521 => "1111111000100010101001",
			522 => "0000000000100010101001",
			523 => "0011000100000000001000",
			524 => "0011001100001000000100",
			525 => "0000001000100010101001",
			526 => "0000001000100010101001",
			527 => "0000000000100010101001",
			528 => "0011001000111100000100",
			529 => "1111111000100010101001",
			530 => "0000111111011100001100",
			531 => "0001110101101100000100",
			532 => "1111111000100010101001",
			533 => "0001010001101000000100",
			534 => "0000001000100010101001",
			535 => "0000000000100010101001",
			536 => "0000110100000100001000",
			537 => "0011000011011100000100",
			538 => "0000001000100010101001",
			539 => "0000000000100010101001",
			540 => "0011010001101000000100",
			541 => "0000000000100010101001",
			542 => "0000000000100010101001",
			543 => "0011011000000000001000",
			544 => "0011101000011000000100",
			545 => "0000000000100010101001",
			546 => "0000001000100010101001",
			547 => "0001100100111100000100",
			548 => "1111111000100010101001",
			549 => "0000101111010100001000",
			550 => "0001010110100100000100",
			551 => "0000000000100010101001",
			552 => "0000001000100010101001",
			553 => "1111111000100010101001",
			554 => "0011000110000110001000",
			555 => "0000010000011000001100",
			556 => "0001100100110100000100",
			557 => "1111111000100111100101",
			558 => "0001110111111000000100",
			559 => "0000001000100111100101",
			560 => "1111111000100111100101",
			561 => "0010011001111001000000",
			562 => "0000110100000000100000",
			563 => "0010011001111000010000",
			564 => "0000110100010100001000",
			565 => "0011000000110000000100",
			566 => "0000001000100111100101",
			567 => "0000000000100111100101",
			568 => "0011110110100100000100",
			569 => "0000010000100111100101",
			570 => "0000000000100111100101",
			571 => "0000011110100000001000",
			572 => "0011000111111000000100",
			573 => "0000000000100111100101",
			574 => "1111111000100111100101",
			575 => "0011111010001100000100",
			576 => "0000001000100111100101",
			577 => "1111111000100111100101",
			578 => "0011110101100100010000",
			579 => "0011100000110000001000",
			580 => "0010100001010000000100",
			581 => "0000000000100111100101",
			582 => "0000001000100111100101",
			583 => "0000001111000100000100",
			584 => "0000000000100111100101",
			585 => "0000010000100111100101",
			586 => "0010001001101000001000",
			587 => "0011100100010100000100",
			588 => "1111111000100111100101",
			589 => "0000000000100111100101",
			590 => "0000111001110000000100",
			591 => "0000000000100111100101",
			592 => "0000001000100111100101",
			593 => "0011101000111100011100",
			594 => "0000111110001100010000",
			595 => "0000111100101100001000",
			596 => "0000111100101100000100",
			597 => "0000000000100111100101",
			598 => "1111111000100111100101",
			599 => "0000101001011100000100",
			600 => "0000001000100111100101",
			601 => "0000000000100111100101",
			602 => "0010001010101100001000",
			603 => "0011110101100100000100",
			604 => "0000000000100111100101",
			605 => "1111111000100111100101",
			606 => "0000010000100111100101",
			607 => "0010011101101000010000",
			608 => "0000100010000000001000",
			609 => "0001111100001000000100",
			610 => "0000000000100111100101",
			611 => "0000001000100111100101",
			612 => "0001101100011000000100",
			613 => "0000000000100111100101",
			614 => "0000000000100111100101",
			615 => "0011101101111000001000",
			616 => "0011011101111000000100",
			617 => "0000001000100111100101",
			618 => "0000000000100111100101",
			619 => "0010011111001100000100",
			620 => "0000000000100111100101",
			621 => "0000000000100111100101",
			622 => "0011001010111100010100",
			623 => "0011011001010000010000",
			624 => "0001111101111000001100",
			625 => "0001111110001100000100",
			626 => "1111111000100111100101",
			627 => "0011000110000100000100",
			628 => "0000000000100111100101",
			629 => "0000000000100111100101",
			630 => "1111111000100111100101",
			631 => "0000010000100111100101",
			632 => "1111111000100111100101",
			633 => "0001110101101101101100",
			634 => "0000011100100000000100",
			635 => "1111111000101101000001",
			636 => "0001001110111000111000",
			637 => "0001111001110000100000",
			638 => "0001101101111100010000",
			639 => "0000100111111100001000",
			640 => "0011101000111100000100",
			641 => "0000000000101101000001",
			642 => "0000001000101101000001",
			643 => "0000000010111100000100",
			644 => "1111111000101101000001",
			645 => "0000000000101101000001",
			646 => "0001111100001000001000",
			647 => "0011111011110100000100",
			648 => "0000001000101101000001",
			649 => "0000001000101101000001",
			650 => "0011100110000100000100",
			651 => "0000000000101101000001",
			652 => "0000001000101101000001",
			653 => "0010000111000100001100",
			654 => "0001101001100100001000",
			655 => "0011111010010100000100",
			656 => "1111111000101101000001",
			657 => "0000001000101101000001",
			658 => "1111111000101101000001",
			659 => "0001001001001100001000",
			660 => "0000100110111100000100",
			661 => "1111111000101101000001",
			662 => "0000000000101101000001",
			663 => "0000000000101101000001",
			664 => "0010010110101000010100",
			665 => "0001100111101000000100",
			666 => "1111111000101101000001",
			667 => "0011101011000100001000",
			668 => "0001110111111000000100",
			669 => "0000001000101101000001",
			670 => "0000000000101101000001",
			671 => "0000101100010100000100",
			672 => "0000001000101101000001",
			673 => "0000001000101101000001",
			674 => "0000110101101100001100",
			675 => "0011010110000100000100",
			676 => "0000001000101101000001",
			677 => "0000101111010000000100",
			678 => "0000000000101101000001",
			679 => "1111111000101101000001",
			680 => "0001101100011000001000",
			681 => "0011101001110000000100",
			682 => "0000000000101101000001",
			683 => "1111111000101101000001",
			684 => "0001001111100000000100",
			685 => "0000000000101101000001",
			686 => "0000000000101101000001",
			687 => "0001111100101000100100",
			688 => "0011101001001000000100",
			689 => "1111111000101101000001",
			690 => "0000100111010100011100",
			691 => "0011010111010000001100",
			692 => "0011100100000100001000",
			693 => "0000001101010000000100",
			694 => "1111111000101101000001",
			695 => "0000001000101101000001",
			696 => "1111111000101101000001",
			697 => "0001100100110100001000",
			698 => "0010111010111000000100",
			699 => "1111111000101101000001",
			700 => "0000000000101101000001",
			701 => "0010111101010100000100",
			702 => "0000010000101101000001",
			703 => "0000000000101101000001",
			704 => "1111111000101101000001",
			705 => "0010000110011100011100",
			706 => "0001001011110000010000",
			707 => "0001110001111100001100",
			708 => "0001110001111100001000",
			709 => "0001111100101000000100",
			710 => "0000000000101101000001",
			711 => "0000000000101101000001",
			712 => "0000000000101101000001",
			713 => "1111111000101101000001",
			714 => "0000000111000100000100",
			715 => "0000010000101101000001",
			716 => "0001001000110100000100",
			717 => "1111111000101101000001",
			718 => "0000001000101101000001",
			719 => "1111111000101101000001",
			720 => "0010011001111001101000",
			721 => "0011000100010100111000",
			722 => "0011000100010100110100",
			723 => "0001000001101100011100",
			724 => "0011101111000100001100",
			725 => "0010110100010100001000",
			726 => "0000100010110100000100",
			727 => "0000000000110011011101",
			728 => "0000000000110011011101",
			729 => "1111111000110011011101",
			730 => "0011110000011100001000",
			731 => "0010000111000100000100",
			732 => "0000000000110011011101",
			733 => "0000001000110011011101",
			734 => "0011000111111000000100",
			735 => "0000000000110011011101",
			736 => "0000001000110011011101",
			737 => "0010100001010100001100",
			738 => "0000101101000100000100",
			739 => "0000011000110011011101",
			740 => "0001001100111100000100",
			741 => "0000001000110011011101",
			742 => "0000000000110011011101",
			743 => "0010100001110000000100",
			744 => "1111111000110011011101",
			745 => "0001000011111000000100",
			746 => "0000000000110011011101",
			747 => "0000000000110011011101",
			748 => "1111111000110011011101",
			749 => "0000010110000000001000",
			750 => "0011100000111000000100",
			751 => "1111111000110011011101",
			752 => "0000000000110011011101",
			753 => "0000100001000000010100",
			754 => "0000101110101000001100",
			755 => "0001110100010100001000",
			756 => "0001100001111000000100",
			757 => "0000001000110011011101",
			758 => "1111111000110011011101",
			759 => "0000001000110011011101",
			760 => "0001001110111000000100",
			761 => "1111111000110011011101",
			762 => "0000000000110011011101",
			763 => "0011000100010100001100",
			764 => "0011011101100000000100",
			765 => "0000010000110011011101",
			766 => "0011100000111000000100",
			767 => "0000000000110011011101",
			768 => "0000001000110011011101",
			769 => "0010101100011100000100",
			770 => "0000001000110011011101",
			771 => "0000000000110011011101",
			772 => "0000011110100000101000",
			773 => "0011000000110000000100",
			774 => "0000001000110011011101",
			775 => "0000101001011100010100",
			776 => "0001001011100000010000",
			777 => "0011100100010100001000",
			778 => "0010110100010100000100",
			779 => "0000000000110011011101",
			780 => "0000000000110011011101",
			781 => "0001100001111000000100",
			782 => "0000001000110011011101",
			783 => "0000000000110011011101",
			784 => "0000001000110011011101",
			785 => "0010011001111000001100",
			786 => "0010100001010000000100",
			787 => "1111111000110011011101",
			788 => "0000000100010100000100",
			789 => "0000000000110011011101",
			790 => "1111111000110011011101",
			791 => "1111111000110011011101",
			792 => "0001110111111000000100",
			793 => "0000001000110011011101",
			794 => "0011001000111000100000",
			795 => "0010101001000100010000",
			796 => "0010101001000100001000",
			797 => "0011101000111100000100",
			798 => "0000000000110011011101",
			799 => "0000000000110011011101",
			800 => "0001001000110100000100",
			801 => "1111111000110011011101",
			802 => "0000000000110011011101",
			803 => "0010001011010100001000",
			804 => "0011111110101100000100",
			805 => "0000001000110011011101",
			806 => "0000000000110011011101",
			807 => "0010100110011000000100",
			808 => "0000000000110011011101",
			809 => "0000000000110011011101",
			810 => "0001001110111000010000",
			811 => "0001000011110000001000",
			812 => "0010001011010100000100",
			813 => "0000000000110011011101",
			814 => "1111111000110011011101",
			815 => "0000001110111100000100",
			816 => "0000000000110011011101",
			817 => "1111111000110011011101",
			818 => "0010000001110100000100",
			819 => "1111111000110011011101",
			820 => "0000000100010100000100",
			821 => "0000000000110011011101",
			822 => "1111111000110011011101",
			823 => "0000100010110101100100",
			824 => "0000100001001000101000",
			825 => "0000001000110000011000",
			826 => "0000111101100000001100",
			827 => "0000010110000000000100",
			828 => "0000000000111011011001",
			829 => "0011100000111000000100",
			830 => "0000000000111011011001",
			831 => "0000001000111011011001",
			832 => "0011111010011100000100",
			833 => "1111111000111011011001",
			834 => "0001001110010000000100",
			835 => "0000000000111011011001",
			836 => "0000000000111011011001",
			837 => "0011001010000000001100",
			838 => "0001110111111000001000",
			839 => "0001111110111100000100",
			840 => "0000000000111011011001",
			841 => "0000001000111011011001",
			842 => "1111111000111011011001",
			843 => "1111111000111011011001",
			844 => "0010101000010100011000",
			845 => "0001001110100100010000",
			846 => "0000111000111100000100",
			847 => "1111111000111011011001",
			848 => "0000001000110000001000",
			849 => "0000101110101100000100",
			850 => "0000000000111011011001",
			851 => "0000001000111011011001",
			852 => "0000001000111011011001",
			853 => "0000011110100000000100",
			854 => "0000000000111011011001",
			855 => "0000010000111011011001",
			856 => "0010101001000100001000",
			857 => "0001000010110000000100",
			858 => "1111111000111011011001",
			859 => "0000000000111011011001",
			860 => "0001100001111000001100",
			861 => "0011001010000000001000",
			862 => "0011001010000000000100",
			863 => "0000000000111011011001",
			864 => "0000001000111011011001",
			865 => "1111111000111011011001",
			866 => "0011001010000000001000",
			867 => "0000010000011000000100",
			868 => "0000000000111011011001",
			869 => "1111111000111011011001",
			870 => "0001110111111000000100",
			871 => "0000010000111011011001",
			872 => "0000001000111011011001",
			873 => "0011101111000101011000",
			874 => "0011110110100100100100",
			875 => "0000110111111000011000",
			876 => "0000010110000000010000",
			877 => "0000110011111100001000",
			878 => "0011010100000000000100",
			879 => "0000000000111011011001",
			880 => "1111111000111011011001",
			881 => "0010100110011100000100",
			882 => "0000000000111011011001",
			883 => "0000001000111011011001",
			884 => "0001001001001100000100",
			885 => "0000000000111011011001",
			886 => "1111111000111011011001",
			887 => "0000110111111000000100",
			888 => "0000001000111011011001",
			889 => "0001101100011000000100",
			890 => "0000000000111011011001",
			891 => "0000000000111011011001",
			892 => "0011101000110000100000",
			893 => "0011111000011000010000",
			894 => "0001100001111000001000",
			895 => "0010101010110000000100",
			896 => "0000000000111011011001",
			897 => "0000001000111011011001",
			898 => "0011100111000100000100",
			899 => "0000000000111011011001",
			900 => "1111111000111011011001",
			901 => "0000001011000100001000",
			902 => "0000001110111100000100",
			903 => "0000000000111011011001",
			904 => "0000001000111011011001",
			905 => "0001111011000100000100",
			906 => "0000000000111011011001",
			907 => "0000000000111011011001",
			908 => "0000011110100000001100",
			909 => "0010011100110100001000",
			910 => "0011111111011100000100",
			911 => "0000001000111011011001",
			912 => "1111111000111011011001",
			913 => "1111111000111011011001",
			914 => "0001001111100000000100",
			915 => "0000000000111011011001",
			916 => "0000000000111011011001",
			917 => "0011110110100100000100",
			918 => "0000001000111011011001",
			919 => "0010101001000100100000",
			920 => "0010101000010100010000",
			921 => "0001101100011000001000",
			922 => "0000000010111100000100",
			923 => "0000000000111011011001",
			924 => "0000000000111011011001",
			925 => "0011001000111000000100",
			926 => "0000001000111011011001",
			927 => "0000000000111011011001",
			928 => "0001101101111100001000",
			929 => "0010001001101000000100",
			930 => "0000001000111011011001",
			931 => "0000000000111011011001",
			932 => "0011010100001000000100",
			933 => "1111111000111011011001",
			934 => "0000000000111011011001",
			935 => "0011000100010100010000",
			936 => "0000011100110100001000",
			937 => "0001111011000100000100",
			938 => "0000000000111011011001",
			939 => "0000000000111011011001",
			940 => "0010000110001000000100",
			941 => "0000000000111011011001",
			942 => "0000001000111011011001",
			943 => "0011000100010100001000",
			944 => "0000011100110100000100",
			945 => "0000000000111011011001",
			946 => "0000000000111011011001",
			947 => "0011000100010100000100",
			948 => "0000000000111011011001",
			949 => "0000000000111011011001",
			950 => "0001111101111010000000",
			951 => "0001000011111001111100",
			952 => "0001110100010100111100",
			953 => "0000110000101000100000",
			954 => "0010011100110100010000",
			955 => "0000110000111000001000",
			956 => "0000101101000100000100",
			957 => "0000000000111111111101",
			958 => "0000001000111111111101",
			959 => "0001100111101000000100",
			960 => "1111111000111111111101",
			961 => "0000001000111111111101",
			962 => "0000101110101100001000",
			963 => "0000111110111100000100",
			964 => "0000000000111111111101",
			965 => "0000001000111111111101",
			966 => "0010100101000100000100",
			967 => "0000000000111111111101",
			968 => "0000001000111111111101",
			969 => "0010101001000100010000",
			970 => "0000100111100000001000",
			971 => "0010111011000100000100",
			972 => "0000000000111111111101",
			973 => "0000001000111111111101",
			974 => "0010101000010100000100",
			975 => "0000000000111111111101",
			976 => "1111111000111111111101",
			977 => "0000101110101000000100",
			978 => "0000010000111111111101",
			979 => "0010010010001100000100",
			980 => "0000001000111111111101",
			981 => "0000000000111111111101",
			982 => "0001100100110100100000",
			983 => "0000101010001000010000",
			984 => "0001110100000000001000",
			985 => "0011100101101100000100",
			986 => "0000000000111111111101",
			987 => "0000001000111111111101",
			988 => "0001001000001000000100",
			989 => "0000000000111111111101",
			990 => "1111111000111111111101",
			991 => "0010011001111000001000",
			992 => "0010001111001000000100",
			993 => "0000000000111111111101",
			994 => "0000010000111111111101",
			995 => "0010111000111100000100",
			996 => "0000000000111111111101",
			997 => "1111111000111111111101",
			998 => "0010010110101000010000",
			999 => "0011011110001100001000",
			1000 => "0000101001010000000100",
			1001 => "0000001000111111111101",
			1002 => "0000000000111111111101",
			1003 => "0010100101000100000100",
			1004 => "0000001000111111111101",
			1005 => "1111111000111111111101",
			1006 => "0000111100101100001000",
			1007 => "0010100110011000000100",
			1008 => "1111110000111111111101",
			1009 => "0000000000111111111101",
			1010 => "0010010111100100000100",
			1011 => "0000001000111111111101",
			1012 => "0000000000111111111101",
			1013 => "1111111000111111111101",
			1014 => "0010100111110100010000",
			1015 => "0011111000101000001100",
			1016 => "0001110001111100001000",
			1017 => "0001101011111100000100",
			1018 => "1111111000111111111101",
			1019 => "0000001000111111111101",
			1020 => "1111111000111111111101",
			1021 => "0000010000111111111101",
			1022 => "1111111000111111111101",
			1023 => "0011101100110010101000",
			1024 => "0011010001111101110100",
			1025 => "0011110101110101000000",
			1026 => "0011100100000000100000",
			1027 => "0011110101100100010000",
			1028 => "0000111100001000001000",
			1029 => "0010110100010100000100",
			1030 => "0000000001001000001001",
			1031 => "0000000001001000001001",
			1032 => "0010011001111000000100",
			1033 => "0000001001001000001001",
			1034 => "0000000001001000001001",
			1035 => "0000011100110100001000",
			1036 => "0011100100010100000100",
			1037 => "0000000001001000001001",
			1038 => "0000000001001000001001",
			1039 => "0011101100001000000100",
			1040 => "0000000001001000001001",
			1041 => "1111111001001000001001",
			1042 => "0001001100001100010000",
			1043 => "0011110010001000001000",
			1044 => "0001100111101000000100",
			1045 => "1111111001001000001001",
			1046 => "0000001001001000001001",
			1047 => "0001111100001000000100",
			1048 => "0000000001001000001001",
			1049 => "1111111001001000001001",
			1050 => "0011000000101000001000",
			1051 => "0001110100000000000100",
			1052 => "0000001001001000001001",
			1053 => "1111111001001000001001",
			1054 => "0010111000111000000100",
			1055 => "0000001001001000001001",
			1056 => "0000000001001000001001",
			1057 => "0011000000101000100000",
			1058 => "0011001110111100010000",
			1059 => "0011001010000000001000",
			1060 => "0011110000110100000100",
			1061 => "0000000001001000001001",
			1062 => "0000001001001000001001",
			1063 => "0001101100011000000100",
			1064 => "0000001001001000001001",
			1065 => "0000000001001000001001",
			1066 => "0010001011010100001000",
			1067 => "0011011100101100000100",
			1068 => "1111111001001000001001",
			1069 => "0000000001001000001001",
			1070 => "0000000011010000000100",
			1071 => "0000001001001000001001",
			1072 => "0000000001001000001001",
			1073 => "0011000000101000000100",
			1074 => "0000010001001000001001",
			1075 => "0011000100000000001000",
			1076 => "0011110111110000000100",
			1077 => "0000000001001000001001",
			1078 => "1111111001001000001001",
			1079 => "0011101000111000000100",
			1080 => "0000000001001000001001",
			1081 => "0000001001001000001001",
			1082 => "0011001000111000100100",
			1083 => "0011110000110100011100",
			1084 => "0000110100001000010000",
			1085 => "0011101100001000001000",
			1086 => "0011100000101000000100",
			1087 => "0000000001001000001001",
			1088 => "0000000001001000001001",
			1089 => "0011000100000000000100",
			1090 => "1111111001001000001001",
			1091 => "1111111001001000001001",
			1092 => "0001110100000000000100",
			1093 => "0000001001001000001001",
			1094 => "0011100011011100000100",
			1095 => "0000000001001000001001",
			1096 => "1111111001001000001001",
			1097 => "0010011011101000000100",
			1098 => "0000000001001000001001",
			1099 => "0000001001001000001001",
			1100 => "0011110111110000001000",
			1101 => "0000100110100000000100",
			1102 => "0000001001001000001001",
			1103 => "1111111001001000001001",
			1104 => "0011100011011100000100",
			1105 => "0000011001001000001001",
			1106 => "0000000001001000001001",
			1107 => "0011010000001100100000",
			1108 => "0000100110010000010100",
			1109 => "0000011110100000000100",
			1110 => "1111111001001000001001",
			1111 => "0001110100010100000100",
			1112 => "0000000001001000001001",
			1113 => "0010111000111100001000",
			1114 => "0010110100000000000100",
			1115 => "0000001001001000001001",
			1116 => "0000000001001000001001",
			1117 => "0000001001001000001001",
			1118 => "0011111100100100001000",
			1119 => "0001111100001000000100",
			1120 => "0000001001001000001001",
			1121 => "1111111001001000001001",
			1122 => "1111111001001000001001",
			1123 => "0000110000001100001100",
			1124 => "0010110100000000000100",
			1125 => "0000000001001000001001",
			1126 => "0000010010001100000100",
			1127 => "1111110001001000001001",
			1128 => "0000000001001000001001",
			1129 => "0010001010101100011000",
			1130 => "0001000010100100010000",
			1131 => "0000001111000100001000",
			1132 => "0001001000110100000100",
			1133 => "0000000001001000001001",
			1134 => "1111111001001000001001",
			1135 => "0010001001101000000100",
			1136 => "0000001001001000001001",
			1137 => "0000000001001000001001",
			1138 => "0011010100001000000100",
			1139 => "0000000001001000001001",
			1140 => "1111111001001000001001",
			1141 => "0011000100000000001100",
			1142 => "0011111110101100000100",
			1143 => "0000011001001000001001",
			1144 => "0011111100100100000100",
			1145 => "0000000001001000001001",
			1146 => "0000001001001000001001",
			1147 => "0011100110100100001000",
			1148 => "0001111000111000000100",
			1149 => "0000000001001000001001",
			1150 => "1111111001001000001001",
			1151 => "0001101000010000000100",
			1152 => "0000001001001000001001",
			1153 => "0000000001001000001001",
			1154 => "0011000110000110101100",
			1155 => "0010011001111001011000",
			1156 => "0000111000111100111100",
			1157 => "0010000110001000100000",
			1158 => "0001000010111000010000",
			1159 => "0011000111111000001000",
			1160 => "0010001011010100000100",
			1161 => "0000001001001101110101",
			1162 => "0000000001001101110101",
			1163 => "0011100011010000000100",
			1164 => "1111111001001101110101",
			1165 => "0000000001001101110101",
			1166 => "0001011001110000001000",
			1167 => "0000101110101000000100",
			1168 => "0000000001001101110101",
			1169 => "1111111001001101110101",
			1170 => "0001010011011100000100",
			1171 => "0000010001001101110101",
			1172 => "0000000001001101110101",
			1173 => "0001011100110000010000",
			1174 => "0010010010001100001000",
			1175 => "0000111010000000000100",
			1176 => "0000000001001101110101",
			1177 => "0000000001001101110101",
			1178 => "0010001111001000000100",
			1179 => "1111111001001101110101",
			1180 => "0000000001001101110101",
			1181 => "0010000010101000000100",
			1182 => "0000011001001101110101",
			1183 => "0011011100101100000100",
			1184 => "0000000001001101110101",
			1185 => "0000001001001101110101",
			1186 => "0010111100001000011000",
			1187 => "0000100010011100001100",
			1188 => "0000000010011000000100",
			1189 => "1111111001001101110101",
			1190 => "0010000110001000000100",
			1191 => "0000010001001101110101",
			1192 => "0000001001001101110101",
			1193 => "0000000000111000000100",
			1194 => "1111111001001101110101",
			1195 => "0001011100110000000100",
			1196 => "0000000001001101110101",
			1197 => "0000001001001101110101",
			1198 => "1111111001001101110101",
			1199 => "0000011110100000011000",
			1200 => "0001010011011100000100",
			1201 => "0000000001001101110101",
			1202 => "0000011110100000001000",
			1203 => "0011100111111000000100",
			1204 => "1111111001001101110101",
			1205 => "1111110001001101110101",
			1206 => "0011100100010100001000",
			1207 => "0000000100010100000100",
			1208 => "1111111001001101110101",
			1209 => "0000000001001101110101",
			1210 => "0000000001001101110101",
			1211 => "0011000111111000100000",
			1212 => "0010011001111000010000",
			1213 => "0001011101100000001000",
			1214 => "0011000111111000000100",
			1215 => "0000000001001101110101",
			1216 => "1111111001001101110101",
			1217 => "0010001111001000000100",
			1218 => "0000001001001101110101",
			1219 => "0000001001001101110101",
			1220 => "0000100011001000001000",
			1221 => "0000100100101000000100",
			1222 => "0000000001001101110101",
			1223 => "0000000001001101110101",
			1224 => "0001011101100000000100",
			1225 => "0000001001001101110101",
			1226 => "0000000001001101110101",
			1227 => "0011000100010100010000",
			1228 => "0001011110001100001000",
			1229 => "0010010110101000000100",
			1230 => "0000000001001101110101",
			1231 => "0000001001001101110101",
			1232 => "0010111000111100000100",
			1233 => "1111111001001101110101",
			1234 => "0000001001001101110101",
			1235 => "0001010011011100000100",
			1236 => "0000001001001101110101",
			1237 => "0010111011000100000100",
			1238 => "1111111001001101110101",
			1239 => "0000000001001101110101",
			1240 => "0010100111110100001000",
			1241 => "0000100001011100000100",
			1242 => "1111111001001101110101",
			1243 => "0000001001001101110101",
			1244 => "1111111001001101110101",
			1245 => "0010001001101010001100",
			1246 => "0010001001101001000000",
			1247 => "0011010101101100100100",
			1248 => "0001110100010100010100",
			1249 => "0001100001111000010000",
			1250 => "0011101110111100001000",
			1251 => "0010110100010100000100",
			1252 => "0000000001010110100001",
			1253 => "1111111001010110100001",
			1254 => "0001001110000000000100",
			1255 => "0000000001010110100001",
			1256 => "0000001001010110100001",
			1257 => "1111111001010110100001",
			1258 => "0000101101000100001100",
			1259 => "0000110100010100000100",
			1260 => "0000000001010110100001",
			1261 => "0000100010110100000100",
			1262 => "0000001001010110100001",
			1263 => "0000001001010110100001",
			1264 => "0000000001010110100001",
			1265 => "0011100000110000000100",
			1266 => "1111111001010110100001",
			1267 => "0001110100010100001000",
			1268 => "0000011110100000000100",
			1269 => "0000000001010110100001",
			1270 => "0000001001010110100001",
			1271 => "0010110000101000001000",
			1272 => "0001000110001100000100",
			1273 => "1111111001010110100001",
			1274 => "0000000001010110100001",
			1275 => "0001011100101100000100",
			1276 => "0000000001010110100001",
			1277 => "0000000001010110100001",
			1278 => "0000100010011100101000",
			1279 => "0010101000010100010000",
			1280 => "0010101000010100000100",
			1281 => "0000000001010110100001",
			1282 => "0001100001111000001000",
			1283 => "0010111100001000000100",
			1284 => "1111111001010110100001",
			1285 => "0000000001010110100001",
			1286 => "1111111001010110100001",
			1287 => "0000011110100000001000",
			1288 => "0010011001111000000100",
			1289 => "0000000001010110100001",
			1290 => "1111111001010110100001",
			1291 => "0001011101111000001000",
			1292 => "0011000000101000000100",
			1293 => "0000000001010110100001",
			1294 => "0000001001010110100001",
			1295 => "0001010000001100000100",
			1296 => "1111111001010110100001",
			1297 => "0000000001010110100001",
			1298 => "0010110100010100001000",
			1299 => "0011000000111000000100",
			1300 => "0000000001010110100001",
			1301 => "0000001001010110100001",
			1302 => "0000011100110100001100",
			1303 => "0001111011000100000100",
			1304 => "1111111001010110100001",
			1305 => "0011101000111100000100",
			1306 => "1111111001010110100001",
			1307 => "0000000001010110100001",
			1308 => "0011010000001100001000",
			1309 => "0000011100110100000100",
			1310 => "0000000001010110100001",
			1311 => "0000001001010110100001",
			1312 => "0000011001111000000100",
			1313 => "1111111001010110100001",
			1314 => "0000000001010110100001",
			1315 => "0010001011010100110100",
			1316 => "0001101010011000101000",
			1317 => "0001001000001000010100",
			1318 => "0011011110001100001100",
			1319 => "0010110000101000000100",
			1320 => "0000001001010110100001",
			1321 => "0001000110001100000100",
			1322 => "0000001001010110100001",
			1323 => "1111111001010110100001",
			1324 => "0000101010001000000100",
			1325 => "0000001001010110100001",
			1326 => "0000001001010110100001",
			1327 => "0000100101110000001100",
			1328 => "0001000011001100000100",
			1329 => "0000000001010110100001",
			1330 => "0001100001111000000100",
			1331 => "0000000001010110100001",
			1332 => "0000001001010110100001",
			1333 => "0001110100010100000100",
			1334 => "0000001001010110100001",
			1335 => "1111111001010110100001",
			1336 => "0000101111010100000100",
			1337 => "1111111001010110100001",
			1338 => "0000111101000100000100",
			1339 => "0000001001010110100001",
			1340 => "0000000001010110100001",
			1341 => "0001010100011001000000",
			1342 => "0010011011101000100000",
			1343 => "0000010010001100010000",
			1344 => "0000100010000000001000",
			1345 => "0000111101111000000100",
			1346 => "0000000001010110100001",
			1347 => "0000000001010110100001",
			1348 => "0001110100000000000100",
			1349 => "0000000001010110100001",
			1350 => "0000000001010110100001",
			1351 => "0010110100000000001000",
			1352 => "0010011101101000000100",
			1353 => "1111111001010110100001",
			1354 => "0000000001010110100001",
			1355 => "0010011101101000000100",
			1356 => "0000001001010110100001",
			1357 => "0000000001010110100001",
			1358 => "0011101101010100010000",
			1359 => "0011001000111000001000",
			1360 => "0010001011010100000100",
			1361 => "1111111001010110100001",
			1362 => "0000000001010110100001",
			1363 => "0001001110111000000100",
			1364 => "0000001001010110100001",
			1365 => "1111111001010110100001",
			1366 => "0010011111001100001000",
			1367 => "0001101010011000000100",
			1368 => "0000000001010110100001",
			1369 => "0000001001010110100001",
			1370 => "0010100001010000000100",
			1371 => "0000000001010110100001",
			1372 => "0000000001010110100001",
			1373 => "0001000010100100010100",
			1374 => "0011101101010100000100",
			1375 => "0000010001010110100001",
			1376 => "0001001000001000001000",
			1377 => "0001111001110000000100",
			1378 => "0000001001010110100001",
			1379 => "0000000001010110100001",
			1380 => "0011000100000000000100",
			1381 => "0000000001010110100001",
			1382 => "0000001001010110100001",
			1383 => "1111111001010110100001",
			1384 => "0001010011100010110000",
			1385 => "0001000011010101100000",
			1386 => "0011100100010100110000",
			1387 => "0011101010000000010100",
			1388 => "0001000111010100000100",
			1389 => "0000011001011101110101",
			1390 => "0001101101111100001000",
			1391 => "0010110100010100000100",
			1392 => "0000001001011101110101",
			1393 => "0000000001011101110101",
			1394 => "0000000100010100000100",
			1395 => "0000010001011101110101",
			1396 => "1111111001011101110101",
			1397 => "0010001100000100001100",
			1398 => "0001100001111000001000",
			1399 => "0001010101101100000100",
			1400 => "0000000001011101110101",
			1401 => "1111111001011101110101",
			1402 => "0000010001011101110101",
			1403 => "0000101110101000001000",
			1404 => "0000000010111100000100",
			1405 => "0000001001011101110101",
			1406 => "0000100001011101110101",
			1407 => "0010011001111000000100",
			1408 => "0000010001011101110101",
			1409 => "0000001001011101110101",
			1410 => "0001100111101000010000",
			1411 => "0010000001010100001100",
			1412 => "0000111101100000000100",
			1413 => "0000000001011101110101",
			1414 => "0011000111111000000100",
			1415 => "1111111001011101110101",
			1416 => "1111111001011101110101",
			1417 => "0000001001011101110101",
			1418 => "0001001010110100010000",
			1419 => "0001101001100100001000",
			1420 => "0001101101111100000100",
			1421 => "0000001001011101110101",
			1422 => "0000010001011101110101",
			1423 => "0010101100011100000100",
			1424 => "1111111001011101110101",
			1425 => "0000001001011101110101",
			1426 => "0011000100000000001000",
			1427 => "0011101100110000000100",
			1428 => "0000001001011101110101",
			1429 => "0000010001011101110101",
			1430 => "0000101100010000000100",
			1431 => "0000000001011101110101",
			1432 => "0000001001011101110101",
			1433 => "0001101101111100010100",
			1434 => "0001000011110100000100",
			1435 => "0000001001011101110101",
			1436 => "0000010000011000000100",
			1437 => "1111111001011101110101",
			1438 => "0010010010001100001000",
			1439 => "0001000011101100000100",
			1440 => "1111111001011101110101",
			1441 => "0000000001011101110101",
			1442 => "1111111001011101110101",
			1443 => "0010111100001000100000",
			1444 => "0000001011000100010000",
			1445 => "0011000111111000001000",
			1446 => "0001000011110100000100",
			1447 => "0000010001011101110101",
			1448 => "0000100001011101110101",
			1449 => "0001010101101100000100",
			1450 => "0000001001011101110101",
			1451 => "0000000001011101110101",
			1452 => "0001000001101100001000",
			1453 => "0010011100110100000100",
			1454 => "0000010001011101110101",
			1455 => "0000000001011101110101",
			1456 => "0010101100000100000100",
			1457 => "0000010001011101110101",
			1458 => "1111111001011101110101",
			1459 => "0011111100100100010000",
			1460 => "0000101001011100001000",
			1461 => "0000110101101100000100",
			1462 => "0000000001011101110101",
			1463 => "0000010001011101110101",
			1464 => "0011000111111000000100",
			1465 => "0000001001011101110101",
			1466 => "1111111001011101110101",
			1467 => "0000000100010100000100",
			1468 => "1111111001011101110101",
			1469 => "0001000011101100000100",
			1470 => "0000010001011101110101",
			1471 => "0000000001011101110101",
			1472 => "0011000110000100100100",
			1473 => "0001010100010000100000",
			1474 => "0000111000011000000100",
			1475 => "1111111001011101110101",
			1476 => "0001101101011000001100",
			1477 => "0001100001111000000100",
			1478 => "1111111001011101110101",
			1479 => "0000101100010100000100",
			1480 => "0000011001011101110101",
			1481 => "0000001001011101110101",
			1482 => "0001101001100100001000",
			1483 => "0000101100010000000100",
			1484 => "1111111001011101110101",
			1485 => "0000000001011101110101",
			1486 => "0011001100001000000100",
			1487 => "0000000001011101110101",
			1488 => "1111111001011101110101",
			1489 => "0000011001011101110101",
			1490 => "0011000110000100010100",
			1491 => "0010001111001000010000",
			1492 => "0010000110001000001100",
			1493 => "0010000110011100000100",
			1494 => "1111111001011101110101",
			1495 => "0010001100000100000100",
			1496 => "0000000001011101110101",
			1497 => "1111111001011101110101",
			1498 => "0000001001011101110101",
			1499 => "1111111001011101110101",
			1500 => "1111111001011101110101",
			1501 => "0000101100010110001100",
			1502 => "0001000011011001100000",
			1503 => "0001101010011001000000",
			1504 => "0001101100011000100000",
			1505 => "0001101100011000010000",
			1506 => "0000101110101000001000",
			1507 => "0001100001111000000100",
			1508 => "0000000001100110011001",
			1509 => "0000000001100110011001",
			1510 => "0001101101111100000100",
			1511 => "0000000001100110011001",
			1512 => "0000000001100110011001",
			1513 => "0001000011001100001000",
			1514 => "0000011100110100000100",
			1515 => "1111111001100110011001",
			1516 => "0000000001100110011001",
			1517 => "0010001111001000000100",
			1518 => "1111111001100110011001",
			1519 => "0000000001100110011001",
			1520 => "0000111101111000010000",
			1521 => "0000011100110100001000",
			1522 => "0000111100101100000100",
			1523 => "0000000001100110011001",
			1524 => "0000001001100110011001",
			1525 => "0010000001110100000100",
			1526 => "1111111001100110011001",
			1527 => "0000000001100110011001",
			1528 => "0011000100000000001000",
			1529 => "0011101001110000000100",
			1530 => "0000000001100110011001",
			1531 => "0000001001100110011001",
			1532 => "0001101010011000000100",
			1533 => "0000000001100110011001",
			1534 => "1111111001100110011001",
			1535 => "0010001011010100001100",
			1536 => "0011001000111000001000",
			1537 => "0010001001101000000100",
			1538 => "0000000001100110011001",
			1539 => "1111110001100110011001",
			1540 => "0000000001100110011001",
			1541 => "0010100001010000000100",
			1542 => "0000010001100110011001",
			1543 => "0001110100000000001000",
			1544 => "0000100011001000000100",
			1545 => "0000000001100110011001",
			1546 => "0000001001100110011001",
			1547 => "0011011100101000000100",
			1548 => "0000001001100110011001",
			1549 => "1111111001100110011001",
			1550 => "0000011110100000100100",
			1551 => "0011010110000100011100",
			1552 => "0000001100110000010000",
			1553 => "0000111110111100001000",
			1554 => "0010100101000100000100",
			1555 => "0000000001100110011001",
			1556 => "0000001001100110011001",
			1557 => "0001100001111000000100",
			1558 => "0000000001100110011001",
			1559 => "0000010001100110011001",
			1560 => "0001000110110000000100",
			1561 => "1111111001100110011001",
			1562 => "0001000011111000000100",
			1563 => "0000001001100110011001",
			1564 => "1111111001100110011001",
			1565 => "0011100011111100000100",
			1566 => "1111111001100110011001",
			1567 => "0000000001100110011001",
			1568 => "0011000000101000000100",
			1569 => "0000011001100110011001",
			1570 => "1111111001100110011001",
			1571 => "0001101100011001001100",
			1572 => "0011111110101000101000",
			1573 => "0011101101111000100000",
			1574 => "0000000000110000010000",
			1575 => "0010110000101000001000",
			1576 => "0011001010000000000100",
			1577 => "0000000001100110011001",
			1578 => "0000000001100110011001",
			1579 => "0001111100001000000100",
			1580 => "1111111001100110011001",
			1581 => "1111111001100110011001",
			1582 => "0001111100001000001000",
			1583 => "0011011100101100000100",
			1584 => "0000000001100110011001",
			1585 => "0000001001100110011001",
			1586 => "0001110100000000000100",
			1587 => "1111111001100110011001",
			1588 => "0000000001100110011001",
			1589 => "0000010010001100000100",
			1590 => "0000001001100110011001",
			1591 => "0000000001100110011001",
			1592 => "0011100011011100000100",
			1593 => "0000010001100110011001",
			1594 => "0011011010111000010000",
			1595 => "0011000000101000001000",
			1596 => "0010001100000100000100",
			1597 => "0000001001100110011001",
			1598 => "1111111001100110011001",
			1599 => "0000000000110000000100",
			1600 => "1111110001100110011001",
			1601 => "1111111001100110011001",
			1602 => "0001101100011000001000",
			1603 => "0001000001011100000100",
			1604 => "0000000001100110011001",
			1605 => "1111111001100110011001",
			1606 => "0000101110110100000100",
			1607 => "0000001001100110011001",
			1608 => "0000000001100110011001",
			1609 => "0001101111000000110000",
			1610 => "0011110000110100010000",
			1611 => "0001101010011000001000",
			1612 => "0000111110001100000100",
			1613 => "1111111001100110011001",
			1614 => "0000001001100110011001",
			1615 => "0000010010001100000100",
			1616 => "1111111001100110011001",
			1617 => "0000000001100110011001",
			1618 => "0010001111001000010000",
			1619 => "0001001000001000001000",
			1620 => "0011011010111000000100",
			1621 => "0000001001100110011001",
			1622 => "0000000001100110011001",
			1623 => "0000100010000000000100",
			1624 => "0000000001100110011001",
			1625 => "1111111001100110011001",
			1626 => "0001001110111000001000",
			1627 => "0011110101110000000100",
			1628 => "0000000001100110011001",
			1629 => "0000001001100110011001",
			1630 => "0000001110111100000100",
			1631 => "0000000001100110011001",
			1632 => "0000000001100110011001",
			1633 => "0011011011000000001000",
			1634 => "0000101111010100000100",
			1635 => "0000000001100110011001",
			1636 => "0000001001100110011001",
			1637 => "1111111001100110011001",
			1638 => "0011000100000010101100",
			1639 => "0011000000101001110000",
			1640 => "0000100110010000111000",
			1641 => "0000010010001100100000",
			1642 => "0001111100001000010000",
			1643 => "0001110000101000001000",
			1644 => "0001110000101000000100",
			1645 => "0000000001110000001101",
			1646 => "0000000001110000001101",
			1647 => "0011101101111000000100",
			1648 => "0000000001110000001101",
			1649 => "0000001001110000001101",
			1650 => "0001111100001000001000",
			1651 => "0010101100011100000100",
			1652 => "1111111001110000001101",
			1653 => "0000000001110000001101",
			1654 => "0010000001110100000100",
			1655 => "0000000001110000001101",
			1656 => "0000000001110000001101",
			1657 => "0010011101011100010000",
			1658 => "0001111000111000001000",
			1659 => "0001001000101000000100",
			1660 => "0000000001110000001101",
			1661 => "0000001001110000001101",
			1662 => "0010100001010000000100",
			1663 => "1111111001110000001101",
			1664 => "0000000001110000001101",
			1665 => "0011101000000000000100",
			1666 => "1111111001110000001101",
			1667 => "0000000001110000001101",
			1668 => "0010011101101000100000",
			1669 => "0011111101000100010000",
			1670 => "0010101100011100001000",
			1671 => "0010000110001000000100",
			1672 => "0000000001110000001101",
			1673 => "1111111001110000001101",
			1674 => "0011101000111100000100",
			1675 => "1111111001110000001101",
			1676 => "0000000001110000001101",
			1677 => "0011111110000100001000",
			1678 => "0011000100010100000100",
			1679 => "0000000001110000001101",
			1680 => "0000001001110000001101",
			1681 => "0011110010011100000100",
			1682 => "1111111001110000001101",
			1683 => "0000000001110000001101",
			1684 => "0001000010110000001000",
			1685 => "0001000110001100000100",
			1686 => "1111111001110000001101",
			1687 => "0000001001110000001101",
			1688 => "0010000111000100001000",
			1689 => "0000011001111000000100",
			1690 => "1111111001110000001101",
			1691 => "0000000001110000001101",
			1692 => "0001000100001100000100",
			1693 => "0000000001110000001101",
			1694 => "1111111001110000001101",
			1695 => "0011000000101000011000",
			1696 => "0001001101001000001100",
			1697 => "0000110000001100000100",
			1698 => "1111111001110000001101",
			1699 => "0011100001111100000100",
			1700 => "0000001001110000001101",
			1701 => "0000000001110000001101",
			1702 => "0010111000111000001000",
			1703 => "0010000001110100000100",
			1704 => "0000010001110000001101",
			1705 => "0000001001110000001101",
			1706 => "0000000001110000001101",
			1707 => "0010000001110000010000",
			1708 => "0010100111110100001000",
			1709 => "0010011111001100000100",
			1710 => "1111111001110000001101",
			1711 => "0000001001110000001101",
			1712 => "0000010010001100000100",
			1713 => "0000001001110000001101",
			1714 => "0000001001110000001101",
			1715 => "0010101000010100001000",
			1716 => "0010101000100100000100",
			1717 => "0000000001110000001101",
			1718 => "1111110001110000001101",
			1719 => "0010101000010100000100",
			1720 => "0000001001110000001101",
			1721 => "0010001011010100000100",
			1722 => "0000000001110000001101",
			1723 => "0000000001110000001101",
			1724 => "0011000100000000111000",
			1725 => "0001110100000000001100",
			1726 => "0001110100000000000100",
			1727 => "1111111001110000001101",
			1728 => "0011110001001000000100",
			1729 => "0000000001110000001101",
			1730 => "0000001001110000001101",
			1731 => "0000011001111000011000",
			1732 => "0000100110010000010000",
			1733 => "0010011101101000001000",
			1734 => "0010111000111000000100",
			1735 => "1111111001110000001101",
			1736 => "1111110001110000001101",
			1737 => "0000010010001100000100",
			1738 => "0000000001110000001101",
			1739 => "1111111001110000001101",
			1740 => "0001011100101000000100",
			1741 => "1111111001110000001101",
			1742 => "0000000001110000001101",
			1743 => "0011101110110000001000",
			1744 => "0001111001110000000100",
			1745 => "0000001001110000001101",
			1746 => "0000000001110000001101",
			1747 => "0011111001011100001000",
			1748 => "0000000010011000000100",
			1749 => "1111110001110000001101",
			1750 => "1111111001110000001101",
			1751 => "0000000001110000001101",
			1752 => "0011000100000000011100",
			1753 => "0001010000001100001000",
			1754 => "0001011101111000000100",
			1755 => "0000001001110000001101",
			1756 => "0000001001110000001101",
			1757 => "0001010100001000000100",
			1758 => "1111111001110000001101",
			1759 => "0001011010111000001000",
			1760 => "0011101100101000000100",
			1761 => "0000000001110000001101",
			1762 => "0000001001110000001101",
			1763 => "0011110100101000000100",
			1764 => "1111111001110000001101",
			1765 => "0000000001110000001101",
			1766 => "0011001000111100011100",
			1767 => "0011001000111100010000",
			1768 => "0011101010111000001000",
			1769 => "0001111000111000000100",
			1770 => "0000000001110000001101",
			1771 => "1111111001110000001101",
			1772 => "0000100110010000000100",
			1773 => "0000001001110000001101",
			1774 => "1111111001110000001101",
			1775 => "0011101110001100000100",
			1776 => "0000000001110000001101",
			1777 => "0000101100000000000100",
			1778 => "1111111001110000001101",
			1779 => "0000000001110000001101",
			1780 => "0011001000111000010000",
			1781 => "0000110001011000001000",
			1782 => "0011100000001100000100",
			1783 => "0000000001110000001101",
			1784 => "0000001001110000001101",
			1785 => "0000011101101000000100",
			1786 => "1111111001110000001101",
			1787 => "0000001001110000001101",
			1788 => "0011001000111000001000",
			1789 => "0000101000001100000100",
			1790 => "1111111001110000001101",
			1791 => "0000001001110000001101",
			1792 => "0001011101010100000100",
			1793 => "0000000001110000001101",
			1794 => "0000000001110000001101",
			1795 => "0011001000111011011100",
			1796 => "0011000111111001110100",
			1797 => "0010010110101001000000",
			1798 => "0000111001110000100000",
			1799 => "0010011001111000010000",
			1800 => "0000111011000100001000",
			1801 => "0011110111010000000100",
			1802 => "0000000001111001011001",
			1803 => "1111111001111001011001",
			1804 => "0001010011011100000100",
			1805 => "0000000001111001011001",
			1806 => "0000000001111001011001",
			1807 => "0001000011110000001000",
			1808 => "0011100000110000000100",
			1809 => "0000000001111001011001",
			1810 => "0000001001111001011001",
			1811 => "0010100001010000000100",
			1812 => "1111111001111001011001",
			1813 => "0000000001111001011001",
			1814 => "0011110010001000010000",
			1815 => "0011100100010100001000",
			1816 => "0001110100010100000100",
			1817 => "0000000001111001011001",
			1818 => "0000001001111001011001",
			1819 => "0001100111101000000100",
			1820 => "0000000001111001011001",
			1821 => "0000001001111001011001",
			1822 => "0010100001010000001000",
			1823 => "0011100100000000000100",
			1824 => "1111111001111001011001",
			1825 => "0000000001111001011001",
			1826 => "0010101100011100000100",
			1827 => "0000001001111001011001",
			1828 => "1111111001111001011001",
			1829 => "0001011100110000010100",
			1830 => "0010110000101000001100",
			1831 => "0011000111111000001000",
			1832 => "0011100000101000000100",
			1833 => "1111111001111001011001",
			1834 => "0000000001111001011001",
			1835 => "0000000001111001011001",
			1836 => "0010010110101000000100",
			1837 => "1111111001111001011001",
			1838 => "1111110001111001011001",
			1839 => "0010101001000100010000",
			1840 => "0001001000110100001000",
			1841 => "0010101000100100000100",
			1842 => "0000000001111001011001",
			1843 => "0000001001111001011001",
			1844 => "0000100101001000000100",
			1845 => "1111111001111001011001",
			1846 => "0000000001111001011001",
			1847 => "0011000111111000001000",
			1848 => "0001011100101100000100",
			1849 => "0000001001111001011001",
			1850 => "1111111001111001011001",
			1851 => "0000100010011100000100",
			1852 => "0000000001111001011001",
			1853 => "0000000001111001011001",
			1854 => "0011000100010100101000",
			1855 => "0001001000001000010100",
			1856 => "0011000111111000001100",
			1857 => "0001110100010100000100",
			1858 => "0000001001111001011001",
			1859 => "0001111100001000000100",
			1860 => "1111111001111001011001",
			1861 => "0000000001111001011001",
			1862 => "0010010110101000000100",
			1863 => "0000000001111001011001",
			1864 => "0000001001111001011001",
			1865 => "0010111110111100000100",
			1866 => "1111111001111001011001",
			1867 => "0000100011001000001000",
			1868 => "0011100100010100000100",
			1869 => "0000001001111001011001",
			1870 => "0000001001111001011001",
			1871 => "0011101001110000000100",
			1872 => "1111111001111001011001",
			1873 => "0000001001111001011001",
			1874 => "0000111100110000100000",
			1875 => "0010010110101000010000",
			1876 => "0011011110001100001000",
			1877 => "0001010110000100000100",
			1878 => "0000000001111001011001",
			1879 => "1111111001111001011001",
			1880 => "0011110101100100000100",
			1881 => "0000001001111001011001",
			1882 => "1111111001111001011001",
			1883 => "0011110100000100001000",
			1884 => "0000111001110000000100",
			1885 => "1111111001111001011001",
			1886 => "0000000001111001011001",
			1887 => "0000101001010000000100",
			1888 => "1111111001111001011001",
			1889 => "0000000001111001011001",
			1890 => "0010010111100100010000",
			1891 => "0011000100010100001000",
			1892 => "0011010000001100000100",
			1893 => "0000000001111001011001",
			1894 => "1111111001111001011001",
			1895 => "0001010101101100000100",
			1896 => "0000001001111001011001",
			1897 => "0000000001111001011001",
			1898 => "0011101000111100001000",
			1899 => "0010100001010000000100",
			1900 => "0000000001111001011001",
			1901 => "1111111001111001011001",
			1902 => "0011111010010100000100",
			1903 => "0000000001111001011001",
			1904 => "0000000001111001011001",
			1905 => "0011111101000100011000",
			1906 => "0001011000000000001100",
			1907 => "0011100110000100001000",
			1908 => "0001001010110100000100",
			1909 => "0000001001111001011001",
			1910 => "1111111001111001011001",
			1911 => "1111111001111001011001",
			1912 => "0001011000000000001000",
			1913 => "0001101100011000000100",
			1914 => "0000000001111001011001",
			1915 => "0000010001111001011001",
			1916 => "1111111001111001011001",
			1917 => "0001101101011000011000",
			1918 => "0001001000001000010100",
			1919 => "0000100011001000001000",
			1920 => "0001110100001000000100",
			1921 => "0000001001111001011001",
			1922 => "0000000001111001011001",
			1923 => "0010011001100100000100",
			1924 => "1111111001111001011001",
			1925 => "0010100010101100000100",
			1926 => "0000000001111001011001",
			1927 => "0000001001111001011001",
			1928 => "0000001001111001011001",
			1929 => "0010100110011100010000",
			1930 => "0010111101111000000100",
			1931 => "1111111001111001011001",
			1932 => "0010010101011100000100",
			1933 => "0000001001111001011001",
			1934 => "0000101100000000000100",
			1935 => "0000000001111001011001",
			1936 => "1111111001111001011001",
			1937 => "0011110010011100001000",
			1938 => "0001110101101100000100",
			1939 => "0000010001111001011001",
			1940 => "0000000001111001011001",
			1941 => "1111111001111001011001",
			1942 => "0010011001111010001000",
			1943 => "0001011101100001001000",
			1944 => "0001010011011101000000",
			1945 => "0000101001010000100000",
			1946 => "0000110100010100010000",
			1947 => "0010111011000100001000",
			1948 => "0010100101000100000100",
			1949 => "0000000010000010111101",
			1950 => "0000001010000010111101",
			1951 => "0001100001111000000100",
			1952 => "0000000010000010111101",
			1953 => "1111111010000010111101",
			1954 => "0001110111111000001000",
			1955 => "0000111100001000000100",
			1956 => "1111111010000010111101",
			1957 => "0000000010000010111101",
			1958 => "0010110100010100000100",
			1959 => "0000001010000010111101",
			1960 => "0000000010000010111101",
			1961 => "0000010110000000010000",
			1962 => "0000111100001000001000",
			1963 => "0011001010000000000100",
			1964 => "0000000010000010111101",
			1965 => "1111111010000010111101",
			1966 => "0000111100001000000100",
			1967 => "0000001010000010111101",
			1968 => "0000000010000010111101",
			1969 => "0010110100010100001000",
			1970 => "0010000001110100000100",
			1971 => "1111111010000010111101",
			1972 => "0000000010000010111101",
			1973 => "0011000111111000000100",
			1974 => "0000000010000010111101",
			1975 => "1111111010000010111101",
			1976 => "0011110110100100000100",
			1977 => "0000000010000010111101",
			1978 => "1111111010000010111101",
			1979 => "0001101101111100100100",
			1980 => "0011011101100000001100",
			1981 => "0011000100010100001000",
			1982 => "0010001011010100000100",
			1983 => "0000001010000010111101",
			1984 => "1111111010000010111101",
			1985 => "0000001010000010111101",
			1986 => "0000010110000000010000",
			1987 => "0010001011010100001000",
			1988 => "0000100110100000000100",
			1989 => "0000000010000010111101",
			1990 => "0000001010000010111101",
			1991 => "0000100010000000000100",
			1992 => "1111111010000010111101",
			1993 => "0000000010000010111101",
			1994 => "0010111011000100000100",
			1995 => "1111111010000010111101",
			1996 => "0000000010000010111101",
			1997 => "0001111100001000011000",
			1998 => "0011100000111000001100",
			1999 => "0011110101100100001000",
			2000 => "0000101110000100000100",
			2001 => "0000000010000010111101",
			2002 => "0000001010000010111101",
			2003 => "1111111010000010111101",
			2004 => "0011011101100000000100",
			2005 => "0000000010000010111101",
			2006 => "0011010101101100000100",
			2007 => "0000001010000010111101",
			2008 => "0000001010000010111101",
			2009 => "1111111010000010111101",
			2010 => "0000110101101101001100",
			2011 => "0000110101101100110100",
			2012 => "0000111100110000100000",
			2013 => "0010010111100100010000",
			2014 => "0011000111111000001000",
			2015 => "0010110000101000000100",
			2016 => "0000000010000010111101",
			2017 => "1111111010000010111101",
			2018 => "0011000100010100000100",
			2019 => "0000000010000010111101",
			2020 => "0000000010000010111101",
			2021 => "0010010111100100001000",
			2022 => "0010101010110000000100",
			2023 => "1111111010000010111101",
			2024 => "0000000010000010111101",
			2025 => "0011111011011100000100",
			2026 => "0000000010000010111101",
			2027 => "1111111010000010111101",
			2028 => "0001100100110100001100",
			2029 => "0011000100010100001000",
			2030 => "0011000100010100000100",
			2031 => "0000000010000010111101",
			2032 => "1111111010000010111101",
			2033 => "0000001010000010111101",
			2034 => "0000101110010000000100",
			2035 => "0000001010000010111101",
			2036 => "0000000010000010111101",
			2037 => "0010100110011000001000",
			2038 => "0001100001111000000100",
			2039 => "1111111010000010111101",
			2040 => "0000000010000010111101",
			2041 => "0010101010110000001000",
			2042 => "0010111100001000000100",
			2043 => "1111111010000010111101",
			2044 => "1111111010000010111101",
			2045 => "0000101001011100000100",
			2046 => "0000000010000010111101",
			2047 => "1111111010000010111101",
			2048 => "0010010110101000110000",
			2049 => "0011110101110100010100",
			2050 => "0010101000010100001000",
			2051 => "0011111011011100000100",
			2052 => "0000000010000010111101",
			2053 => "0000000010000010111101",
			2054 => "0010010110101000000100",
			2055 => "0000000010000010111101",
			2056 => "0010111100001000000100",
			2057 => "0000001010000010111101",
			2058 => "0000001010000010111101",
			2059 => "0001011100101100010000",
			2060 => "0011000111111000001000",
			2061 => "0000111100101100000100",
			2062 => "0000001010000010111101",
			2063 => "0000000010000010111101",
			2064 => "0011000100010100000100",
			2065 => "0000000010000010111101",
			2066 => "0000001010000010111101",
			2067 => "0010010110101000000100",
			2068 => "0000000010000010111101",
			2069 => "0011101000111000000100",
			2070 => "1111111010000010111101",
			2071 => "0000000010000010111101",
			2072 => "0011000111111000010100",
			2073 => "0010010110101000000100",
			2074 => "1111111010000010111101",
			2075 => "0011111010010100001000",
			2076 => "0011011110001100000100",
			2077 => "0000001010000010111101",
			2078 => "0000000010000010111101",
			2079 => "0000101110010000000100",
			2080 => "1111111010000010111101",
			2081 => "0000000010000010111101",
			2082 => "0011000111111000001100",
			2083 => "0001111011000100000100",
			2084 => "0000000010000010111101",
			2085 => "0001011110001100000100",
			2086 => "0000000010000010111101",
			2087 => "0000001010000010111101",
			2088 => "0000111100101100001000",
			2089 => "0000111100101100000100",
			2090 => "0000000010000010111101",
			2091 => "1111111010000010111101",
			2092 => "0010010111100100000100",
			2093 => "0000000010000010111101",
			2094 => "0000000010000010111101",
			2095 => "0011100101101110100100",
			2096 => "0011110101100101010100",
			2097 => "0001100111101000100100",
			2098 => "0011011100101100011000",
			2099 => "0000111000111000010000",
			2100 => "0001100111101000001000",
			2101 => "0011011100110000000100",
			2102 => "0000001010001101000001",
			2103 => "0000000010001101000001",
			2104 => "0001110111111000000100",
			2105 => "0000001010001101000001",
			2106 => "1111111010001101000001",
			2107 => "0011101110111100000100",
			2108 => "0000000010001101000001",
			2109 => "0000001010001101000001",
			2110 => "0011101000111000000100",
			2111 => "1111111010001101000001",
			2112 => "0011100011011100000100",
			2113 => "0000000010001101000001",
			2114 => "0000000010001101000001",
			2115 => "0000110101101100100000",
			2116 => "0000100010110100010000",
			2117 => "0000100000110100001000",
			2118 => "0001110100010100000100",
			2119 => "1111111010001101000001",
			2120 => "0000000010001101000001",
			2121 => "0011111001001000000100",
			2122 => "0000000010001101000001",
			2123 => "0000001010001101000001",
			2124 => "0010010111100100001000",
			2125 => "0000111101100000000100",
			2126 => "0000000010001101000001",
			2127 => "0000001010001101000001",
			2128 => "0011110100000100000100",
			2129 => "0000000010001101000001",
			2130 => "1111111010001101000001",
			2131 => "0011010001111100001100",
			2132 => "0010010110101000000100",
			2133 => "0000000010001101000001",
			2134 => "0000011100110100000100",
			2135 => "0000001010001101000001",
			2136 => "0000001010001101000001",
			2137 => "0000000010001101000001",
			2138 => "0010011011101000111100",
			2139 => "0000110011011100011100",
			2140 => "0010011001111000001100",
			2141 => "0001110000101000001000",
			2142 => "0000111000111000000100",
			2143 => "0000000010001101000001",
			2144 => "0000000010001101000001",
			2145 => "1111111010001101000001",
			2146 => "0000011110100000001000",
			2147 => "0011110110110100000100",
			2148 => "0000000010001101000001",
			2149 => "1111111010001101000001",
			2150 => "0011011100101100000100",
			2151 => "0000000010001101000001",
			2152 => "1111111010001101000001",
			2153 => "0010010110101000010000",
			2154 => "0010100001010000001000",
			2155 => "0000101001010000000100",
			2156 => "0000000010001101000001",
			2157 => "0000000010001101000001",
			2158 => "0000100010000000000100",
			2159 => "0000000010001101000001",
			2160 => "0000000010001101000001",
			2161 => "0000110110000100001000",
			2162 => "0011110100010000000100",
			2163 => "0000000010001101000001",
			2164 => "1111111010001101000001",
			2165 => "0011111010010100000100",
			2166 => "0000000010001101000001",
			2167 => "0000000010001101000001",
			2168 => "0000010010001100000100",
			2169 => "1111111010001101000001",
			2170 => "0011110000110100001000",
			2171 => "0011101100110000000100",
			2172 => "1111111010001101000001",
			2173 => "0000000010001101000001",
			2174 => "0000101011101100000100",
			2175 => "0000010010001101000001",
			2176 => "0000000010001101000001",
			2177 => "0000001111000101010100",
			2178 => "0001001011110000101100",
			2179 => "0000001101010000011100",
			2180 => "0010000001110000010000",
			2181 => "0010100111110100001000",
			2182 => "0001001011101100000100",
			2183 => "0000000010001101000001",
			2184 => "1111111010001101000001",
			2185 => "0001111000111000000100",
			2186 => "0000001010001101000001",
			2187 => "0000000010001101000001",
			2188 => "0010011011101000000100",
			2189 => "1111110010001101000001",
			2190 => "0011100001101000000100",
			2191 => "0000000010001101000001",
			2192 => "1111111010001101000001",
			2193 => "0001000011000000000100",
			2194 => "1111111010001101000001",
			2195 => "0001010000001100000100",
			2196 => "0000000010001101000001",
			2197 => "0000101001100000000100",
			2198 => "0000001010001101000001",
			2199 => "0000000010001101000001",
			2200 => "0001111000111000010100",
			2201 => "0001011010111100010000",
			2202 => "0000111010111100001000",
			2203 => "0010000001110000000100",
			2204 => "1111111010001101000001",
			2205 => "0000000010001101000001",
			2206 => "0010001100000100000100",
			2207 => "1111111010001101000001",
			2208 => "1111110010001101000001",
			2209 => "0000000010001101000001",
			2210 => "0001011101010100000100",
			2211 => "0000001010001101000001",
			2212 => "0000100010000100001000",
			2213 => "0001001000000100000100",
			2214 => "0000000010001101000001",
			2215 => "1111111010001101000001",
			2216 => "0001110110100100000100",
			2217 => "0000000010001101000001",
			2218 => "1111111010001101000001",
			2219 => "0010001001101000010100",
			2220 => "0001000110001100001100",
			2221 => "0000010010001100001000",
			2222 => "0011111110101100000100",
			2223 => "0000001010001101000001",
			2224 => "0000000010001101000001",
			2225 => "0000001010001101000001",
			2226 => "0000000010111100000100",
			2227 => "1111111010001101000001",
			2228 => "0000001010001101000001",
			2229 => "0010011011101000011100",
			2230 => "0000000011111100001100",
			2231 => "0000101110010000001000",
			2232 => "0011100110000100000100",
			2233 => "1111111010001101000001",
			2234 => "0000000010001101000001",
			2235 => "1111111010001101000001",
			2236 => "0000101001100000001000",
			2237 => "0011111101000100000100",
			2238 => "0000000010001101000001",
			2239 => "0000001010001101000001",
			2240 => "0010000111000100000100",
			2241 => "0000000010001101000001",
			2242 => "0000000010001101000001",
			2243 => "0000111000000000010000",
			2244 => "0000000011111100001000",
			2245 => "0011111110101100000100",
			2246 => "0000001010001101000001",
			2247 => "0000000010001101000001",
			2248 => "0001001111100000000100",
			2249 => "1111111010001101000001",
			2250 => "0000001010001101000001",
			2251 => "0011111001100000001000",
			2252 => "0011010100000100000100",
			2253 => "0000000010001101000001",
			2254 => "0000010010001101000001",
			2255 => "1111111010001101000001",
			2256 => "0001010011100011000000",
			2257 => "0001000011010101110100",
			2258 => "0011100100010100110100",
			2259 => "0000111001110000010100",
			2260 => "0000000100010100010000",
			2261 => "0001101101111100001000",
			2262 => "0010110100010100000100",
			2263 => "0000001010010101010101",
			2264 => "0000000010010101010101",
			2265 => "0000001010000000000100",
			2266 => "0000010010010101010101",
			2267 => "0000001010010101010101",
			2268 => "1111111010010101010101",
			2269 => "0010010110101000010000",
			2270 => "0001101101111100001000",
			2271 => "0000101100100100000100",
			2272 => "0000010010010101010101",
			2273 => "0000000010010101010101",
			2274 => "0011110010001000000100",
			2275 => "0000011010010101010101",
			2276 => "0000001010010101010101",
			2277 => "0000000000111000001000",
			2278 => "0010000001110000000100",
			2279 => "0000000010010101010101",
			2280 => "0000001010010101010101",
			2281 => "0000111100110000000100",
			2282 => "0000000010010101010101",
			2283 => "0000001010010101010101",
			2284 => "0001100111101000100000",
			2285 => "0010000001010100010000",
			2286 => "0010100011101000001000",
			2287 => "0011000100010100000100",
			2288 => "0000000010010101010101",
			2289 => "1111111010010101010101",
			2290 => "0001001111101000000100",
			2291 => "0000010010010101010101",
			2292 => "1111111010010101010101",
			2293 => "0010010110101000001000",
			2294 => "0001001100001100000100",
			2295 => "0000011010010101010101",
			2296 => "1111111010010101010101",
			2297 => "0011000100010100000100",
			2298 => "1111111010010101010101",
			2299 => "0000000010010101010101",
			2300 => "0000100101110000010000",
			2301 => "0011100100000000001000",
			2302 => "0010010111100100000100",
			2303 => "0000010010010101010101",
			2304 => "0000001010010101010101",
			2305 => "0001101010011000000100",
			2306 => "0000010010010101010101",
			2307 => "0000000010010101010101",
			2308 => "0011101101100000001000",
			2309 => "0011000100010100000100",
			2310 => "0000001010010101010101",
			2311 => "0000000010010101010101",
			2312 => "0010110011011100000100",
			2313 => "0000010010010101010101",
			2314 => "0000001010010101010101",
			2315 => "0001101101111100010000",
			2316 => "0001000011110100000100",
			2317 => "0000001010010101010101",
			2318 => "0000010000011000000100",
			2319 => "1111111010010101010101",
			2320 => "0010000001110100000100",
			2321 => "1111111010010101010101",
			2322 => "0000000010010101010101",
			2323 => "0010111100001000100000",
			2324 => "0000100101001000010000",
			2325 => "0010110100010100001000",
			2326 => "0000111110111100000100",
			2327 => "0000000010010101010101",
			2328 => "0000010010010101010101",
			2329 => "0000110100010100000100",
			2330 => "1111111010010101010101",
			2331 => "0000000010010101010101",
			2332 => "0010010010001100001000",
			2333 => "0001100100110100000100",
			2334 => "0000011010010101010101",
			2335 => "0000000010010101010101",
			2336 => "0011000000101000000100",
			2337 => "0000001010010101010101",
			2338 => "0000011010010101010101",
			2339 => "0011111001010000010000",
			2340 => "0000101001011100001000",
			2341 => "0000000000101000000100",
			2342 => "0000001010010101010101",
			2343 => "1111111010010101010101",
			2344 => "0010100110011100000100",
			2345 => "1111111010010101010101",
			2346 => "0000000010010101010101",
			2347 => "0010110110000100001000",
			2348 => "0000110001101000000100",
			2349 => "0000000010010101010101",
			2350 => "0000011010010101010101",
			2351 => "1111111010010101010101",
			2352 => "0011000110000100110100",
			2353 => "0000111000011000000100",
			2354 => "1111111010010101010101",
			2355 => "0001101101011000010100",
			2356 => "0001100001111000000100",
			2357 => "1111111010010101010101",
			2358 => "0001011000000000001000",
			2359 => "0001101101011000000100",
			2360 => "0000001010010101010101",
			2361 => "0000000010010101010101",
			2362 => "0010111010111000000100",
			2363 => "0000010010010101010101",
			2364 => "0000011010010101010101",
			2365 => "0001101001100100010000",
			2366 => "0000101100010000001000",
			2367 => "0010010001000100000100",
			2368 => "1111111010010101010101",
			2369 => "0000000010010101010101",
			2370 => "0000101000001100000100",
			2371 => "0000001010010101010101",
			2372 => "1111111010010101010101",
			2373 => "0011001100001000000100",
			2374 => "0000000010010101010101",
			2375 => "0001101111000000000100",
			2376 => "1111111010010101010101",
			2377 => "1111111010010101010101",
			2378 => "0011000110000100010100",
			2379 => "0010001111001000010000",
			2380 => "0010000110001000001100",
			2381 => "0010000110011100000100",
			2382 => "1111111010010101010101",
			2383 => "0010001100000100000100",
			2384 => "0000000010010101010101",
			2385 => "1111111010010101010101",
			2386 => "0000001010010101010101",
			2387 => "1111111010010101010101",
			2388 => "1111111010010101010101",
			2389 => "0010010110101010000000",
			2390 => "0000011100110101110000",
			2391 => "0001011100101101000000",
			2392 => "0010110000101000100000",
			2393 => "0010000111000000010000",
			2394 => "0001001011100000001000",
			2395 => "0000001011000100000100",
			2396 => "0000000010011101011001",
			2397 => "0000000010011101011001",
			2398 => "0011110110100100000100",
			2399 => "1111111010011101011001",
			2400 => "0000001010011101011001",
			2401 => "0011110111010000001000",
			2402 => "0000101111010000000100",
			2403 => "0000000010011101011001",
			2404 => "0000001010011101011001",
			2405 => "0000010000011000000100",
			2406 => "0000000010011101011001",
			2407 => "1111111010011101011001",
			2408 => "0011101010000000010000",
			2409 => "0010011001111000001000",
			2410 => "0010101010110000000100",
			2411 => "0000000010011101011001",
			2412 => "0000001010011101011001",
			2413 => "0001110100010100000100",
			2414 => "0000000010011101011001",
			2415 => "1111111010011101011001",
			2416 => "0000101110010000001000",
			2417 => "0001100100110100000100",
			2418 => "0000001010011101011001",
			2419 => "0000001010011101011001",
			2420 => "0001100100110100000100",
			2421 => "1111111010011101011001",
			2422 => "0000000010011101011001",
			2423 => "0001100100110100010100",
			2424 => "0011011100101100000100",
			2425 => "0000000010011101011001",
			2426 => "0001111100001000001000",
			2427 => "0001000101000000000100",
			2428 => "0000000010011101011001",
			2429 => "1111111010011101011001",
			2430 => "0001000101010100000100",
			2431 => "0000000010011101011001",
			2432 => "1111111010011101011001",
			2433 => "0000100101110000001100",
			2434 => "0000100001000000000100",
			2435 => "0000000010011101011001",
			2436 => "0010001110001100000100",
			2437 => "0000001010011101011001",
			2438 => "0000000010011101011001",
			2439 => "0000100010000100001000",
			2440 => "0000101110010000000100",
			2441 => "0000000010011101011001",
			2442 => "1111111010011101011001",
			2443 => "0010100010101000000100",
			2444 => "0000010010011101011001",
			2445 => "0000000010011101011001",
			2446 => "0001010101101100000100",
			2447 => "0000000010011101011001",
			2448 => "0000100101110000001000",
			2449 => "0010111100001000000100",
			2450 => "0000001010011101011001",
			2451 => "0000000010011101011001",
			2452 => "0000010010011101011001",
			2453 => "0000011110100000001100",
			2454 => "0010111100001000001000",
			2455 => "0001110100010100000100",
			2456 => "0000000010011101011001",
			2457 => "1111111010011101011001",
			2458 => "1111110010011101011001",
			2459 => "0011100100010100111100",
			2460 => "0010110000101000011100",
			2461 => "0001000101010100010000",
			2462 => "0001000010110000001000",
			2463 => "0001111011000100000100",
			2464 => "0000000010011101011001",
			2465 => "1111111010011101011001",
			2466 => "0000011110100000000100",
			2467 => "0000001010011101011001",
			2468 => "0000010010011101011001",
			2469 => "0001000011010100001000",
			2470 => "0011110010001000000100",
			2471 => "1111111010011101011001",
			2472 => "0000000010011101011001",
			2473 => "0000000010011101011001",
			2474 => "0011110001011000010000",
			2475 => "0001000100001100001000",
			2476 => "0011100111111000000100",
			2477 => "1111111010011101011001",
			2478 => "0000000010011101011001",
			2479 => "0010100110011100000100",
			2480 => "0000010010011101011001",
			2481 => "1111111010011101011001",
			2482 => "0000101110000100001000",
			2483 => "0011110101100100000100",
			2484 => "1111111010011101011001",
			2485 => "1111111010011101011001",
			2486 => "0001001001001100000100",
			2487 => "0000000010011101011001",
			2488 => "1111111010011101011001",
			2489 => "0000101110000100011100",
			2490 => "0001100001111000010000",
			2491 => "0011100100000000001000",
			2492 => "0001000010010100000100",
			2493 => "0000000010011101011001",
			2494 => "1111111010011101011001",
			2495 => "0010100011101000000100",
			2496 => "1111111010011101011001",
			2497 => "0000001010011101011001",
			2498 => "0001000010111000001000",
			2499 => "0000000011010000000100",
			2500 => "0000000010011101011001",
			2501 => "1111111010011101011001",
			2502 => "0000001010011101011001",
			2503 => "0010000001110100010000",
			2504 => "0010010110101000001000",
			2505 => "0011110101110100000100",
			2506 => "0000001010011101011001",
			2507 => "0000000010011101011001",
			2508 => "0011101000111000000100",
			2509 => "0000000010011101011001",
			2510 => "0000000010011101011001",
			2511 => "0000000111111000001000",
			2512 => "0001101011001100000100",
			2513 => "0000010010011101011001",
			2514 => "0000000010011101011001",
			2515 => "0000011001111000000100",
			2516 => "0000000010011101011001",
			2517 => "1111111010011101011001",
			2518 => "0011000100001010101100",
			2519 => "0000111011000100111000",
			2520 => "0011110001011000110100",
			2521 => "0001110111111000011000",
			2522 => "0010001001101000001000",
			2523 => "0000111010000000000100",
			2524 => "0000001010100010110101",
			2525 => "0000010010100010110101",
			2526 => "0001110111111000001000",
			2527 => "0011000111111000000100",
			2528 => "0000000010100010110101",
			2529 => "0000001010100010110101",
			2530 => "0011000111111000000100",
			2531 => "0000001010100010110101",
			2532 => "1111111010100010110101",
			2533 => "0000110111111000010000",
			2534 => "0010100110011100001000",
			2535 => "0001100001111000000100",
			2536 => "0000000010100010110101",
			2537 => "1111111010100010110101",
			2538 => "0010100001110000000100",
			2539 => "0000000010100010110101",
			2540 => "1111111010100010110101",
			2541 => "0010111110111100000100",
			2542 => "0000001010100010110101",
			2543 => "0001000000010100000100",
			2544 => "0000000010100010110101",
			2545 => "0000000010100010110101",
			2546 => "1111111010100010110101",
			2547 => "0011110010001000111100",
			2548 => "0001010011011100011100",
			2549 => "0010101010110000010000",
			2550 => "0011011100110000001000",
			2551 => "0010111011000100000100",
			2552 => "0000000010100010110101",
			2553 => "1111111010100010110101",
			2554 => "0000110100000000000100",
			2555 => "0000001010100010110101",
			2556 => "0000010010100010110101",
			2557 => "0001010011011100001000",
			2558 => "0011000111111000000100",
			2559 => "0000010010100010110101",
			2560 => "0000000010100010110101",
			2561 => "0000010010100010110101",
			2562 => "0000110100000000010000",
			2563 => "0011110110100100001000",
			2564 => "0011011100101100000100",
			2565 => "0000010010100010110101",
			2566 => "0000000010100010110101",
			2567 => "0000011110100000000100",
			2568 => "0000000010100010110101",
			2569 => "0000001010100010110101",
			2570 => "0011011100101000001000",
			2571 => "0000111100110000000100",
			2572 => "0000000010100010110101",
			2573 => "0000000010100010110101",
			2574 => "0000111110001100000100",
			2575 => "1111111010100010110101",
			2576 => "0000000010100010110101",
			2577 => "0000110101101100011000",
			2578 => "0000110101101100010000",
			2579 => "0000111100110000001000",
			2580 => "0011010110000100000100",
			2581 => "0000000010100010110101",
			2582 => "1111111010100010110101",
			2583 => "0011000100010100000100",
			2584 => "0000001010100010110101",
			2585 => "0000000010100010110101",
			2586 => "0011110101110100000100",
			2587 => "1111111010100010110101",
			2588 => "1111111010100010110101",
			2589 => "0010000010101000010000",
			2590 => "0001000000010100001000",
			2591 => "0010000111000100000100",
			2592 => "0000000010100010110101",
			2593 => "0000000010100010110101",
			2594 => "0010101010110000000100",
			2595 => "0000000010100010110101",
			2596 => "0000000010100010110101",
			2597 => "0000100010000000001000",
			2598 => "0001101010011000000100",
			2599 => "0000010010100010110101",
			2600 => "0000000010100010110101",
			2601 => "0001000010100100000100",
			2602 => "0000001010100010110101",
			2603 => "0000000010100010110101",
			2604 => "1111111010100010110101",
			2605 => "0011110000110111100100",
			2606 => "0011101010000001101100",
			2607 => "0010110100010100110100",
			2608 => "0000011110100000011100",
			2609 => "0010011001111000010000",
			2610 => "0011000111111000001000",
			2611 => "0001110111111000000100",
			2612 => "0000000010101110100011",
			2613 => "0000000010101110100011",
			2614 => "0001111010000000000100",
			2615 => "1111111010101110100011",
			2616 => "0000000010101110100011",
			2617 => "0010110100010100001000",
			2618 => "0011000111111000000100",
			2619 => "0000000010101110100011",
			2620 => "1111111010101110100011",
			2621 => "0000000010101110100011",
			2622 => "0011000111111000001100",
			2623 => "0010011001111000000100",
			2624 => "0000001010101110100011",
			2625 => "0000111100001000000100",
			2626 => "1111111010101110100011",
			2627 => "0000000010101110100011",
			2628 => "0001111011000100001000",
			2629 => "0011010101101100000100",
			2630 => "0000001010101110100011",
			2631 => "0000000010101110100011",
			2632 => "0000000010101110100011",
			2633 => "0001101100011000011000",
			2634 => "0000100010000000010000",
			2635 => "0010010010001100001000",
			2636 => "0000010110000000000100",
			2637 => "0000000010101110100011",
			2638 => "0000010010101110100011",
			2639 => "0011100000111000000100",
			2640 => "1111111010101110100011",
			2641 => "0000000010101110100011",
			2642 => "0000100010000000000100",
			2643 => "0000100010101110100011",
			2644 => "0000000010101110100011",
			2645 => "0011110100000100010000",
			2646 => "0011111000011000001000",
			2647 => "0000101111010000000100",
			2648 => "1111111010101110100011",
			2649 => "0000001010101110100011",
			2650 => "0001111100001000000100",
			2651 => "0000001010101110100011",
			2652 => "1111111010101110100011",
			2653 => "0011011110001100001000",
			2654 => "0001011101100000000100",
			2655 => "0000000010101110100011",
			2656 => "1111111010101110100011",
			2657 => "0010010110101000000100",
			2658 => "0000001010101110100011",
			2659 => "1111111010101110100011",
			2660 => "0011011100101100111100",
			2661 => "0010110000101000100000",
			2662 => "0000110101101100010000",
			2663 => "0011110101110100001000",
			2664 => "0011000100010100000100",
			2665 => "0000000010101110100011",
			2666 => "0000001010101110100011",
			2667 => "0001110100010100000100",
			2668 => "0000000010101110100011",
			2669 => "1111111010101110100011",
			2670 => "0001001010110100001000",
			2671 => "0011111010010100000100",
			2672 => "0000000010101110100011",
			2673 => "1111111010101110100011",
			2674 => "0001000000010100000100",
			2675 => "0000010010101110100011",
			2676 => "0000001010101110100011",
			2677 => "0010100001010000010000",
			2678 => "0010100110011000001000",
			2679 => "0001110100010100000100",
			2680 => "0000001010101110100011",
			2681 => "0000000010101110100011",
			2682 => "0000100100101000000100",
			2683 => "0000000010101110100011",
			2684 => "0000001010101110100011",
			2685 => "0011111011011100000100",
			2686 => "0000010010101110100011",
			2687 => "0011100100010100000100",
			2688 => "0000000010101110100011",
			2689 => "0000001010101110100011",
			2690 => "0011101101100000100000",
			2691 => "0010010111100100010000",
			2692 => "0000011100110100001000",
			2693 => "0010010110101000000100",
			2694 => "0000000010101110100011",
			2695 => "0000000010101110100011",
			2696 => "0011000100000000000100",
			2697 => "0000000010101110100011",
			2698 => "0000001010101110100011",
			2699 => "0001000011001100001000",
			2700 => "0000111110001100000100",
			2701 => "1111111010101110100011",
			2702 => "0000000010101110100011",
			2703 => "0001101010011000000100",
			2704 => "1111111010101110100011",
			2705 => "0000000010101110100011",
			2706 => "0010011011101000010000",
			2707 => "0011000100010100001000",
			2708 => "0011000100010100000100",
			2709 => "0000000010101110100011",
			2710 => "1111111010101110100011",
			2711 => "0010110100000000000100",
			2712 => "0000001010101110100011",
			2713 => "0000000010101110100011",
			2714 => "0010101010110000001000",
			2715 => "0000011001111000000100",
			2716 => "0000000010101110100011",
			2717 => "0000000010101110100011",
			2718 => "1111111010101110100011",
			2719 => "0001110100000001011100",
			2720 => "0010101100011100101100",
			2721 => "0001001010110100011000",
			2722 => "0011000100000000001100",
			2723 => "0001101101111100000100",
			2724 => "1111111010101110100011",
			2725 => "0000100010000000000100",
			2726 => "0000000010101110100011",
			2727 => "0000000010101110100011",
			2728 => "0011011010111000001000",
			2729 => "0010100001010000000100",
			2730 => "1111111010101110100011",
			2731 => "0000000010101110100011",
			2732 => "0000000010101110100011",
			2733 => "0011010101101100001000",
			2734 => "0001110111111000000100",
			2735 => "1111111010101110100011",
			2736 => "0000001010101110100011",
			2737 => "0000100011001000000100",
			2738 => "0000000010101110100011",
			2739 => "0011000100000000000100",
			2740 => "1111111010101110100011",
			2741 => "0000000010101110100011",
			2742 => "0010111001110000100000",
			2743 => "0001000011010100010000",
			2744 => "0001010000001100001000",
			2745 => "0000100110010000000100",
			2746 => "0000001010101110100011",
			2747 => "0000000010101110100011",
			2748 => "0001101010011000000100",
			2749 => "0000010010101110100011",
			2750 => "0000001010101110100011",
			2751 => "0001111100001000001000",
			2752 => "0011101000111000000100",
			2753 => "1111111010101110100011",
			2754 => "0000000010101110100011",
			2755 => "0011000100010100000100",
			2756 => "0000000010101110100011",
			2757 => "1111111010101110100011",
			2758 => "0011000000101000000100",
			2759 => "0000001010101110100011",
			2760 => "0011101100101100000100",
			2761 => "0000000010101110100011",
			2762 => "0001011010111100000100",
			2763 => "1111111010101110100011",
			2764 => "1111111010101110100011",
			2765 => "0001111000111000011100",
			2766 => "0011110000110100000100",
			2767 => "1111111010101110100011",
			2768 => "0000010010001100001100",
			2769 => "0010111000111000000100",
			2770 => "0000000010101110100011",
			2771 => "0000010010001100000100",
			2772 => "0000001010101110100011",
			2773 => "0000001010101110100011",
			2774 => "0001101101011000001000",
			2775 => "0001000011110000000100",
			2776 => "0000001010101110100011",
			2777 => "0000000010101110100011",
			2778 => "0000001010101110100011",
			2779 => "0000110100001000000100",
			2780 => "0000001010101110100011",
			2781 => "0010010111100100001000",
			2782 => "0011111110101100000100",
			2783 => "1111111010101110100011",
			2784 => "1111110010101110100011",
			2785 => "0011000000101000001000",
			2786 => "0001101010011000000100",
			2787 => "0000000010101110100011",
			2788 => "1111111010101110100011",
			2789 => "0000100101110000000100",
			2790 => "1111111010101110100011",
			2791 => "0000000010101110100011",
			2792 => "0001011000000001110100",
			2793 => "0001111101100001011000",
			2794 => "0001111101100000111100",
			2795 => "0001110000101000100000",
			2796 => "0001110100010100010000",
			2797 => "0001110100010100001000",
			2798 => "0000011100110100000100",
			2799 => "0000000010110100010101",
			2800 => "0000001010110100010101",
			2801 => "0010110100010100000100",
			2802 => "1111111010110100010101",
			2803 => "0000000010110100010101",
			2804 => "0001010011011100001000",
			2805 => "0001111011000100000100",
			2806 => "0000001010110100010101",
			2807 => "0000000010110100010101",
			2808 => "0000100010000100000100",
			2809 => "0000000010110100010101",
			2810 => "0000001010110100010101",
			2811 => "0001110000101000001100",
			2812 => "0001100111101000000100",
			2813 => "0000001010110100010101",
			2814 => "0001011110001100000100",
			2815 => "1111111010110100010101",
			2816 => "0000000010110100010101",
			2817 => "0010100111110100001000",
			2818 => "0000101001010000000100",
			2819 => "0000000010110100010101",
			2820 => "1111111010110100010101",
			2821 => "0001111100001000000100",
			2822 => "0000000010110100010101",
			2823 => "0000000010110100010101",
			2824 => "0011101010111000001100",
			2825 => "0001111101100000001000",
			2826 => "0010000110001000000100",
			2827 => "0000001010110100010101",
			2828 => "0000010010110100010101",
			2829 => "0000000010110100010101",
			2830 => "0001101101011000000100",
			2831 => "1111111010110100010101",
			2832 => "0011001000111100001000",
			2833 => "0010111100101100000100",
			2834 => "1111111010110100010101",
			2835 => "0000000010110100010101",
			2836 => "0000001010110100010101",
			2837 => "0010100110011000010000",
			2838 => "0011001000111000000100",
			2839 => "1111111010110100010101",
			2840 => "0011001001110000001000",
			2841 => "0010101100011000000100",
			2842 => "0000000010110100010101",
			2843 => "0000001010110100010101",
			2844 => "1111111010110100010101",
			2845 => "0011111001010000000100",
			2846 => "1111111010110100010101",
			2847 => "0000110000011100000100",
			2848 => "0000000010110100010101",
			2849 => "1111111010110100010101",
			2850 => "0011101001010100101100",
			2851 => "0010101100011100101000",
			2852 => "0010001111001000011000",
			2853 => "0001011000011000001100",
			2854 => "0000101100010000001000",
			2855 => "0010100001010000000100",
			2856 => "0000001010110100010101",
			2857 => "1111111010110100010101",
			2858 => "1111111010110100010101",
			2859 => "0001011010001100001000",
			2860 => "0000101100100100000100",
			2861 => "0000000010110100010101",
			2862 => "0000001010110100010101",
			2863 => "0000000010110100010101",
			2864 => "0000100111011000000100",
			2865 => "0000001010110100010101",
			2866 => "0011110010000000001000",
			2867 => "0001111110001100000100",
			2868 => "0000010010110100010101",
			2869 => "0000000010110100010101",
			2870 => "0000000010110100010101",
			2871 => "1111111010110100010101",
			2872 => "0000011101101000001000",
			2873 => "0000100110010000000100",
			2874 => "0000000010110100010101",
			2875 => "1111111010110100010101",
			2876 => "0011001010111100010000",
			2877 => "0001101111000000001100",
			2878 => "0000100010000100000100",
			2879 => "0000000010110100010101",
			2880 => "0011001100110000000100",
			2881 => "0000001010110100010101",
			2882 => "0000000010110100010101",
			2883 => "1111111010110100010101",
			2884 => "1111111010110100010101",
			2885 => "0001111101100001111000",
			2886 => "0000011100100000001000",
			2887 => "0001101101111100000100",
			2888 => "1111111010111001111001",
			2889 => "0000001010111001111001",
			2890 => "0010000111000101000000",
			2891 => "0001101101111100100000",
			2892 => "0000101010001000010000",
			2893 => "0000110100000000001000",
			2894 => "0010110111111000000100",
			2895 => "0000001010111001111001",
			2896 => "0000000010111001111001",
			2897 => "0010100111110100000100",
			2898 => "0000000010111001111001",
			2899 => "0000001010111001111001",
			2900 => "0010000110001000001000",
			2901 => "0000111110001100000100",
			2902 => "1111111010111001111001",
			2903 => "0000000010111001111001",
			2904 => "0001110100010100000100",
			2905 => "0000001010111001111001",
			2906 => "1111111010111001111001",
			2907 => "0000101001100000010000",
			2908 => "0010001111001000001000",
			2909 => "0011000100000000000100",
			2910 => "0000001010111001111001",
			2911 => "0000001010111001111001",
			2912 => "0010100001010000000100",
			2913 => "0000000010111001111001",
			2914 => "0000001010111001111001",
			2915 => "0011100001111100001000",
			2916 => "0000101110110100000100",
			2917 => "0000000010111001111001",
			2918 => "1111111010111001111001",
			2919 => "0001011010111000000100",
			2920 => "0000001010111001111001",
			2921 => "0000000010111001111001",
			2922 => "0001110111111000010100",
			2923 => "0000101101000100001000",
			2924 => "0010111110111100000100",
			2925 => "0000001010111001111001",
			2926 => "0000000010111001111001",
			2927 => "0000011110100000001000",
			2928 => "0010000010101000000100",
			2929 => "0000001010111001111001",
			2930 => "0000010010111001111001",
			2931 => "0000000010111001111001",
			2932 => "0010000111000000010000",
			2933 => "0000110100010100001000",
			2934 => "0001101100011000000100",
			2935 => "1111111010111001111001",
			2936 => "0000001010111001111001",
			2937 => "0001111100001000000100",
			2938 => "0000001010111001111001",
			2939 => "0000000010111001111001",
			2940 => "0001100100110100000100",
			2941 => "0000001010111001111001",
			2942 => "0000011110100000000100",
			2943 => "0000000010111001111001",
			2944 => "1111111010111001111001",
			2945 => "0011001100110000101100",
			2946 => "0000110001101000010000",
			2947 => "0000111001110100000100",
			2948 => "1111111010111001111001",
			2949 => "0000100011001000001000",
			2950 => "0001011001110100000100",
			2951 => "0000001010111001111001",
			2952 => "1111111010111001111001",
			2953 => "1111111010111001111001",
			2954 => "0001101011001100010000",
			2955 => "0001100001111000000100",
			2956 => "1111111010111001111001",
			2957 => "0011111110101000000100",
			2958 => "0000010010111001111001",
			2959 => "0000101100010000000100",
			2960 => "0000000010111001111001",
			2961 => "0000001010111001111001",
			2962 => "0011010111010000000100",
			2963 => "1111111010111001111001",
			2964 => "0000100000010000000100",
			2965 => "0000011010111001111001",
			2966 => "1111111010111001111001",
			2967 => "0001111101111000001100",
			2968 => "0001111110001100000100",
			2969 => "1111111010111001111001",
			2970 => "0011000110000100000100",
			2971 => "0000001010111001111001",
			2972 => "1111111010111001111001",
			2973 => "1111111010111001111001",
			2974 => "0011000011011101101100",
			2975 => "0001000011111001101000",
			2976 => "0001111001110001000000",
			2977 => "0011101101100000100000",
			2978 => "0010011101101000010000",
			2979 => "0000101010001000001000",
			2980 => "0011100100010100000100",
			2981 => "0000000010111110100101",
			2982 => "0000000010111110100101",
			2983 => "0010100001010000000100",
			2984 => "0000000010111110100101",
			2985 => "0000000010111110100101",
			2986 => "0001000011001100001000",
			2987 => "0000111110001100000100",
			2988 => "1111111010111110100101",
			2989 => "0000000010111110100101",
			2990 => "0010000110001000000100",
			2991 => "1111111010111110100101",
			2992 => "0000000010111110100101",
			2993 => "0010011101101000010000",
			2994 => "0001001111100000001000",
			2995 => "0010100110011100000100",
			2996 => "0000001010111110100101",
			2997 => "0000010010111110100101",
			2998 => "0011101110001100000100",
			2999 => "1111111010111110100101",
			3000 => "0000000010111110100101",
			3001 => "0011100110000100001000",
			3002 => "0000100111111100000100",
			3003 => "0000000010111110100101",
			3004 => "1111111010111110100101",
			3005 => "0001001101001000000100",
			3006 => "0000001010111110100101",
			3007 => "0000000010111110100101",
			3008 => "0001101111000000100000",
			3009 => "0000100111011000010000",
			3010 => "0010101100011100001000",
			3011 => "0001100001111000000100",
			3012 => "1111111010111110100101",
			3013 => "0000000010111110100101",
			3014 => "0010011011101000000100",
			3015 => "0000000010111110100101",
			3016 => "1111111010111110100101",
			3017 => "0000001010000000001000",
			3018 => "0001111101100000000100",
			3019 => "1111111010111110100101",
			3020 => "0000001010111110100101",
			3021 => "0010110110000100000100",
			3022 => "0000010010111110100101",
			3023 => "0000000010111110100101",
			3024 => "0010110001111100000100",
			3025 => "1111111010111110100101",
			3026 => "0000000010111110100101",
			3027 => "1111111010111110100101",
			3028 => "0011000110000100011000",
			3029 => "0010111000000000010100",
			3030 => "0010011101011100000100",
			3031 => "1111111010111110100101",
			3032 => "0010011101011100000100",
			3033 => "0000001010111110100101",
			3034 => "0010111010111100001000",
			3035 => "0011010111010000000100",
			3036 => "1111111010111110100101",
			3037 => "0000001010111110100101",
			3038 => "1111111010111110100101",
			3039 => "0000001010111110100101",
			3040 => "0011001010111100010000",
			3041 => "0010000110011100001100",
			3042 => "0010001100011100000100",
			3043 => "1111111010111110100101",
			3044 => "0011000100001000000100",
			3045 => "0000000010111110100101",
			3046 => "0000010010111110100101",
			3047 => "1111111010111110100101",
			3048 => "1111111010111110100101",
			3049 => "0011000011011101111000",
			3050 => "0001000011111001110100",
			3051 => "0010011111001100111100",
			3052 => "0001101010011000100000",
			3053 => "0011110010110100010000",
			3054 => "0011100110000100001000",
			3055 => "0010011101101000000100",
			3056 => "0000000011000100000001",
			3057 => "0000000011000100000001",
			3058 => "0010110011011100000100",
			3059 => "0000001011000100000001",
			3060 => "0000000011000100000001",
			3061 => "0001101100011000001000",
			3062 => "0011111110101000000100",
			3063 => "0000000011000100000001",
			3064 => "1111111011000100000001",
			3065 => "0001001101001000000100",
			3066 => "0000001011000100000001",
			3067 => "0000000011000100000001",
			3068 => "0000001011000100010000",
			3069 => "0010011101101000001000",
			3070 => "0001001111100000000100",
			3071 => "0000001011000100000001",
			3072 => "0000000011000100000001",
			3073 => "0000110100011000000100",
			3074 => "0000000011000100000001",
			3075 => "0000001011000100000001",
			3076 => "0001101010011000000100",
			3077 => "0000010011000100000001",
			3078 => "0011100000001100000100",
			3079 => "1111111011000100000001",
			3080 => "0000001011000100000001",
			3081 => "0011100111001000011100",
			3082 => "0000000011010000010000",
			3083 => "0011111010010100001000",
			3084 => "0010110110000100000100",
			3085 => "1111110011000100000001",
			3086 => "1111111011000100000001",
			3087 => "0010111100110000000100",
			3088 => "0000000011000100000001",
			3089 => "0000001011000100000001",
			3090 => "0000111001110100001000",
			3091 => "0001111101100000000100",
			3092 => "1111111011000100000001",
			3093 => "1111111011000100000001",
			3094 => "0000000011000100000001",
			3095 => "0011000000101000001100",
			3096 => "0001001000000100000100",
			3097 => "0000000011000100000001",
			3098 => "0010111101100000000100",
			3099 => "1111110011000100000001",
			3100 => "1111111011000100000001",
			3101 => "0001111000111000001000",
			3102 => "0010011001011000000100",
			3103 => "0000001011000100000001",
			3104 => "0000000011000100000001",
			3105 => "0001001000100000000100",
			3106 => "0000001011000100000001",
			3107 => "0000000011000100000001",
			3108 => "1111111011000100000001",
			3109 => "0011000110000100100100",
			3110 => "0010011011111100010000",
			3111 => "0001110101101100000100",
			3112 => "1111111011000100000001",
			3113 => "0001110101101100000100",
			3114 => "0000001011000100000001",
			3115 => "0010111100101100000100",
			3116 => "0000000011000100000001",
			3117 => "1111111011000100000001",
			3118 => "0000000010101000001000",
			3119 => "0011111100100100000100",
			3120 => "1111111011000100000001",
			3121 => "0000001011000100000001",
			3122 => "0010010111101000001000",
			3123 => "0010011110010100000100",
			3124 => "0000000011000100000001",
			3125 => "0000001011000100000001",
			3126 => "1111111011000100000001",
			3127 => "0011001010111100010000",
			3128 => "0010000110011100001100",
			3129 => "0010001100011100000100",
			3130 => "1111111011000100000001",
			3131 => "0011000100001000000100",
			3132 => "0000000011000100000001",
			3133 => "0000001011000100000001",
			3134 => "1111111011000100000001",
			3135 => "1111111011000100000001",
			3136 => "0011001000111001111000",
			3137 => "0010010110000000000100",
			3138 => "1111111011001001100101",
			3139 => "0011101100001000111000",
			3140 => "0001111100001000011100",
			3141 => "0011100011010000001100",
			3142 => "0010000101000100000100",
			3143 => "0000010011001001100101",
			3144 => "0010011100110100000100",
			3145 => "0000001011001001100101",
			3146 => "0000000011001001100101",
			3147 => "0011110010001000001000",
			3148 => "0010000101000100000100",
			3149 => "1111111011001001100101",
			3150 => "0000001011001001100101",
			3151 => "0011011100101100000100",
			3152 => "0000000011001001100101",
			3153 => "0000000011001001100101",
			3154 => "0000111101100000010000",
			3155 => "0010010110101000001000",
			3156 => "0000111100001000000100",
			3157 => "1111111011001001100101",
			3158 => "0000000011001001100101",
			3159 => "0010101000010100000100",
			3160 => "0000000011001001100101",
			3161 => "1111111011001001100101",
			3162 => "0010010110101000000100",
			3163 => "0000010011001001100101",
			3164 => "0011110000011100000100",
			3165 => "0000001011001001100101",
			3166 => "0000000011001001100101",
			3167 => "0000101010001000100000",
			3168 => "0001100001111000010000",
			3169 => "0010110100000000001000",
			3170 => "0011011110001100000100",
			3171 => "0000000011001001100101",
			3172 => "0000001011001001100101",
			3173 => "0001100111101000000100",
			3174 => "1111111011001001100101",
			3175 => "0000000011001001100101",
			3176 => "0010011101101000001000",
			3177 => "0011110010001000000100",
			3178 => "0000010011001001100101",
			3179 => "0000001011001001100101",
			3180 => "0010000111000100000100",
			3181 => "0000001011001001100101",
			3182 => "1111111011001001100101",
			3183 => "0000110001011000010000",
			3184 => "0011100110000100001000",
			3185 => "0010111100001000000100",
			3186 => "0000001011001001100101",
			3187 => "0000000011001001100101",
			3188 => "0001110100000000000100",
			3189 => "0000001011001001100101",
			3190 => "0000001011001001100101",
			3191 => "0001010001101000001000",
			3192 => "0011011000000000000100",
			3193 => "0000000011001001100101",
			3194 => "1111111011001001100101",
			3195 => "0000001011001001100101",
			3196 => "0011001100110000101100",
			3197 => "0011111101000100010000",
			3198 => "0001111001110000000100",
			3199 => "0000000011001001100101",
			3200 => "0011110010110100000100",
			3201 => "1111111011001001100101",
			3202 => "0011110110100000000100",
			3203 => "0000000011001001100101",
			3204 => "1111111011001001100101",
			3205 => "0000101000001100010100",
			3206 => "0011010100000100001100",
			3207 => "0000010111100100001000",
			3208 => "0011010001101000000100",
			3209 => "0000000011001001100101",
			3210 => "0000001011001001100101",
			3211 => "1111111011001001100101",
			3212 => "0000110110100000000100",
			3213 => "0000010011001001100101",
			3214 => "0000000011001001100101",
			3215 => "0010100001010000000100",
			3216 => "0000000011001001100101",
			3217 => "1111111011001001100101",
			3218 => "0001111101111000001100",
			3219 => "0001111110001100000100",
			3220 => "1111111011001001100101",
			3221 => "0011000110000100000100",
			3222 => "0000001011001001100101",
			3223 => "1111111011001001100101",
			3224 => "1111111011001001100101",
			3225 => "0011000110000101111000",
			3226 => "0001000011111001110100",
			3227 => "0000101110000100111100",
			3228 => "0001100111101000011100",
			3229 => "0001010101101100010000",
			3230 => "0000111000111100001000",
			3231 => "0010000001110000000100",
			3232 => "0000001011001110001001",
			3233 => "0000000011001110001001",
			3234 => "0001110100010100000100",
			3235 => "0000000011001110001001",
			3236 => "0000010011001110001001",
			3237 => "0011111010001100000100",
			3238 => "1111111011001110001001",
			3239 => "0010011011101000000100",
			3240 => "0000000011001110001001",
			3241 => "0000001011001110001001",
			3242 => "0011011100110000010000",
			3243 => "0001001001001100001000",
			3244 => "0010001011010100000100",
			3245 => "0000000011001110001001",
			3246 => "1111111011001110001001",
			3247 => "0010100001010000000100",
			3248 => "0000010011001110001001",
			3249 => "0000000011001110001001",
			3250 => "0010101001000100001000",
			3251 => "0000111101100000000100",
			3252 => "0000000011001110001001",
			3253 => "0000000011001110001001",
			3254 => "0001101101111100000100",
			3255 => "0000001011001110001001",
			3256 => "0000000011001110001001",
			3257 => "0010101100011100011100",
			3258 => "0000101110000100001100",
			3259 => "0001001110100100000100",
			3260 => "1111111011001110001001",
			3261 => "0001000011110000000100",
			3262 => "0000001011001110001001",
			3263 => "1111111011001110001001",
			3264 => "0001001110111000001000",
			3265 => "0010100001010000000100",
			3266 => "0000000011001110001001",
			3267 => "0000000011001110001001",
			3268 => "0000010110000000000100",
			3269 => "0000001011001110001001",
			3270 => "0000000011001110001001",
			3271 => "0011110111010000001100",
			3272 => "0000100101001000000100",
			3273 => "0000000011001110001001",
			3274 => "0000110100010100000100",
			3275 => "0000001011001110001001",
			3276 => "0000010011001110001001",
			3277 => "0010000111000000001000",
			3278 => "0001000011011000000100",
			3279 => "0000000011001110001001",
			3280 => "0000010011001110001001",
			3281 => "0000100100101000000100",
			3282 => "1111111011001110001001",
			3283 => "0000000011001110001001",
			3284 => "1111111011001110001001",
			3285 => "0011001010111100011000",
			3286 => "0000111100111000010000",
			3287 => "0001111101111000001100",
			3288 => "0001101011001100000100",
			3289 => "1111111011001110001001",
			3290 => "0001101001100100000100",
			3291 => "0000001011001110001001",
			3292 => "0000000011001110001001",
			3293 => "1111111011001110001001",
			3294 => "0001000011001100000100",
			3295 => "0000010011001110001001",
			3296 => "0000000011001110001001",
			3297 => "1111111011001110001001",
			3298 => "0001110101101110000000",
			3299 => "0010011110100000001000",
			3300 => "0001101101111100000100",
			3301 => "1111111011010100001101",
			3302 => "0000001011010100001101",
			3303 => "0001001110111001000000",
			3304 => "0001101101111100100000",
			3305 => "0000100101110000010000",
			3306 => "0011111010011100001000",
			3307 => "0010110000101000000100",
			3308 => "0000000011010100001101",
			3309 => "1111111011010100001101",
			3310 => "0000110011011100000100",
			3311 => "0000000011010100001101",
			3312 => "0000001011010100001101",
			3313 => "0000001111000100001000",
			3314 => "0001001011110000000100",
			3315 => "0000000011010100001101",
			3316 => "1111111011010100001101",
			3317 => "0000111101111000000100",
			3318 => "0000000011010100001101",
			3319 => "0000001011010100001101",
			3320 => "0010110101101100010000",
			3321 => "0001000011001100001000",
			3322 => "0010100001010000000100",
			3323 => "0000001011010100001101",
			3324 => "0000001011010100001101",
			3325 => "0010100110011000000100",
			3326 => "0000000011010100001101",
			3327 => "0000001011010100001101",
			3328 => "0001101101011000001000",
			3329 => "0001000010010100000100",
			3330 => "0000010011010100001101",
			3331 => "0000000011010100001101",
			3332 => "0010010101011100000100",
			3333 => "0000000011010100001101",
			3334 => "1111111011010100001101",
			3335 => "0010010110101000011100",
			3336 => "0000100110100000010000",
			3337 => "0001101101111100001000",
			3338 => "0001100001111000000100",
			3339 => "1111111011010100001101",
			3340 => "0000011011010100001101",
			3341 => "0001110100010100000100",
			3342 => "1111111011010100001101",
			3343 => "0000000011010100001101",
			3344 => "0010100110011000000100",
			3345 => "1111111011010100001101",
			3346 => "0011000000110000000100",
			3347 => "0000010011010100001101",
			3348 => "0000001011010100001101",
			3349 => "0011101011000100001100",
			3350 => "0010000010101000001000",
			3351 => "0011110110110100000100",
			3352 => "0000000011010100001101",
			3353 => "1111111011010100001101",
			3354 => "1111111011010100001101",
			3355 => "0001001111100000001000",
			3356 => "0010000001110100000100",
			3357 => "0000000011010100001101",
			3358 => "0000001011010100001101",
			3359 => "0001111011000100000100",
			3360 => "0000001011010100001101",
			3361 => "0000000011010100001101",
			3362 => "0011000110000100101100",
			3363 => "0011010111010000011000",
			3364 => "0011101000000000000100",
			3365 => "1111111011010100001101",
			3366 => "0001000110001100001100",
			3367 => "0011110111100000001000",
			3368 => "0011100110100100000100",
			3369 => "1111111011010100001101",
			3370 => "0000000011010100001101",
			3371 => "1111111011010100001101",
			3372 => "0011000011011100000100",
			3373 => "0000001011010100001101",
			3374 => "1111111011010100001101",
			3375 => "0001001001001100010000",
			3376 => "0001101111000000001000",
			3377 => "0000001001101000000100",
			3378 => "1111111011010100001101",
			3379 => "0000010011010100001101",
			3380 => "0010001111001000000100",
			3381 => "1111111011010100001101",
			3382 => "0000000011010100001101",
			3383 => "1111111011010100001101",
			3384 => "0011001010111100010100",
			3385 => "0001110110100100010000",
			3386 => "0001111101111000001100",
			3387 => "0001111110001100000100",
			3388 => "1111111011010100001101",
			3389 => "0011000110000100000100",
			3390 => "0000000011010100001101",
			3391 => "1111111011010100001101",
			3392 => "1111111011010100001101",
			3393 => "0000100011010100001101",
			3394 => "1111111011010100001101",
			3395 => "0010000111000010011000",
			3396 => "0010100110011101111000",
			3397 => "0010100001010000111100",
			3398 => "0010000110001000100000",
			3399 => "0010010110101000010000",
			3400 => "0001110111111000001000",
			3401 => "0010001011010100000100",
			3402 => "0000000011011011011001",
			3403 => "1111111011011011011001",
			3404 => "0001000101010100000100",
			3405 => "0000000011011011011001",
			3406 => "0000001011011011011001",
			3407 => "0010010110101000001000",
			3408 => "0001100001111000000100",
			3409 => "1111111011011011011001",
			3410 => "0000000011011011011001",
			3411 => "0010010110101000000100",
			3412 => "0000000011011011011001",
			3413 => "0000000011011011011001",
			3414 => "0001001110111000010000",
			3415 => "0010100001010000001000",
			3416 => "0011000111111000000100",
			3417 => "1111111011011011011001",
			3418 => "0000000011011011011001",
			3419 => "0001110100010100000100",
			3420 => "0000000011011011011001",
			3421 => "1111111011011011011001",
			3422 => "0010001111001000000100",
			3423 => "1111111011011011011001",
			3424 => "0001100001111000000100",
			3425 => "1111111011011011011001",
			3426 => "0000001011011011011001",
			3427 => "0001000101010100100000",
			3428 => "0011011010111100010000",
			3429 => "0001101101111100001000",
			3430 => "0010010110101000000100",
			3431 => "0000000011011011011001",
			3432 => "1111111011011011011001",
			3433 => "0011110101110100000100",
			3434 => "0000001011011011011001",
			3435 => "0000000011011011011001",
			3436 => "0011111101000100001000",
			3437 => "0011011101010100000100",
			3438 => "1111111011011011011001",
			3439 => "0000000011011011011001",
			3440 => "0011100001111100000100",
			3441 => "0000001011011011011001",
			3442 => "0000000011011011011001",
			3443 => "0011000111111000001100",
			3444 => "0011110010110100001000",
			3445 => "0011000111111000000100",
			3446 => "0000000011011011011001",
			3447 => "0000000011011011011001",
			3448 => "0000001011011011011001",
			3449 => "0000000000110000001000",
			3450 => "0010010111100100000100",
			3451 => "0000001011011011011001",
			3452 => "1111111011011011011001",
			3453 => "0011011010111100000100",
			3454 => "0000000011011011011001",
			3455 => "0000000011011011011001",
			3456 => "0010010110101000000100",
			3457 => "0000001011011011011001",
			3458 => "0010111000111100001000",
			3459 => "0011100011011100000100",
			3460 => "1111111011011011011001",
			3461 => "0000000011011011011001",
			3462 => "0010011011101000001000",
			3463 => "0011101101100000000100",
			3464 => "0000000011011011011001",
			3465 => "0000001011011011011001",
			3466 => "0011111001010000000100",
			3467 => "1111111011011011011001",
			3468 => "0000011001111000000100",
			3469 => "0000001011011011011001",
			3470 => "1111111011011011011001",
			3471 => "0011000111111000011100",
			3472 => "0000001000111100000100",
			3473 => "1111111011011011011001",
			3474 => "0010110100010100010000",
			3475 => "0010011100110100001100",
			3476 => "0011110100001000000100",
			3477 => "0000000011011011011001",
			3478 => "0011001010000000000100",
			3479 => "0000001011011011011001",
			3480 => "0000000011011011011001",
			3481 => "1111111011011011011001",
			3482 => "0011010011011100000100",
			3483 => "0000000011011011011001",
			3484 => "0000001011011011011001",
			3485 => "0001111011000100010100",
			3486 => "0001000010010000001000",
			3487 => "0011011001110000000100",
			3488 => "0000000011011011011001",
			3489 => "1111111011011011011001",
			3490 => "0001100100110100001000",
			3491 => "0000001101111000000100",
			3492 => "0000001011011011011001",
			3493 => "0000000011011011011001",
			3494 => "0000000011011011011001",
			3495 => "0000011110100000010000",
			3496 => "0010100101000100000100",
			3497 => "1111111011011011011001",
			3498 => "0010100001010100000100",
			3499 => "0000001011011011011001",
			3500 => "0010010010001100000100",
			3501 => "1111111011011011011001",
			3502 => "0000000011011011011001",
			3503 => "0000000000101000000100",
			3504 => "0000001011011011011001",
			3505 => "0010111100001000000100",
			3506 => "0000000011011011011001",
			3507 => "0001001111100000000100",
			3508 => "0000000011011011011001",
			3509 => "1111111011011011011001",
			3510 => "0011000110000101111100",
			3511 => "0001000011111001111000",
			3512 => "0011000000101001000000",
			3513 => "0011000100010100100000",
			3514 => "0011000100010100010000",
			3515 => "0001111011000100001000",
			3516 => "0010110100000000000100",
			3517 => "0000000011100000011101",
			3518 => "0000001011100000011101",
			3519 => "0001110000101000000100",
			3520 => "0000000011100000011101",
			3521 => "0000000011100000011101",
			3522 => "0001111100001000001000",
			3523 => "0001111100001000000100",
			3524 => "0000000011100000011101",
			3525 => "0000001011100000011101",
			3526 => "0001111100001000000100",
			3527 => "1111111011100000011101",
			3528 => "0000000011100000011101",
			3529 => "0011000100010100010000",
			3530 => "0001111100001000001000",
			3531 => "0001110000101000000100",
			3532 => "0000001011100000011101",
			3533 => "0000000011100000011101",
			3534 => "0010111100001000000100",
			3535 => "0000010011100000011101",
			3536 => "0000001011100000011101",
			3537 => "0001000100001100001000",
			3538 => "0011000100010100000100",
			3539 => "1111111011100000011101",
			3540 => "0000000011100000011101",
			3541 => "0000011110100000000100",
			3542 => "0000001011100000011101",
			3543 => "1111111011100000011101",
			3544 => "0011000000101000011000",
			3545 => "0011011010111100010000",
			3546 => "0001101100011000001000",
			3547 => "0000100111111100000100",
			3548 => "0000000011100000011101",
			3549 => "1111111011100000011101",
			3550 => "0011100110000100000100",
			3551 => "1111111011100000011101",
			3552 => "0000001011100000011101",
			3553 => "0011010111001000000100",
			3554 => "1111110011100000011101",
			3555 => "1111111011100000011101",
			3556 => "0001100100110100010000",
			3557 => "0001000110001100001000",
			3558 => "0010101000010100000100",
			3559 => "0000000011100000011101",
			3560 => "0000001011100000011101",
			3561 => "0011100101101100000100",
			3562 => "0000000011100000011101",
			3563 => "1111111011100000011101",
			3564 => "0010100110011000001000",
			3565 => "0001000011001100000100",
			3566 => "0000001011100000011101",
			3567 => "0000000011100000011101",
			3568 => "0010011111001100000100",
			3569 => "0000000011100000011101",
			3570 => "0000000011100000011101",
			3571 => "1111111011100000011101",
			3572 => "0011001010111100100100",
			3573 => "0001111011000000011000",
			3574 => "0001110100011000010000",
			3575 => "0001111101111000001100",
			3576 => "0001111110001100000100",
			3577 => "1111111011100000011101",
			3578 => "0011000110000100000100",
			3579 => "0000000011100000011101",
			3580 => "0000000011100000011101",
			3581 => "1111111011100000011101",
			3582 => "0011000100001000000100",
			3583 => "0000010011100000011101",
			3584 => "1111111011100000011101",
			3585 => "0001000010010100000100",
			3586 => "1111111011100000011101",
			3587 => "0010100001010000000100",
			3588 => "0000010011100000011101",
			3589 => "0000000011100000011101",
			3590 => "1111111011100000011101",
			3591 => "0011000110000110101100",
			3592 => "0010101001000101101000",
			3593 => "0001001100001100101100",
			3594 => "0001001100001100100000",
			3595 => "0001001110000000010000",
			3596 => "0010001001101000001000",
			3597 => "0010100011101000000100",
			3598 => "0000000011100110010001",
			3599 => "0000000011100110010001",
			3600 => "0000101111010000000100",
			3601 => "0000000011100110010001",
			3602 => "1111110011100110010001",
			3603 => "0000001111000100001000",
			3604 => "0000011100110100000100",
			3605 => "0000000011100110010001",
			3606 => "1111111011100110010001",
			3607 => "0011101000111000000100",
			3608 => "0000000011100110010001",
			3609 => "0000000011100110010001",
			3610 => "0010010111100100001000",
			3611 => "0010110000101000000100",
			3612 => "0000010011100110010001",
			3613 => "1111111011100110010001",
			3614 => "0000001011100110010001",
			3615 => "0011111011011100011100",
			3616 => "0000011110100000001100",
			3617 => "0011101110111100001000",
			3618 => "0001110000101000000100",
			3619 => "0000000011100110010001",
			3620 => "1111111011100110010001",
			3621 => "0000010011100110010001",
			3622 => "0011000100010100001000",
			3623 => "0011110001011000000100",
			3624 => "0000000011100110010001",
			3625 => "1111111011100110010001",
			3626 => "0010001001101000000100",
			3627 => "0000000011100110010001",
			3628 => "0000010011100110010001",
			3629 => "0011011100101100010000",
			3630 => "0010110100010100001000",
			3631 => "0000000011111100000100",
			3632 => "1111111011100110010001",
			3633 => "0000001011100110010001",
			3634 => "0011100000101000000100",
			3635 => "1111111011100110010001",
			3636 => "1111111011100110010001",
			3637 => "0011000000101000001000",
			3638 => "0011101100101100000100",
			3639 => "0000000011100110010001",
			3640 => "1111111011100110010001",
			3641 => "0011000000101000000100",
			3642 => "1111111011100110010001",
			3643 => "0000000011100110010001",
			3644 => "0000001111000100010100",
			3645 => "0011010100011000000100",
			3646 => "1111110011100110010001",
			3647 => "0000100010000000000100",
			3648 => "0000001011100110010001",
			3649 => "0010001001101000001000",
			3650 => "0010001001101000000100",
			3651 => "1111111011100110010001",
			3652 => "0000000011100110010001",
			3653 => "1111111011100110010001",
			3654 => "0001000011001100010000",
			3655 => "0000000000110000001100",
			3656 => "0000010110000000000100",
			3657 => "1111111011100110010001",
			3658 => "0011001010000000000100",
			3659 => "1111111011100110010001",
			3660 => "0000000011100110010001",
			3661 => "1111111011100110010001",
			3662 => "0001111100001000010000",
			3663 => "0001110000101000001000",
			3664 => "0001110000101000000100",
			3665 => "0000000011100110010001",
			3666 => "0000000011100110010001",
			3667 => "0011111011011100000100",
			3668 => "0000001011100110010001",
			3669 => "0000000011100110010001",
			3670 => "0010000110001000001000",
			3671 => "0011111001010100000100",
			3672 => "0000000011100110010001",
			3673 => "1111111011100110010001",
			3674 => "0001111100001000000100",
			3675 => "0000000011100110010001",
			3676 => "0000000011100110010001",
			3677 => "0011001010111100001100",
			3678 => "0000000111000100001000",
			3679 => "0000001111001000000100",
			3680 => "1111111011100110010001",
			3681 => "0000001011100110010001",
			3682 => "1111111011100110010001",
			3683 => "1111111011100110010001",
			3684 => "0000110100000010000000",
			3685 => "0001000011010100111000",
			3686 => "0000000100010100101000",
			3687 => "0000110100000000011000",
			3688 => "0000101111010000010000",
			3689 => "0011110100000100001000",
			3690 => "0010000111000100000100",
			3691 => "0000000011101110000101",
			3692 => "0000000011101110000101",
			3693 => "0001011001110000000100",
			3694 => "1111111011101110000101",
			3695 => "0000001011101110000101",
			3696 => "0011011001110000000100",
			3697 => "0000000011101110000101",
			3698 => "1111111011101110000101",
			3699 => "0001110111111000000100",
			3700 => "0000000011101110000101",
			3701 => "0011110100000100001000",
			3702 => "0011010101101100000100",
			3703 => "0000000011101110000101",
			3704 => "1111111011101110000101",
			3705 => "1111111011101110000101",
			3706 => "0001100100110100000100",
			3707 => "1111111011101110000101",
			3708 => "0011011101100000000100",
			3709 => "0000001011101110000101",
			3710 => "0011011100101100000100",
			3711 => "1111111011101110000101",
			3712 => "0000000011101110000101",
			3713 => "0001000011110100010100",
			3714 => "0000011110100000010000",
			3715 => "0010101100011100001100",
			3716 => "0010000001110100001000",
			3717 => "0001101101111100000100",
			3718 => "0000001011101110000101",
			3719 => "0000000011101110000101",
			3720 => "0000000011101110000101",
			3721 => "0000001011101110000101",
			3722 => "1111111011101110000101",
			3723 => "0000010110000000011100",
			3724 => "0011111110110000010000",
			3725 => "0011010100000000001000",
			3726 => "0011001010000000000100",
			3727 => "0000000011101110000101",
			3728 => "0000000011101110000101",
			3729 => "0000101100100100000100",
			3730 => "1111111011101110000101",
			3731 => "0000000011101110000101",
			3732 => "0011000100010100001000",
			3733 => "0011110000011100000100",
			3734 => "0000001011101110000101",
			3735 => "0000000011101110000101",
			3736 => "1111111011101110000101",
			3737 => "0000101100100100001100",
			3738 => "0000110111111000001000",
			3739 => "0010100101000100000100",
			3740 => "1111111011101110000101",
			3741 => "0000000011101110000101",
			3742 => "0000001011101110000101",
			3743 => "0010010110101000001000",
			3744 => "0001000011011000000100",
			3745 => "0000000011101110000101",
			3746 => "0000000011101110000101",
			3747 => "0000001011101110000101",
			3748 => "0010010010001100010100",
			3749 => "0001100001111000000100",
			3750 => "1111111011101110000101",
			3751 => "0001101101111100000100",
			3752 => "0000001011101110000101",
			3753 => "0001100100110100000100",
			3754 => "0000000011101110000101",
			3755 => "0000111001110000000100",
			3756 => "0000000011101110000101",
			3757 => "0000001011101110000101",
			3758 => "0011110001011000101100",
			3759 => "0010010110101000010000",
			3760 => "0000011110100000001100",
			3761 => "0001010101101100001000",
			3762 => "0001111011000100000100",
			3763 => "0000000011101110000101",
			3764 => "0000001011101110000101",
			3765 => "1111111011101110000101",
			3766 => "0000001011101110000101",
			3767 => "0011011110001100010000",
			3768 => "0011110000011100001000",
			3769 => "0010001001101000000100",
			3770 => "1111111011101110000101",
			3771 => "0000000011101110000101",
			3772 => "0000110011011100000100",
			3773 => "0000001011101110000101",
			3774 => "0000000011101110000101",
			3775 => "0011000111111000000100",
			3776 => "1111111011101110000101",
			3777 => "0011011101111000000100",
			3778 => "0000001011101110000101",
			3779 => "0000000011101110000101",
			3780 => "0001101101111100100000",
			3781 => "0000111110001100010000",
			3782 => "0001011100101100001000",
			3783 => "0001000010111000000100",
			3784 => "0000000011101110000101",
			3785 => "0000000011101110000101",
			3786 => "0001001110000000000100",
			3787 => "0000000011101110000101",
			3788 => "1111111011101110000101",
			3789 => "0000111010111100001000",
			3790 => "0011000100000000000100",
			3791 => "0000000011101110000101",
			3792 => "1111111011101110000101",
			3793 => "0000011001111000000100",
			3794 => "1111111011101110000101",
			3795 => "0000000011101110000101",
			3796 => "0000101100100100001100",
			3797 => "0001011110001100000100",
			3798 => "1111111011101110000101",
			3799 => "0010001100000100000100",
			3800 => "1111111011101110000101",
			3801 => "0000000011101110000101",
			3802 => "0011010101101100001000",
			3803 => "0000100101001000000100",
			3804 => "0000001011101110000101",
			3805 => "0000000011101110000101",
			3806 => "0000110011011100000100",
			3807 => "0000000011101110000101",
			3808 => "0000000011101110000101",
			3809 => "0000100110010010010100",
			3810 => "0001000011011001010100",
			3811 => "0000001100001000110100",
			3812 => "0001011000111100010100",
			3813 => "0001011000111100010000",
			3814 => "0000101110000100001000",
			3815 => "0001100001111000000100",
			3816 => "0000000011110111000001",
			3817 => "1111111011110111000001",
			3818 => "0000110100010100000100",
			3819 => "0000001011110111000001",
			3820 => "0000001011110111000001",
			3821 => "0000010011110111000001",
			3822 => "0010110111111000010000",
			3823 => "0001000000010100001000",
			3824 => "0011011101100000000100",
			3825 => "1111111011110111000001",
			3826 => "0000000011110111000001",
			3827 => "0001110111111000000100",
			3828 => "0000000011110111000001",
			3829 => "1111111011110111000001",
			3830 => "0010011001111000001000",
			3831 => "0000111100001000000100",
			3832 => "0000000011110111000001",
			3833 => "0000001011110111000001",
			3834 => "0001100100110100000100",
			3835 => "0000000011110111000001",
			3836 => "0000000011110111000001",
			3837 => "0011100000101000011000",
			3838 => "0010110111111000001100",
			3839 => "0001011000111100001000",
			3840 => "0001011000111100000100",
			3841 => "1111111011110111000001",
			3842 => "0000000011110111000001",
			3843 => "0000001011110111000001",
			3844 => "0010100001010100001000",
			3845 => "0001110000101000000100",
			3846 => "1111111011110111000001",
			3847 => "0000000011110111000001",
			3848 => "0000000011110111000001",
			3849 => "0011100100000000000100",
			3850 => "0000010011110111000001",
			3851 => "1111111011110111000001",
			3852 => "0001000001100100100100",
			3853 => "0010100110011100001100",
			3854 => "0010110111111000001000",
			3855 => "0001111010000000000100",
			3856 => "0000000011110111000001",
			3857 => "0000010011110111000001",
			3858 => "1111111011110111000001",
			3859 => "0010100101000100001000",
			3860 => "0011000100010100000100",
			3861 => "0000001011110111000001",
			3862 => "0000010011110111000001",
			3863 => "0001000000100000001000",
			3864 => "0010001000110000000100",
			3865 => "1111111011110111000001",
			3866 => "0000000011110111000001",
			3867 => "0000100001000000000100",
			3868 => "0000001011110111000001",
			3869 => "0000000011110111000001",
			3870 => "0000101001010000001100",
			3871 => "0001011000111100001000",
			3872 => "0011100101000100000100",
			3873 => "1111111011110111000001",
			3874 => "0000001011110111000001",
			3875 => "1111111011110111000001",
			3876 => "0000101010001000001100",
			3877 => "0011100010101000001000",
			3878 => "0001100100110100000100",
			3879 => "0000001011110111000001",
			3880 => "1111111011110111000001",
			3881 => "0000001011110111000001",
			3882 => "1111111011110111000001",
			3883 => "0001101010011001000000",
			3884 => "0001011101100000010100",
			3885 => "0001001011100000001000",
			3886 => "0000000011111100000100",
			3887 => "0000000011110111000001",
			3888 => "0000001011110111000001",
			3889 => "0000000000101000001000",
			3890 => "0001110111111000000100",
			3891 => "0000000011110111000001",
			3892 => "0000000011110111000001",
			3893 => "1111111011110111000001",
			3894 => "0001111000111000011000",
			3895 => "0011000100000000010000",
			3896 => "0001011100101000001000",
			3897 => "0010111000111100000100",
			3898 => "0000000011110111000001",
			3899 => "1111111011110111000001",
			3900 => "0000101001100000000100",
			3901 => "0000001011110111000001",
			3902 => "0000000011110111000001",
			3903 => "0000101110110100000100",
			3904 => "1111111011110111000001",
			3905 => "1111111011110111000001",
			3906 => "0000000011111100001100",
			3907 => "0000101110110100000100",
			3908 => "1111111011110111000001",
			3909 => "0001101010011000000100",
			3910 => "0000000011110111000001",
			3911 => "0000001011110111000001",
			3912 => "0001001111100000000100",
			3913 => "0000001011110111000001",
			3914 => "1111111011110111000001",
			3915 => "0001101010011000001100",
			3916 => "0001110101101100000100",
			3917 => "0000001011110111000001",
			3918 => "0010011010011000000100",
			3919 => "1111111011110111000001",
			3920 => "0000000011110111000001",
			3921 => "0010001111001000100000",
			3922 => "0001101101011000010000",
			3923 => "0001000010110000001000",
			3924 => "0000100010000100000100",
			3925 => "0000000011110111000001",
			3926 => "1111111011110111000001",
			3927 => "0000100111011000000100",
			3928 => "1111111011110111000001",
			3929 => "0000000011110111000001",
			3930 => "0000110000011100001000",
			3931 => "0011000100000000000100",
			3932 => "0000000011110111000001",
			3933 => "0000001011110111000001",
			3934 => "0001011000011000000100",
			3935 => "1111111011110111000001",
			3936 => "0000000011110111000001",
			3937 => "0001001001001100010000",
			3938 => "0001111001110000001000",
			3939 => "0011000100000000000100",
			3940 => "0000000011110111000001",
			3941 => "0000001011110111000001",
			3942 => "0010000111000100000100",
			3943 => "0000001011110111000001",
			3944 => "1111111011110111000001",
			3945 => "0000001110111100001000",
			3946 => "0000101100010000000100",
			3947 => "1111111011110111000001",
			3948 => "0000000011110111000001",
			3949 => "0001000100001100000100",
			3950 => "0000000011110111000001",
			3951 => "0000000011110111000001",
			3952 => "0011001000111010111000",
			3953 => "0011000111111001101100",
			3954 => "0011000111111001000000",
			3955 => "0011000111111000100000",
			3956 => "0000101110010000010000",
			3957 => "0001110100010100001000",
			3958 => "0001110100010100000100",
			3959 => "0000000011111110111101",
			3960 => "0000000011111110111101",
			3961 => "0000101001010000000100",
			3962 => "0000000011111110111101",
			3963 => "1111111011111110111101",
			3964 => "0001001011100000001000",
			3965 => "0011111011110100000100",
			3966 => "0000010011111110111101",
			3967 => "0000000011111110111101",
			3968 => "0001100100110100000100",
			3969 => "0000000011111110111101",
			3970 => "1111111011111110111101",
			3971 => "0011000111111000010000",
			3972 => "0010010110101000001000",
			3973 => "0011011001110000000100",
			3974 => "0000000011111110111101",
			3975 => "0000001011111110111101",
			3976 => "0011011110001100000100",
			3977 => "0000000011111110111101",
			3978 => "0000001011111110111101",
			3979 => "0001110100010100001000",
			3980 => "0001110111111000000100",
			3981 => "0000000011111110111101",
			3982 => "0000010011111110111101",
			3983 => "0001110100010100000100",
			3984 => "1111111011111110111101",
			3985 => "0000000011111110111101",
			3986 => "0011000111111000010000",
			3987 => "0001110111111000000100",
			3988 => "0000001011111110111101",
			3989 => "0010010111100100001000",
			3990 => "0000110101101100000100",
			3991 => "0000000011111110111101",
			3992 => "1111111011111110111101",
			3993 => "0000000011111110111101",
			3994 => "0001110000101000010000",
			3995 => "0001110111111000001000",
			3996 => "0000010110000000000100",
			3997 => "0000000011111110111101",
			3998 => "1111111011111110111101",
			3999 => "0000100010110100000100",
			4000 => "1111111011111110111101",
			4001 => "0000000011111110111101",
			4002 => "0001110000101000000100",
			4003 => "1111111011111110111101",
			4004 => "0010110000101000000100",
			4005 => "0000000011111110111101",
			4006 => "0000000011111110111101",
			4007 => "0011000100010100100000",
			4008 => "0000001000110000000100",
			4009 => "1111111011111110111101",
			4010 => "0000011100110100010000",
			4011 => "0001110000101000001000",
			4012 => "0011011100110000000100",
			4013 => "0000000011111110111101",
			4014 => "0000001011111110111101",
			4015 => "0000000000111000000100",
			4016 => "1111111011111110111101",
			4017 => "0000000011111110111101",
			4018 => "0010111000111100001000",
			4019 => "0000110110000100000100",
			4020 => "0000001011111110111101",
			4021 => "0000001011111110111101",
			4022 => "0000000011111110111101",
			4023 => "0000010110000000010000",
			4024 => "0000110011010000001000",
			4025 => "0000101110101000000100",
			4026 => "0000000011111110111101",
			4027 => "0000001011111110111101",
			4028 => "0011010101101100000100",
			4029 => "1111111011111110111101",
			4030 => "0000000011111110111101",
			4031 => "0011011101100000001100",
			4032 => "0011000100010100000100",
			4033 => "1111111011111110111101",
			4034 => "0000101001010000000100",
			4035 => "0000001011111110111101",
			4036 => "0000000011111110111101",
			4037 => "0000111100110000001000",
			4038 => "0011011101111000000100",
			4039 => "0000000011111110111101",
			4040 => "1111111011111110111101",
			4041 => "0010010111100100000100",
			4042 => "0000000011111110111101",
			4043 => "0000000011111110111101",
			4044 => "0011111101000100001100",
			4045 => "0000000011010000001000",
			4046 => "0010111100101100000100",
			4047 => "0000000011111110111101",
			4048 => "1111111011111110111101",
			4049 => "1111111011111110111101",
			4050 => "0000010110101000011100",
			4051 => "0001011001110100010000",
			4052 => "0010100110011100001100",
			4053 => "0010101010110000001000",
			4054 => "0010100001010000000100",
			4055 => "1111111011111110111101",
			4056 => "0000001011111110111101",
			4057 => "1111111011111110111101",
			4058 => "0000001011111110111101",
			4059 => "0010110001111100001000",
			4060 => "0000110001101000000100",
			4061 => "0000000011111110111101",
			4062 => "0000001011111110111101",
			4063 => "0000000011111110111101",
			4064 => "0000000111000100010000",
			4065 => "0011001010111100001100",
			4066 => "0000001001101000000100",
			4067 => "0000000011111110111101",
			4068 => "0000011110010100000100",
			4069 => "0000001011111110111101",
			4070 => "0000000011111110111101",
			4071 => "1111111011111110111101",
			4072 => "0001111110001100000100",
			4073 => "1111111011111110111101",
			4074 => "0001111101111000001000",
			4075 => "0000101011101100000100",
			4076 => "0000001011111110111101",
			4077 => "0000000011111110111101",
			4078 => "1111111011111110111101",
			4079 => "0010100001010010010000",
			4080 => "0010001111001001110000",
			4081 => "0000000011010000111000",
			4082 => "0000100110010000100000",
			4083 => "0010101001000100010000",
			4084 => "0001101010011000001000",
			4085 => "0000011001111000000100",
			4086 => "0000000100000111111001",
			4087 => "0000000100000111111001",
			4088 => "0001010100011000000100",
			4089 => "1111111100000111111001",
			4090 => "0000000100000111111001",
			4091 => "0001101101111100001000",
			4092 => "0011100100010100000100",
			4093 => "0000000100000111111001",
			4094 => "0000001100000111111001",
			4095 => "0000111110001100000100",
			4096 => "1111111100000111111001",
			4097 => "0000000100000111111001",
			4098 => "0011110101001000001000",
			4099 => "0001110100000000000100",
			4100 => "0000000100000111111001",
			4101 => "1111111100000111111001",
			4102 => "0010100110011000001000",
			4103 => "0010100110011000000100",
			4104 => "0000000100000111111001",
			4105 => "0000001100000111111001",
			4106 => "0001011000011000000100",
			4107 => "1111111100000111111001",
			4108 => "0000001100000111111001",
			4109 => "0010111100001000011000",
			4110 => "0010111100001000010000",
			4111 => "0000000000111000001000",
			4112 => "0010000110001000000100",
			4113 => "0000000100000111111001",
			4114 => "0000001100000111111001",
			4115 => "0010001111001000000100",
			4116 => "0000000100000111111001",
			4117 => "0000001100000111111001",
			4118 => "0010000110001000000100",
			4119 => "0000000100000111111001",
			4120 => "0000001100000111111001",
			4121 => "0011100100000000010000",
			4122 => "0011011110001100001000",
			4123 => "0000100101110000000100",
			4124 => "0000000100000111111001",
			4125 => "1111111100000111111001",
			4126 => "0001100100110100000100",
			4127 => "1111111100000111111001",
			4128 => "0000000100000111111001",
			4129 => "0010011011101000001000",
			4130 => "0011011101111000000100",
			4131 => "0000000100000111111001",
			4132 => "0000000100000111111001",
			4133 => "0010110110000100000100",
			4134 => "1111111100000111111001",
			4135 => "0000000100000111111001",
			4136 => "0011011100110000010100",
			4137 => "0001010011011100010000",
			4138 => "0000010110000000001000",
			4139 => "0000000000101000000100",
			4140 => "0000001100000111111001",
			4141 => "0000000100000111111001",
			4142 => "0000001110111100000100",
			4143 => "0000000100000111111001",
			4144 => "1111111100000111111001",
			4145 => "0000000100000111111001",
			4146 => "0001111100001000000100",
			4147 => "1111111100000111111001",
			4148 => "0011110111110000000100",
			4149 => "0000000100000111111001",
			4150 => "1111111100000111111001",
			4151 => "0000111110111100110100",
			4152 => "0010100101000100011000",
			4153 => "0010011100110100010000",
			4154 => "0011110100011000000100",
			4155 => "1111111100000111111001",
			4156 => "0001011000111100001000",
			4157 => "0000110011111100000100",
			4158 => "0000000100000111111001",
			4159 => "0000001100000111111001",
			4160 => "0000000100000111111001",
			4161 => "0011111010111000000100",
			4162 => "0000000100000111111001",
			4163 => "1111111100000111111001",
			4164 => "0001101010011000011000",
			4165 => "0000001100110000001000",
			4166 => "0010001000110000000100",
			4167 => "0000000100000111111001",
			4168 => "0000001100000111111001",
			4169 => "0000110000110000001000",
			4170 => "0001011001110000000100",
			4171 => "0000000100000111111001",
			4172 => "1111111100000111111001",
			4173 => "0000100110010000000100",
			4174 => "0000001100000111111001",
			4175 => "0000000100000111111001",
			4176 => "1111111100000111111001",
			4177 => "0000101111010000101000",
			4178 => "0000001011000100011000",
			4179 => "0011101101010000001000",
			4180 => "0000101100100100000100",
			4181 => "0000010100000111111001",
			4182 => "0000000100000111111001",
			4183 => "0010000001110100001000",
			4184 => "0000011110100000000100",
			4185 => "0000000100000111111001",
			4186 => "0000000100000111111001",
			4187 => "0011110111010000000100",
			4188 => "0000001100000111111001",
			4189 => "0000000100000111111001",
			4190 => "0000111011000100001000",
			4191 => "0000010110000000000100",
			4192 => "0000000100000111111001",
			4193 => "1111111100000111111001",
			4194 => "0000011110100000000100",
			4195 => "0000001100000111111001",
			4196 => "1111111100000111111001",
			4197 => "0000101001010000010100",
			4198 => "0001100100110100001000",
			4199 => "0000101111010000000100",
			4200 => "1111111100000111111001",
			4201 => "0000000100000111111001",
			4202 => "0000011110100000000100",
			4203 => "0000001100000111111001",
			4204 => "0000011100110100000100",
			4205 => "1111111100000111111001",
			4206 => "0000000100000111111001",
			4207 => "0011011100110000010000",
			4208 => "0011100111111000001000",
			4209 => "0001110111111000000100",
			4210 => "0000000100000111111001",
			4211 => "0000000100000111111001",
			4212 => "0000111101100000000100",
			4213 => "1111111100000111111001",
			4214 => "0000000100000111111001",
			4215 => "0010010111100100001000",
			4216 => "0000110101101100000100",
			4217 => "0000000100000111111001",
			4218 => "0000000100000111111001",
			4219 => "0000011100110100000100",
			4220 => "0000000100000111111001",
			4221 => "0000000100000111111001",
			4222 => "0010100110011010101100",
			4223 => "0011000100010101010000",
			4224 => "0001111011000100100000",
			4225 => "0001011100101100011000",
			4226 => "0001101101111100001100",
			4227 => "0001111011000100001000",
			4228 => "0001111011000100000100",
			4229 => "0000000100010000011101",
			4230 => "1111111100010000011101",
			4231 => "0000001100010000011101",
			4232 => "0010111100001000001000",
			4233 => "0001000010110000000100",
			4234 => "1111111100010000011101",
			4235 => "0000000100010000011101",
			4236 => "0000000100010000011101",
			4237 => "0001111011000100000100",
			4238 => "0000000100010000011101",
			4239 => "0000001100010000011101",
			4240 => "0011000100010100100000",
			4241 => "0000011100110100010000",
			4242 => "0001000011001100001000",
			4243 => "0000000010111100000100",
			4244 => "0000000100010000011101",
			4245 => "0000000100010000011101",
			4246 => "0001000010111000000100",
			4247 => "1111111100010000011101",
			4248 => "0000000100010000011101",
			4249 => "0010111000111100001000",
			4250 => "0001100100110100000100",
			4251 => "1111111100010000011101",
			4252 => "0000000100010000011101",
			4253 => "0001111100001000000100",
			4254 => "0000000100010000011101",
			4255 => "0000001100010000011101",
			4256 => "0001111100001000001000",
			4257 => "0000011100110100000100",
			4258 => "1111111100010000011101",
			4259 => "1111111100010000011101",
			4260 => "0010110100000000000100",
			4261 => "0000000100010000011101",
			4262 => "1111111100010000011101",
			4263 => "0011000100010100100100",
			4264 => "0000011110100000010000",
			4265 => "0010111011000100001000",
			4266 => "0010011001111000000100",
			4267 => "0000000100010000011101",
			4268 => "1111111100010000011101",
			4269 => "0001110000101000000100",
			4270 => "0000001100010000011101",
			4271 => "1111111100010000011101",
			4272 => "0010111000111100001100",
			4273 => "0000111101111000001000",
			4274 => "0000111001110000000100",
			4275 => "0000001100010000011101",
			4276 => "0000000100010000011101",
			4277 => "0000001100010000011101",
			4278 => "0001110100000000000100",
			4279 => "0000000100010000011101",
			4280 => "1111111100010000011101",
			4281 => "0000100110100000011000",
			4282 => "0000110100000000001000",
			4283 => "0011010110000100000100",
			4284 => "1111111100010000011101",
			4285 => "0000000100010000011101",
			4286 => "0010100011101000001000",
			4287 => "0000111010011100000100",
			4288 => "1111111100010000011101",
			4289 => "0000000100010000011101",
			4290 => "0011000000101000000100",
			4291 => "0000000100010000011101",
			4292 => "0000001100010000011101",
			4293 => "0000101100100100010000",
			4294 => "0000101110101000001000",
			4295 => "0000101110101000000100",
			4296 => "0000000100010000011101",
			4297 => "0000001100010000011101",
			4298 => "0010101000100100000100",
			4299 => "0000000100010000011101",
			4300 => "1111111100010000011101",
			4301 => "0011010000001100001000",
			4302 => "0000011100110100000100",
			4303 => "0000000100010000011101",
			4304 => "0000001100010000011101",
			4305 => "0001010000001100000100",
			4306 => "1111111100010000011101",
			4307 => "0000000100010000011101",
			4308 => "0010100110011000011000",
			4309 => "0011000100010100000100",
			4310 => "1111111100010000011101",
			4311 => "0011011100101100000100",
			4312 => "0000010100010000011101",
			4313 => "0001001101001000001100",
			4314 => "0001100100110100000100",
			4315 => "0000000100010000011101",
			4316 => "0000001111000100000100",
			4317 => "0000000100010000011101",
			4318 => "0000001100010000011101",
			4319 => "1111111100010000011101",
			4320 => "0011000000111000011000",
			4321 => "0000100110100000000100",
			4322 => "1111111100010000011101",
			4323 => "0001100001111000000100",
			4324 => "0000000100010000011101",
			4325 => "0011000000111000001000",
			4326 => "0000011110011100000100",
			4327 => "0000000100010000011101",
			4328 => "0000000100010000011101",
			4329 => "0000001101111000000100",
			4330 => "0000001100010000011101",
			4331 => "0000000100010000011101",
			4332 => "0000111011000100011100",
			4333 => "0001000100001100010000",
			4334 => "0011001010000000001000",
			4335 => "0011001010000000000100",
			4336 => "1111111100010000011101",
			4337 => "0000001100010000011101",
			4338 => "0010101010110000000100",
			4339 => "1111111100010000011101",
			4340 => "0000000100010000011101",
			4341 => "0000000100010100000100",
			4342 => "0000001100010000011101",
			4343 => "0001001111100000000100",
			4344 => "1111111100010000011101",
			4345 => "0000000100010000011101",
			4346 => "0010001001101000001100",
			4347 => "0001001011110000001000",
			4348 => "0001011000000000000100",
			4349 => "0000000100010000011101",
			4350 => "0000001100010000011101",
			4351 => "1111111100010000011101",
			4352 => "0000101110000100001000",
			4353 => "0000101110000100000100",
			4354 => "0000000100010000011101",
			4355 => "0000001100010000011101",
			4356 => "0001000101010100000100",
			4357 => "0000000100010000011101",
			4358 => "0000000100010000011101",
			4359 => "0010110110000110111100",
			4360 => "0001000100001101100000",
			4361 => "0011100111111000100100",
			4362 => "0001000110101100000100",
			4363 => "1110100100011001100001",
			4364 => "0001101101111100010000",
			4365 => "0001100111101000001000",
			4366 => "0010110100010100000100",
			4367 => "1110000100011001100001",
			4368 => "1101111100011001100001",
			4369 => "0000110100010100000100",
			4370 => "1110000100011001100001",
			4371 => "1110000100011001100001",
			4372 => "0000000000111000001000",
			4373 => "0010011001111000000100",
			4374 => "1110101100011001100001",
			4375 => "1110010100011001100001",
			4376 => "0001010110000100000100",
			4377 => "1110001100011001100001",
			4378 => "1101111100011001100001",
			4379 => "0001100111101000011100",
			4380 => "0010000001010100010000",
			4381 => "0010100011101000001000",
			4382 => "0001101011111100000100",
			4383 => "1101111100011001100001",
			4384 => "1101111100011001100001",
			4385 => "0001000110111000000100",
			4386 => "1110010100011001100001",
			4387 => "1101111100011001100001",
			4388 => "0010010110101000001000",
			4389 => "0001001100001100000100",
			4390 => "1110100100011001100001",
			4391 => "1110000100011001100001",
			4392 => "1101111100011001100001",
			4393 => "0001001101001000010000",
			4394 => "0001101101111100001000",
			4395 => "0000101100100100000100",
			4396 => "1110100100011001100001",
			4397 => "1110010100011001100001",
			4398 => "0001111001110000000100",
			4399 => "1110100100011001100001",
			4400 => "1110001100011001100001",
			4401 => "0001110000101000001000",
			4402 => "0001101100011000000100",
			4403 => "1110011100011001100001",
			4404 => "1110101100011001100001",
			4405 => "0011100110000100000100",
			4406 => "1110001100011001100001",
			4407 => "1110010100011001100001",
			4408 => "0001101101111100011100",
			4409 => "0001000011110100001100",
			4410 => "0000001010000000000100",
			4411 => "1101111100011001100001",
			4412 => "0000000100010100000100",
			4413 => "1110011100011001100001",
			4414 => "1110000100011001100001",
			4415 => "0000010000011000000100",
			4416 => "1101111100011001100001",
			4417 => "0001000011101100000100",
			4418 => "1101111100011001100001",
			4419 => "0010010010001100000100",
			4420 => "1110000100011001100001",
			4421 => "1101111100011001100001",
			4422 => "0010011001111000100000",
			4423 => "0000001011000100010000",
			4424 => "0000111001110000001000",
			4425 => "0001001111100000000100",
			4426 => "1110001100011001100001",
			4427 => "1110010100011001100001",
			4428 => "0001111011000100000100",
			4429 => "1110100100011001100001",
			4430 => "1110010100011001100001",
			4431 => "0001001011100000001000",
			4432 => "0000111100001000000100",
			4433 => "1101111100011001100001",
			4434 => "1110001100011001100001",
			4435 => "0001000011111000000100",
			4436 => "1110001100011001100001",
			4437 => "1101111100011001100001",
			4438 => "0011100110000100010000",
			4439 => "0001010110000100001000",
			4440 => "0000000100010100000100",
			4441 => "1110001100011001100001",
			4442 => "1110000100011001100001",
			4443 => "0000101111010000000100",
			4444 => "1110001100011001100001",
			4445 => "1101111100011001100001",
			4446 => "0001000011010100001000",
			4447 => "0010000001110100000100",
			4448 => "1110000100011001100001",
			4449 => "1110100100011001100001",
			4450 => "0011111001010000000100",
			4451 => "1110000100011001100001",
			4452 => "1110010100011001100001",
			4453 => "0001110101101100111100",
			4454 => "0001101001100100101000",
			4455 => "0000110001101000010000",
			4456 => "0001011010111000000100",
			4457 => "1110001100011001100001",
			4458 => "0000111000000000000100",
			4459 => "1101111100011001100001",
			4460 => "0001111101100000000100",
			4461 => "1110001100011001100001",
			4462 => "1101111100011001100001",
			4463 => "0010101000010100001000",
			4464 => "0001101101111100000100",
			4465 => "1110010100011001100001",
			4466 => "1110101100011001100001",
			4467 => "0010010101011100001000",
			4468 => "0010111101111000000100",
			4469 => "1110001100011001100001",
			4470 => "1110011100011001100001",
			4471 => "0000000010111100000100",
			4472 => "1101111100011001100001",
			4473 => "1110000100011001100001",
			4474 => "0001101001100100010000",
			4475 => "0001111001110000000100",
			4476 => "1110001100011001100001",
			4477 => "0011111001011100000100",
			4478 => "1101111100011001100001",
			4479 => "0000010111100100000100",
			4480 => "1101111100011001100001",
			4481 => "1110000100011001100001",
			4482 => "1101111100011001100001",
			4483 => "0001111101111000011100",
			4484 => "0011101001001000001100",
			4485 => "0010111110001100001000",
			4486 => "0001010011100000000100",
			4487 => "1101111100011001100001",
			4488 => "1110000100011001100001",
			4489 => "1101111100011001100001",
			4490 => "0000100111010100001100",
			4491 => "0000001011010100000100",
			4492 => "1101111100011001100001",
			4493 => "0010110100001000000100",
			4494 => "1110000100011001100001",
			4495 => "1110100100011001100001",
			4496 => "1101111100011001100001",
			4497 => "0010000110011100001100",
			4498 => "0010100010101100000100",
			4499 => "1101111100011001100001",
			4500 => "0010001100011100000100",
			4501 => "1101111100011001100001",
			4502 => "1101111100011001100001",
			4503 => "1101111100011001100001",
			4504 => "0010001001101010101000",
			4505 => "0010001001101001100100",
			4506 => "0011010101101100101100",
			4507 => "0001110100010100011100",
			4508 => "0011000111111000010000",
			4509 => "0000111011000100001000",
			4510 => "0001111110111100000100",
			4511 => "0000000100100010110101",
			4512 => "0000001100100010110101",
			4513 => "0000111000111000000100",
			4514 => "0000000100100010110101",
			4515 => "0000001100100010110101",
			4516 => "0011011100110000001000",
			4517 => "0010010010001100000100",
			4518 => "0000000100100010110101",
			4519 => "1111111100100010110101",
			4520 => "0000000100100010110101",
			4521 => "0000101101000100001100",
			4522 => "0000110100010100000100",
			4523 => "0000000100100010110101",
			4524 => "0011100000110000000100",
			4525 => "0000010100100010110101",
			4526 => "0000001100100010110101",
			4527 => "0000000100100010110101",
			4528 => "0011101000111100011000",
			4529 => "0001110100010100001000",
			4530 => "0000011110100000000100",
			4531 => "0000000100100010110101",
			4532 => "0000001100100010110101",
			4533 => "0010110000101000001000",
			4534 => "0000000010111100000100",
			4535 => "1111111100100010110101",
			4536 => "0000000100100010110101",
			4537 => "0010111100001000000100",
			4538 => "0000000100100010110101",
			4539 => "0000000100100010110101",
			4540 => "0001110000101000010000",
			4541 => "0000100101001000001000",
			4542 => "0001011100101100000100",
			4543 => "0000000100100010110101",
			4544 => "0000001100100010110101",
			4545 => "0001000110001100000100",
			4546 => "0000001100100010110101",
			4547 => "0000010100100010110101",
			4548 => "0001000110001100001000",
			4549 => "0000001111000100000100",
			4550 => "0000000100100010110101",
			4551 => "0000000100100010110101",
			4552 => "0011010001111100000100",
			4553 => "0000000100100010110101",
			4554 => "1111111100100010110101",
			4555 => "0000100101110000100100",
			4556 => "0010101000010100010000",
			4557 => "0000000011111100001100",
			4558 => "0010101000010100000100",
			4559 => "0000000100100010110101",
			4560 => "0010111100001000000100",
			4561 => "1111111100100010110101",
			4562 => "0000000100100010110101",
			4563 => "0000000100100010110101",
			4564 => "0000001111000100000100",
			4565 => "1111111100100010110101",
			4566 => "0000110110000100001000",
			4567 => "0000100111100000000100",
			4568 => "0000000100100010110101",
			4569 => "1111111100100010110101",
			4570 => "0011000000101000000100",
			4571 => "0000001100100010110101",
			4572 => "0000000100100010110101",
			4573 => "0000011001111000010000",
			4574 => "0011101010111100001100",
			4575 => "0011101101111000001000",
			4576 => "0000101100010100000100",
			4577 => "1111111100100010110101",
			4578 => "0000001100100010110101",
			4579 => "0000001100100010110101",
			4580 => "1111110100100010110101",
			4581 => "0010100110011000001100",
			4582 => "0000100010000100001000",
			4583 => "0011101010111000000100",
			4584 => "1111111100100010110101",
			4585 => "0000001100100010110101",
			4586 => "1111111100100010110101",
			4587 => "1111111100100010110101",
			4588 => "0010001011010100101100",
			4589 => "0000101110010000011100",
			4590 => "0011001010000000000100",
			4591 => "0000001100100010110101",
			4592 => "0010101001000100001000",
			4593 => "0010101001000100000100",
			4594 => "0000000100100010110101",
			4595 => "1111111100100010110101",
			4596 => "0001011100101100001000",
			4597 => "0000011100110100000100",
			4598 => "0000001100100010110101",
			4599 => "1111111100100010110101",
			4600 => "0011010100001000000100",
			4601 => "0000001100100010110101",
			4602 => "0000001100100010110101",
			4603 => "0000101110110100001000",
			4604 => "0000011001111000000100",
			4605 => "0000000100100010110101",
			4606 => "1111110100100010110101",
			4607 => "0001110110000100000100",
			4608 => "0000001100100010110101",
			4609 => "0000000100100010110101",
			4610 => "0010001011010100011000",
			4611 => "0000000011010000010100",
			4612 => "0001000010111000001100",
			4613 => "0011100000101000000100",
			4614 => "0000001100100010110101",
			4615 => "0011101110001100000100",
			4616 => "1111111100100010110101",
			4617 => "0000000100100010110101",
			4618 => "0000000011111100000100",
			4619 => "0000000100100010110101",
			4620 => "0000010100100010110101",
			4621 => "1111111100100010110101",
			4622 => "0000000000111000100000",
			4623 => "0010001011010100010000",
			4624 => "0010100110011000001000",
			4625 => "0000011100110100000100",
			4626 => "0000000100100010110101",
			4627 => "1111111100100010110101",
			4628 => "0001000011001100000100",
			4629 => "0000001100100010110101",
			4630 => "0000000100100010110101",
			4631 => "0000101001011100001000",
			4632 => "0001000110001100000100",
			4633 => "0000000100100010110101",
			4634 => "0000001100100010110101",
			4635 => "0001000010111000000100",
			4636 => "0000000100100010110101",
			4637 => "0000000100100010110101",
			4638 => "0001010110000100010000",
			4639 => "0000011100110100001000",
			4640 => "0010010111100100000100",
			4641 => "0000000100100010110101",
			4642 => "1111111100100010110101",
			4643 => "0011000100010100000100",
			4644 => "0000001100100010110101",
			4645 => "0000000100100010110101",
			4646 => "0001000100001100001000",
			4647 => "0011101000111000000100",
			4648 => "0000000100100010110101",
			4649 => "0000000100100010110101",
			4650 => "0010001111001000000100",
			4651 => "0000010100100010110101",
			4652 => "0000000100100010110101",
			4653 => "0011000110000111001100",
			4654 => "0010100001010001100000",
			4655 => "0000101110101000101100",
			4656 => "0000101110101000100000",
			4657 => "0010100011101000010000",
			4658 => "0010111011000100001000",
			4659 => "0011110110100100000100",
			4660 => "0000001100101001101001",
			4661 => "1111111100101001101001",
			4662 => "0011110100010000000100",
			4663 => "1111111100101001101001",
			4664 => "0000000100101001101001",
			4665 => "0000100000110100001000",
			4666 => "0010000001010100000100",
			4667 => "0000001100101001101001",
			4668 => "0000000100101001101001",
			4669 => "0011110110100100000100",
			4670 => "0000001100101001101001",
			4671 => "0000000100101001101001",
			4672 => "0001011101100000000100",
			4673 => "0000000100101001101001",
			4674 => "0011010110000100000100",
			4675 => "0000010100101001101001",
			4676 => "0000001100101001101001",
			4677 => "0001010100011000011100",
			4678 => "0000101110010000010000",
			4679 => "0011101100001000001000",
			4680 => "0010010110101000000100",
			4681 => "0000000100101001101001",
			4682 => "0000000100101001101001",
			4683 => "0010001001101000000100",
			4684 => "0000000100101001101001",
			4685 => "0000000100101001101001",
			4686 => "0011001000111000001000",
			4687 => "0000000000111000000100",
			4688 => "0000000100101001101001",
			4689 => "0000000100101001101001",
			4690 => "0000001100101001101001",
			4691 => "0011100001101000001100",
			4692 => "0011001001110000001000",
			4693 => "0000111000011000000100",
			4694 => "0000001100101001101001",
			4695 => "0000010100101001101001",
			4696 => "0000000100101001101001",
			4697 => "0000010110101000000100",
			4698 => "1111111100101001101001",
			4699 => "0000000001110100000100",
			4700 => "0000001100101001101001",
			4701 => "0000000100101001101001",
			4702 => "0001001001001101000000",
			4703 => "0010011011101000100000",
			4704 => "0000101110010000010000",
			4705 => "0010010110101000001000",
			4706 => "0000001110111100000100",
			4707 => "0000001100101001101001",
			4708 => "0000000100101001101001",
			4709 => "0000000000111000000100",
			4710 => "0000001100101001101001",
			4711 => "0000000100101001101001",
			4712 => "0010111001110000001000",
			4713 => "0010011101101000000100",
			4714 => "0000001100101001101001",
			4715 => "0000000100101001101001",
			4716 => "0010001111001000000100",
			4717 => "0000000100101001101001",
			4718 => "0000001100101001101001",
			4719 => "0000101100010000010000",
			4720 => "0000000000111000001000",
			4721 => "0011010011100000000100",
			4722 => "0000001100101001101001",
			4723 => "0000000100101001101001",
			4724 => "0000111001001000000100",
			4725 => "1111111100101001101001",
			4726 => "0000000100101001101001",
			4727 => "0010110110000100001000",
			4728 => "0001010111001000000100",
			4729 => "0000000100101001101001",
			4730 => "0000001100101001101001",
			4731 => "0010101010110000000100",
			4732 => "0000001100101001101001",
			4733 => "0000000100101001101001",
			4734 => "0000110011111100001100",
			4735 => "0000000011011100000100",
			4736 => "1111111100101001101001",
			4737 => "0001000011111000000100",
			4738 => "0000000100101001101001",
			4739 => "1111111100101001101001",
			4740 => "0011110100000100010000",
			4741 => "0000111000111100001000",
			4742 => "0010011001111000000100",
			4743 => "0000000100101001101001",
			4744 => "1111111100101001101001",
			4745 => "0000011100110100000100",
			4746 => "0000011100101001101001",
			4747 => "0000010100101001101001",
			4748 => "0011001110111100001000",
			4749 => "0011001010000000000100",
			4750 => "0000000100101001101001",
			4751 => "0000001100101001101001",
			4752 => "0000111100001000000100",
			4753 => "1111111100101001101001",
			4754 => "0000000100101001101001",
			4755 => "0011001010111100001100",
			4756 => "0000000111000100001000",
			4757 => "0000001111001000000100",
			4758 => "1111111100101001101001",
			4759 => "0000001100101001101001",
			4760 => "1111111100101001101001",
			4761 => "1111111100101001101001",
			4762 => "0011110010001010000100",
			4763 => "0000110110000101011000",
			4764 => "0011011101111000110100",
			4765 => "0001011110001100100000",
			4766 => "0010110100000000010000",
			4767 => "0000011100110100001000",
			4768 => "0001011100101100000100",
			4769 => "0000000100110011000101",
			4770 => "0000000100110011000101",
			4771 => "0010010111100100000100",
			4772 => "0000000100110011000101",
			4773 => "1111111100110011000101",
			4774 => "0001000101000000001000",
			4775 => "0000011110100000000100",
			4776 => "1111111100110011000101",
			4777 => "0000001100110011000101",
			4778 => "0000011110100000000100",
			4779 => "0000000100110011000101",
			4780 => "1111111100110011000101",
			4781 => "0001001000000100000100",
			4782 => "1111111100110011000101",
			4783 => "0001001010110100001000",
			4784 => "0001000011001100000100",
			4785 => "0000000100110011000101",
			4786 => "0000001100110011000101",
			4787 => "0001001110111000000100",
			4788 => "1111111100110011000101",
			4789 => "0000000100110011000101",
			4790 => "0011111011011100011100",
			4791 => "0011011100101000010000",
			4792 => "0000111100110000001000",
			4793 => "0001111100001000000100",
			4794 => "0000000100110011000101",
			4795 => "1111111100110011000101",
			4796 => "0001101101111100000100",
			4797 => "0000000100110011000101",
			4798 => "0000001100110011000101",
			4799 => "0010111001110000000100",
			4800 => "1111111100110011000101",
			4801 => "0001100100110100000100",
			4802 => "0000000100110011000101",
			4803 => "0000000100110011000101",
			4804 => "0000011110100000000100",
			4805 => "0000000100110011000101",
			4806 => "1111111100110011000101",
			4807 => "0001111100001000010000",
			4808 => "0001110100010100000100",
			4809 => "1111111100110011000101",
			4810 => "0001100001111000000100",
			4811 => "0000000100110011000101",
			4812 => "0011101000111100000100",
			4813 => "0000001100110011000101",
			4814 => "0000001100110011000101",
			4815 => "0010010111100100001100",
			4816 => "0011110101100100000100",
			4817 => "1111111100110011000101",
			4818 => "0000111100101100000100",
			4819 => "0000001100110011000101",
			4820 => "0000001100110011000101",
			4821 => "0010111100001000000100",
			4822 => "1111111100110011000101",
			4823 => "0000110110000100000100",
			4824 => "0000001100110011000101",
			4825 => "0001101101111100000100",
			4826 => "0000000100110011000101",
			4827 => "1111111100110011000101",
			4828 => "0000111100101100110100",
			4829 => "0000111100101100101000",
			4830 => "0001011101111000100000",
			4831 => "0001011100101100010000",
			4832 => "0010110100000000001000",
			4833 => "0011011110001100000100",
			4834 => "0000000100110011000101",
			4835 => "1111111100110011000101",
			4836 => "0001111100001000000100",
			4837 => "0000000100110011000101",
			4838 => "0000001100110011000101",
			4839 => "0000011100110100001000",
			4840 => "0011100000101000000100",
			4841 => "1111111100110011000101",
			4842 => "0000000100110011000101",
			4843 => "0001110100000000000100",
			4844 => "0000001100110011000101",
			4845 => "1111111100110011000101",
			4846 => "0001110100000000000100",
			4847 => "0000001100110011000101",
			4848 => "0000000100110011000101",
			4849 => "0010010111100100001000",
			4850 => "0011010110000100000100",
			4851 => "0000000100110011000101",
			4852 => "1111111100110011000101",
			4853 => "0000000100110011000101",
			4854 => "0001000101010100111000",
			4855 => "0000011100110100100000",
			4856 => "0000000011111100010000",
			4857 => "0001100001111000001000",
			4858 => "0011011101111000000100",
			4859 => "0000001100110011000101",
			4860 => "0000000100110011000101",
			4861 => "0000111101111000000100",
			4862 => "0000000100110011000101",
			4863 => "0000000100110011000101",
			4864 => "0000011100110100001000",
			4865 => "0010110000101000000100",
			4866 => "0000001100110011000101",
			4867 => "0000000100110011000101",
			4868 => "0010111100001000000100",
			4869 => "0000000100110011000101",
			4870 => "0000001100110011000101",
			4871 => "0010110100000000001100",
			4872 => "0000111010111000001000",
			4873 => "0011011101111000000100",
			4874 => "0000000100110011000101",
			4875 => "1111111100110011000101",
			4876 => "0000001100110011000101",
			4877 => "0011011101111000000100",
			4878 => "0000001100110011000101",
			4879 => "0000001110111100000100",
			4880 => "0000000100110011000101",
			4881 => "1111111100110011000101",
			4882 => "0010000111000100100000",
			4883 => "0010111000111100010000",
			4884 => "0000011100110100001000",
			4885 => "0011010101101100000100",
			4886 => "0000001100110011000101",
			4887 => "1111111100110011000101",
			4888 => "0011011101111000000100",
			4889 => "0000001100110011000101",
			4890 => "0000000100110011000101",
			4891 => "0010100001010000001000",
			4892 => "0010001011010100000100",
			4893 => "0000000100110011000101",
			4894 => "0000001100110011000101",
			4895 => "0000000000110000000100",
			4896 => "1111111100110011000101",
			4897 => "0000000100110011000101",
			4898 => "0001000100001100010000",
			4899 => "0001101101011000001000",
			4900 => "0001111000111100000100",
			4901 => "0000000100110011000101",
			4902 => "0000000100110011000101",
			4903 => "0011111101000100000100",
			4904 => "1111111100110011000101",
			4905 => "0000000100110011000101",
			4906 => "0010100110011100001000",
			4907 => "0001010110000100000100",
			4908 => "0000000100110011000101",
			4909 => "1111111100110011000101",
			4910 => "0011110001001000000100",
			4911 => "0000001100110011000101",
			4912 => "0000000100110011000101",
			4913 => "0010100110011010101100",
			4914 => "0010001001101001011000",
			4915 => "0010001100000100110000",
			4916 => "0001001000011100010100",
			4917 => "0000000010011000010000",
			4918 => "0001001000110100001000",
			4919 => "0001001110000000000100",
			4920 => "0000000100111100101001",
			4921 => "0000000100111100101001",
			4922 => "0010111000111100000100",
			4923 => "0000001100111100101001",
			4924 => "0000000100111100101001",
			4925 => "1111111100111100101001",
			4926 => "0010101000010100010000",
			4927 => "0010101000100100001000",
			4928 => "0011100100000000000100",
			4929 => "0000000100111100101001",
			4930 => "0000000100111100101001",
			4931 => "0001000010110000000100",
			4932 => "1111111100111100101001",
			4933 => "0000000100111100101001",
			4934 => "0010101000010100001000",
			4935 => "0000001101010000000100",
			4936 => "0000000100111100101001",
			4937 => "0000001100111100101001",
			4938 => "1111111100111100101001",
			4939 => "0001000110111000001000",
			4940 => "0011011110110000000100",
			4941 => "1111111100111100101001",
			4942 => "0000000100111100101001",
			4943 => "0001000011110000010000",
			4944 => "0000000010111100001000",
			4945 => "0000000010111100000100",
			4946 => "0000000100111100101001",
			4947 => "0000000100111100101001",
			4948 => "0011100100010100000100",
			4949 => "0000000100111100101001",
			4950 => "0000001100111100101001",
			4951 => "0001111011000100001000",
			4952 => "0000111000111000000100",
			4953 => "0000000100111100101001",
			4954 => "0000001100111100101001",
			4955 => "0010111100001000000100",
			4956 => "0000000100111100101001",
			4957 => "1111111100111100101001",
			4958 => "0010101001000100100000",
			4959 => "0011000111111000001100",
			4960 => "0000000011111100000100",
			4961 => "1111111100111100101001",
			4962 => "0001010011011100000100",
			4963 => "0000000100111100101001",
			4964 => "0000001100111100101001",
			4965 => "0001111100001000010000",
			4966 => "0010010110101000001000",
			4967 => "0010011001111000000100",
			4968 => "1111111100111100101001",
			4969 => "0000000100111100101001",
			4970 => "0011000100010100000100",
			4971 => "1111111100111100101001",
			4972 => "1111111100111100101001",
			4973 => "0000000100111100101001",
			4974 => "0011010000001100011000",
			4975 => "0000000011010000001100",
			4976 => "0001001000110100000100",
			4977 => "1111111100111100101001",
			4978 => "0001000101000000000100",
			4979 => "0000001100111100101001",
			4980 => "0000000100111100101001",
			4981 => "0001001000001000000100",
			4982 => "1111111100111100101001",
			4983 => "0011000100010100000100",
			4984 => "0000000100111100101001",
			4985 => "0000001100111100101001",
			4986 => "0001010000001100001100",
			4987 => "0001111011000100000100",
			4988 => "0000000100111100101001",
			4989 => "0001111100001000000100",
			4990 => "1111110100111100101001",
			4991 => "1111111100111100101001",
			4992 => "0001011101010100001000",
			4993 => "0000010010001100000100",
			4994 => "0000000100111100101001",
			4995 => "0000001100111100101001",
			4996 => "0001000011110000000100",
			4997 => "0000000100111100101001",
			4998 => "1111111100111100101001",
			4999 => "0001001000001001001100",
			5000 => "0000000010111100011000",
			5001 => "0000100100101000000100",
			5002 => "1111111100111100101001",
			5003 => "0001000011110000010000",
			5004 => "0001001110100100001000",
			5005 => "0000111001110100000100",
			5006 => "1111111100111100101001",
			5007 => "0000000100111100101001",
			5008 => "0010010000111100000100",
			5009 => "0000001100111100101001",
			5010 => "1111111100111100101001",
			5011 => "1111111100111100101001",
			5012 => "0000000000111000011100",
			5013 => "0011011010111000010000",
			5014 => "0010100001010000001000",
			5015 => "0001000010110000000100",
			5016 => "0000001100111100101001",
			5017 => "0000000100111100101001",
			5018 => "0001000110001100000100",
			5019 => "0000001100111100101001",
			5020 => "0000001100111100101001",
			5021 => "0001011101010100000100",
			5022 => "1111111100111100101001",
			5023 => "0011001000111100000100",
			5024 => "0000001100111100101001",
			5025 => "0000000100111100101001",
			5026 => "0000100100101000001000",
			5027 => "0010100001010000000100",
			5028 => "1111111100111100101001",
			5029 => "0000000100111100101001",
			5030 => "0001111000111000001000",
			5031 => "0010001111001000000100",
			5032 => "0000001100111100101001",
			5033 => "0000000100111100101001",
			5034 => "0000000000111000000100",
			5035 => "0000000100111100101001",
			5036 => "1111111100111100101001",
			5037 => "0000000011111100001000",
			5038 => "0010001011010100000100",
			5039 => "1111111100111100101001",
			5040 => "1111111100111100101001",
			5041 => "0010111100101100100000",
			5042 => "0010011101101000010000",
			5043 => "0010110011011100001000",
			5044 => "0011100110000100000100",
			5045 => "0000000100111100101001",
			5046 => "0000000100111100101001",
			5047 => "0000110111001000000100",
			5048 => "0000001100111100101001",
			5049 => "0000000100111100101001",
			5050 => "0011101100101100001000",
			5051 => "0000000000110000000100",
			5052 => "0000000100111100101001",
			5053 => "1111111100111100101001",
			5054 => "0011000000101000000100",
			5055 => "0000000100111100101001",
			5056 => "0000000100111100101001",
			5057 => "0000101000001100010000",
			5058 => "0011000011011100001000",
			5059 => "0011100111001000000100",
			5060 => "0000010100111100101001",
			5061 => "0000001100111100101001",
			5062 => "0010011001011000000100",
			5063 => "0000000100111100101001",
			5064 => "0000001100111100101001",
			5065 => "1111111100111100101001",
			5066 => "0010011101101011000100",
			5067 => "0001111100001001011000",
			5068 => "0001111100001001000000",
			5069 => "0001110000101000100000",
			5070 => "0001110000101000010000",
			5071 => "0001110000101000001000",
			5072 => "0011000000101000000100",
			5073 => "0000000101000101100101",
			5074 => "0000001101000101100101",
			5075 => "0010001010101100000100",
			5076 => "0000000101000101100101",
			5077 => "0000001101000101100101",
			5078 => "0010010110101000001000",
			5079 => "0010110000101000000100",
			5080 => "1111111101000101100101",
			5081 => "0000000101000101100101",
			5082 => "0011101110111100000100",
			5083 => "0000000101000101100101",
			5084 => "1111111101000101100101",
			5085 => "0010010111100100010000",
			5086 => "0000011100110100001000",
			5087 => "0010110000101000000100",
			5088 => "0000001101000101100101",
			5089 => "0000000101000101100101",
			5090 => "0000101001010000000100",
			5091 => "0000001101000101100101",
			5092 => "0000000101000101100101",
			5093 => "0001111100001000001000",
			5094 => "0010001001101000000100",
			5095 => "0000000101000101100101",
			5096 => "0000000101000101100101",
			5097 => "0000000011010000000100",
			5098 => "0000000101000101100101",
			5099 => "0000000101000101100101",
			5100 => "0000010010001100010100",
			5101 => "0011111101000100010000",
			5102 => "0001101100011000001000",
			5103 => "0011000100010100000100",
			5104 => "1111111101000101100101",
			5105 => "0000000101000101100101",
			5106 => "0011000100010100000100",
			5107 => "0000010101000101100101",
			5108 => "0000000101000101100101",
			5109 => "1111111101000101100101",
			5110 => "1111110101000101100101",
			5111 => "0011101000111000110000",
			5112 => "0010110100000000011000",
			5113 => "0001110100000000010000",
			5114 => "0011101010000000001000",
			5115 => "0000101100100100000100",
			5116 => "0000001101000101100101",
			5117 => "1111111101000101100101",
			5118 => "0011110101110100000100",
			5119 => "0000001101000101100101",
			5120 => "0000000101000101100101",
			5121 => "0001101100011000000100",
			5122 => "1111111101000101100101",
			5123 => "0000000101000101100101",
			5124 => "0000111100110000001000",
			5125 => "0010001001101000000100",
			5126 => "0000000101000101100101",
			5127 => "1111111101000101100101",
			5128 => "0011110001011000001000",
			5129 => "0000110110000100000100",
			5130 => "0000001101000101100101",
			5131 => "0000000101000101100101",
			5132 => "0010010111100100000100",
			5133 => "0000000101000101100101",
			5134 => "1111111101000101100101",
			5135 => "0010010111100100100000",
			5136 => "0010000111000100010000",
			5137 => "0001110100000000001000",
			5138 => "0011100011011100000100",
			5139 => "0000001101000101100101",
			5140 => "0000000101000101100101",
			5141 => "0001110100000000000100",
			5142 => "1111111101000101100101",
			5143 => "0000001101000101100101",
			5144 => "0001000100001100001000",
			5145 => "0011000000101000000100",
			5146 => "0000001101000101100101",
			5147 => "0000010101000101100101",
			5148 => "0000111010111100000100",
			5149 => "0000000101000101100101",
			5150 => "0000001101000101100101",
			5151 => "0011000100010100010000",
			5152 => "0001101100011000001000",
			5153 => "0011110101110100000100",
			5154 => "0000010101000101100101",
			5155 => "0000000101000101100101",
			5156 => "0011111110101100000100",
			5157 => "0000000101000101100101",
			5158 => "0000010101000101100101",
			5159 => "0011001011000100000100",
			5160 => "1111111101000101100101",
			5161 => "0000011100110100000100",
			5162 => "0000000101000101100101",
			5163 => "0000000101000101100101",
			5164 => "0011110110110100010000",
			5165 => "0010001010110000001100",
			5166 => "0000111000000000000100",
			5167 => "1111111101000101100101",
			5168 => "0011100111001000000100",
			5169 => "0000000101000101100101",
			5170 => "0000000101000101100101",
			5171 => "0000010101000101100101",
			5172 => "0000110001111100010100",
			5173 => "0000010010001100000100",
			5174 => "0000000101000101100101",
			5175 => "0000101001010000000100",
			5176 => "0000000101000101100101",
			5177 => "0001001000001000000100",
			5178 => "1111110101000101100101",
			5179 => "0001111000111000000100",
			5180 => "1111111101000101100101",
			5181 => "1111111101000101100101",
			5182 => "0011000100010100011000",
			5183 => "0011000100010100001000",
			5184 => "0000100110010000000100",
			5185 => "0000001101000101100101",
			5186 => "0000000101000101100101",
			5187 => "0001110100000000001000",
			5188 => "0001111100001000000100",
			5189 => "1111111101000101100101",
			5190 => "0000001101000101100101",
			5191 => "0010110011011100000100",
			5192 => "1111111101000101100101",
			5193 => "0000000101000101100101",
			5194 => "0001110100000000010000",
			5195 => "0011101100101000001000",
			5196 => "0000111010111000000100",
			5197 => "0000000101000101100101",
			5198 => "1111111101000101100101",
			5199 => "0001101100011000000100",
			5200 => "0000000101000101100101",
			5201 => "0000001101000101100101",
			5202 => "0001101101111100001000",
			5203 => "0000101001010000000100",
			5204 => "0000000101000101100101",
			5205 => "1111111101000101100101",
			5206 => "0001000011110000000100",
			5207 => "0000000101000101100101",
			5208 => "0000000101000101100101",
			5209 => "0011000110000111010000",
			5210 => "0010100001010001101100",
			5211 => "0000101110101000110000",
			5212 => "0000101101000100011100",
			5213 => "0010100011101000001100",
			5214 => "0010110100010100000100",
			5215 => "0000001101001100100001",
			5216 => "0001100111101000000100",
			5217 => "1111111101001100100001",
			5218 => "0000000101001100100001",
			5219 => "0000100000110100001000",
			5220 => "0010000001010100000100",
			5221 => "0000001101001100100001",
			5222 => "1111111101001100100001",
			5223 => "0001001001001100000100",
			5224 => "0000000101001100100001",
			5225 => "0000001101001100100001",
			5226 => "0011000000101000010000",
			5227 => "0010001011010100001000",
			5228 => "0001001000001000000100",
			5229 => "0000001101001100100001",
			5230 => "0000011101001100100001",
			5231 => "0001000101010100000100",
			5232 => "0000000101001100100001",
			5233 => "0000010101001100100001",
			5234 => "0000000101001100100001",
			5235 => "0001101100011000100000",
			5236 => "0000100011001000010000",
			5237 => "0010100001010000001000",
			5238 => "0001101101111100000100",
			5239 => "0000000101001100100001",
			5240 => "0000000101001100100001",
			5241 => "0011000100010100000100",
			5242 => "1111111101001100100001",
			5243 => "0000000101001100100001",
			5244 => "0000011100110100001000",
			5245 => "0000011100110100000100",
			5246 => "0000000101001100100001",
			5247 => "0000000101001100100001",
			5248 => "0000100011001000000100",
			5249 => "0000000101001100100001",
			5250 => "1111111101001100100001",
			5251 => "0010011101101000001100",
			5252 => "0010001111001000001000",
			5253 => "0001000101010100000100",
			5254 => "0000001101001100100001",
			5255 => "0000000101001100100001",
			5256 => "0000000101001100100001",
			5257 => "0001001010110100001000",
			5258 => "0000001111000100000100",
			5259 => "0000000101001100100001",
			5260 => "0000000101001100100001",
			5261 => "0010111100101100000100",
			5262 => "1111111101001100100001",
			5263 => "0000001101001100100001",
			5264 => "0001001001001101000000",
			5265 => "0010011011101000100000",
			5266 => "0000101110010000010000",
			5267 => "0010010111100100001000",
			5268 => "0010000111000100000100",
			5269 => "0000001101001100100001",
			5270 => "0000000101001100100001",
			5271 => "0000000000110000000100",
			5272 => "0000001101001100100001",
			5273 => "1111111101001100100001",
			5274 => "0011000000101000001000",
			5275 => "0011000000101000000100",
			5276 => "0000001101001100100001",
			5277 => "0000000101001100100001",
			5278 => "0001011100101000000100",
			5279 => "0000001101001100100001",
			5280 => "0000001101001100100001",
			5281 => "0000101100000000010000",
			5282 => "0000000000111000001000",
			5283 => "0011010011100000000100",
			5284 => "0000001101001100100001",
			5285 => "0000000101001100100001",
			5286 => "0011101101010100000100",
			5287 => "1111111101001100100001",
			5288 => "0000000101001100100001",
			5289 => "0011100010001000001000",
			5290 => "0001000011001100000100",
			5291 => "0000011101001100100001",
			5292 => "0000001101001100100001",
			5293 => "0001110110000100000100",
			5294 => "1111111101001100100001",
			5295 => "0000001101001100100001",
			5296 => "0010101100000100100000",
			5297 => "0010001111001000010000",
			5298 => "0001111100001000001000",
			5299 => "0010011001111000000100",
			5300 => "1111111101001100100001",
			5301 => "0000001101001100100001",
			5302 => "0010001111001000000100",
			5303 => "0000000101001100100001",
			5304 => "1111111101001100100001",
			5305 => "0000001010000000001000",
			5306 => "0010000111000100000100",
			5307 => "1111111101001100100001",
			5308 => "0000000101001100100001",
			5309 => "0011101111000100000100",
			5310 => "0000000101001100100001",
			5311 => "0000000101001100100001",
			5312 => "1111111101001100100001",
			5313 => "0011001010111100001100",
			5314 => "0000000111000100001000",
			5315 => "0000001111001000000100",
			5316 => "1111111101001100100001",
			5317 => "0000001101001100100001",
			5318 => "1111111101001100100001",
			5319 => "1111111101001100100001",
			5320 => "0011110000110111010000",
			5321 => "0000111001110001101000",
			5322 => "0010011001111000110000",
			5323 => "0000011110100000011100",
			5324 => "0011010110000100010000",
			5325 => "0000111000111000001000",
			5326 => "0011110110110100000100",
			5327 => "0000000101010111001101",
			5328 => "0000000101010111001101",
			5329 => "0011000000110000000100",
			5330 => "1111111101010111001101",
			5331 => "0000001101010111001101",
			5332 => "0000010110000000001000",
			5333 => "0011100011111100000100",
			5334 => "1111111101010111001101",
			5335 => "0000001101010111001101",
			5336 => "1111111101010111001101",
			5337 => "0000100100101000001100",
			5338 => "0011101110111100001000",
			5339 => "0010000111000100000100",
			5340 => "0000000101010111001101",
			5341 => "0000001101010111001101",
			5342 => "0000001101010111001101",
			5343 => "0000110100000000000100",
			5344 => "0000000101010111001101",
			5345 => "1111111101010111001101",
			5346 => "0000011110100000011000",
			5347 => "0001110100010100001000",
			5348 => "0001011101100000000100",
			5349 => "1111111101010111001101",
			5350 => "0000001101010111001101",
			5351 => "0011000100010100001000",
			5352 => "0001101110010100000100",
			5353 => "0000000101010111001101",
			5354 => "1111111101010111001101",
			5355 => "0001110000101000000100",
			5356 => "0000000101010111001101",
			5357 => "1111111101010111001101",
			5358 => "0011000111111000010000",
			5359 => "0011000111111000001000",
			5360 => "0011110101100100000100",
			5361 => "0000000101010111001101",
			5362 => "1111111101010111001101",
			5363 => "0000111000111100000100",
			5364 => "0000000101010111001101",
			5365 => "1111111101010111001101",
			5366 => "0001010110000100001000",
			5367 => "0010000111000100000100",
			5368 => "0000001101010111001101",
			5369 => "0000000101010111001101",
			5370 => "0001111100001000000100",
			5371 => "1111111101010111001101",
			5372 => "0000000101010111001101",
			5373 => "0001110100010100101100",
			5374 => "0000011110100000011100",
			5375 => "0001001000001000001100",
			5376 => "0001001100001100001000",
			5377 => "0011001010000000000100",
			5378 => "0000001101010111001101",
			5379 => "0000000101010111001101",
			5380 => "1111111101010111001101",
			5381 => "0000101110010000001000",
			5382 => "0010101010110000000100",
			5383 => "0000000101010111001101",
			5384 => "0000001101010111001101",
			5385 => "0010000001110100000100",
			5386 => "1111111101010111001101",
			5387 => "0000000101010111001101",
			5388 => "0000100010011100001100",
			5389 => "0011011100101100000100",
			5390 => "0000000101010111001101",
			5391 => "0001011100101100000100",
			5392 => "0000001101010111001101",
			5393 => "0000000101010111001101",
			5394 => "0000001101010111001101",
			5395 => "0001111000111000100000",
			5396 => "0011000100000000010000",
			5397 => "0011000100000000001000",
			5398 => "0011000000101000000100",
			5399 => "0000000101010111001101",
			5400 => "0000000101010111001101",
			5401 => "0010101010110000000100",
			5402 => "1111111101010111001101",
			5403 => "0000000101010111001101",
			5404 => "0001010000001100001000",
			5405 => "0011010000001100000100",
			5406 => "0000001101010111001101",
			5407 => "0000001101010111001101",
			5408 => "0011101101100000000100",
			5409 => "0000000101010111001101",
			5410 => "0000001101010111001101",
			5411 => "0010001111001000010000",
			5412 => "0001011010111100001000",
			5413 => "0011100110000100000100",
			5414 => "0000000101010111001101",
			5415 => "0000001101010111001101",
			5416 => "0011000000101000000100",
			5417 => "1111111101010111001101",
			5418 => "0000000101010111001101",
			5419 => "0010011101101000001000",
			5420 => "0001011100101000000100",
			5421 => "1111111101010111001101",
			5422 => "0000000101010111001101",
			5423 => "1111111101010111001101",
			5424 => "0011100100001001010000",
			5425 => "0011111101000100110000",
			5426 => "0011110010110100011100",
			5427 => "0000101001011100001100",
			5428 => "0000100111111100001000",
			5429 => "0001100100110100000100",
			5430 => "0000000101010111001101",
			5431 => "0000000101010111001101",
			5432 => "1111111101010111001101",
			5433 => "0001111100001000001000",
			5434 => "0000111110001100000100",
			5435 => "0000000101010111001101",
			5436 => "0000000101010111001101",
			5437 => "0001110100000000000100",
			5438 => "0000000101010111001101",
			5439 => "0000000101010111001101",
			5440 => "0001111001110000010000",
			5441 => "0001101010011000001000",
			5442 => "0010011101101000000100",
			5443 => "0000000101010111001101",
			5444 => "1111111101010111001101",
			5445 => "0000100110010000000100",
			5446 => "0000000101010111001101",
			5447 => "0000000101010111001101",
			5448 => "1111111101010111001101",
			5449 => "0000100110010000000100",
			5450 => "0000001101010111001101",
			5451 => "0010011101101000001100",
			5452 => "0001001011100000001000",
			5453 => "0000010010001100000100",
			5454 => "0000000101010111001101",
			5455 => "0000001101010111001101",
			5456 => "1111111101010111001101",
			5457 => "0011000100000000001000",
			5458 => "0001000000010100000100",
			5459 => "1111111101010111001101",
			5460 => "0000000101010111001101",
			5461 => "0001111001110000000100",
			5462 => "0000000101010111001101",
			5463 => "1111111101010111001101",
			5464 => "0011100001111100011100",
			5465 => "0011000100000000010100",
			5466 => "0001011010111100010000",
			5467 => "0000111110110000001000",
			5468 => "0000110111001000000100",
			5469 => "0000000101010111001101",
			5470 => "1111111101010111001101",
			5471 => "0000100010000100000100",
			5472 => "0000001101010111001101",
			5473 => "0000000101010111001101",
			5474 => "1111111101010111001101",
			5475 => "0010011111001100000100",
			5476 => "0000001101010111001101",
			5477 => "0000000101010111001101",
			5478 => "0001110000101000000100",
			5479 => "0000001101010111001101",
			5480 => "0000011100110100001000",
			5481 => "0001001001001100000100",
			5482 => "0000000101010111001101",
			5483 => "1111111101010111001101",
			5484 => "0011111001011100001000",
			5485 => "0011111110101000000100",
			5486 => "0000000101010111001101",
			5487 => "0000000101010111001101",
			5488 => "0011110010000000000100",
			5489 => "0000000101010111001101",
			5490 => "0000000101010111001101",
			5491 => "0011000100001011010100",
			5492 => "0011111010010101011000",
			5493 => "0011010111001001000000",
			5494 => "0011100111111000100000",
			5495 => "0001111100001000010000",
			5496 => "0000011100110100001000",
			5497 => "0001010101101100000100",
			5498 => "0000000101011101111011",
			5499 => "0000000101011101111011",
			5500 => "0010111100001000000100",
			5501 => "0000010101011101111011",
			5502 => "0000000101011101111011",
			5503 => "0001010110000100001000",
			5504 => "0010100110011100000100",
			5505 => "1111111101011101111011",
			5506 => "0000000101011101111011",
			5507 => "0010010110101000000100",
			5508 => "0000001101011101111011",
			5509 => "1111111101011101111011",
			5510 => "0001001111100000010000",
			5511 => "0010010110101000001000",
			5512 => "0011010101101100000100",
			5513 => "0000000101011101111011",
			5514 => "0000001101011101111011",
			5515 => "0000011110100000000100",
			5516 => "1111111101011101111011",
			5517 => "0000000101011101111011",
			5518 => "0000101001011100001000",
			5519 => "0010100110011100000100",
			5520 => "0000010101011101111011",
			5521 => "1111111101011101111011",
			5522 => "0011110111110000000100",
			5523 => "0000000101011101111011",
			5524 => "0000001101011101111011",
			5525 => "0000010010001100001000",
			5526 => "0011010011100000000100",
			5527 => "1111110101011101111011",
			5528 => "1111111101011101111011",
			5529 => "0001001000001000001100",
			5530 => "0010101000010100001000",
			5531 => "0001001000101000000100",
			5532 => "0000000101011101111011",
			5533 => "1111111101011101111011",
			5534 => "0000001101011101111011",
			5535 => "1111111101011101111011",
			5536 => "0001101100011000111100",
			5537 => "0011101101100000100000",
			5538 => "0010010110101000010000",
			5539 => "0010100110011000001000",
			5540 => "0011101001110000000100",
			5541 => "1111111101011101111011",
			5542 => "0000000101011101111011",
			5543 => "0000101100010100000100",
			5544 => "0000000101011101111011",
			5545 => "0000000101011101111011",
			5546 => "0000011100110100001000",
			5547 => "0000101110010000000100",
			5548 => "1111110101011101111011",
			5549 => "1111111101011101111011",
			5550 => "0010011101101000000100",
			5551 => "0000000101011101111011",
			5552 => "1111111101011101111011",
			5553 => "0000100110010000010000",
			5554 => "0011010000001100001000",
			5555 => "0011001010000000000100",
			5556 => "1111101101011101111011",
			5557 => "0000000101011101111011",
			5558 => "0001101100011000000100",
			5559 => "0000000101011101111011",
			5560 => "1111111101011101111011",
			5561 => "0011000100010100000100",
			5562 => "0000000101011101111011",
			5563 => "0000000010111100000100",
			5564 => "0000000101011101111011",
			5565 => "1111111101011101111011",
			5566 => "0010011101101000100000",
			5567 => "0001001111100000010000",
			5568 => "0010101100011100001000",
			5569 => "0011011101010100000100",
			5570 => "0000000101011101111011",
			5571 => "0000001101011101111011",
			5572 => "0010111000111100000100",
			5573 => "0000000101011101111011",
			5574 => "0000001101011101111011",
			5575 => "0010010110101000001000",
			5576 => "0000101001100000000100",
			5577 => "0000000101011101111011",
			5578 => "0000001101011101111011",
			5579 => "0001101101011000000100",
			5580 => "1111111101011101111011",
			5581 => "0000000101011101111011",
			5582 => "0000100111011000010000",
			5583 => "0000001110111100001000",
			5584 => "0011000100010100000100",
			5585 => "0000000101011101111011",
			5586 => "0000000101011101111011",
			5587 => "0010111000111000000100",
			5588 => "0000000101011101111011",
			5589 => "0000000101011101111011",
			5590 => "0000100111011000001000",
			5591 => "0011100100011000000100",
			5592 => "0000010101011101111011",
			5593 => "0000001101011101111011",
			5594 => "0001001011100000000100",
			5595 => "0000000101011101111011",
			5596 => "1111111101011101111011",
			5597 => "1111111101011101111011",
			5598 => "0001111101111001110100",
			5599 => "0001000001001101101000",
			5600 => "0000000100010100110000",
			5601 => "0001100001000100010000",
			5602 => "0000110000111000000100",
			5603 => "0000001101100010000101",
			5604 => "0000110111111000001000",
			5605 => "0000111110111100000100",
			5606 => "1111111101100010000101",
			5607 => "0000000101100010000101",
			5608 => "1111111101100010000101",
			5609 => "0001111100001000010000",
			5610 => "0000111101100000001000",
			5611 => "0001110111111000000100",
			5612 => "0000001101100010000101",
			5613 => "0000000101100010000101",
			5614 => "0000100100101000000100",
			5615 => "0000001101100010000101",
			5616 => "0000000101100010000101",
			5617 => "0001111100001000001000",
			5618 => "0011011100101000000100",
			5619 => "0000000101100010000101",
			5620 => "1111111101100010000101",
			5621 => "0001100001111000000100",
			5622 => "1111111101100010000101",
			5623 => "0000000101100010000101",
			5624 => "0001101010011000100000",
			5625 => "0010100110011100010000",
			5626 => "0001011000111100001000",
			5627 => "0000100001000000000100",
			5628 => "0000000101100010000101",
			5629 => "0000001101100010000101",
			5630 => "0011110101100100000100",
			5631 => "0000000101100010000101",
			5632 => "0000000101100010000101",
			5633 => "0001000001101100001000",
			5634 => "0010000111000000000100",
			5635 => "0000001101100010000101",
			5636 => "1111111101100010000101",
			5637 => "0001101100011000000100",
			5638 => "0000010101100010000101",
			5639 => "0000000101100010000101",
			5640 => "0000101100010000001100",
			5641 => "0010000010101000000100",
			5642 => "0000000101100010000101",
			5643 => "0011011110110000000100",
			5644 => "1111111101100010000101",
			5645 => "0000000101100010000101",
			5646 => "0010111101100000001000",
			5647 => "0000010010001100000100",
			5648 => "0000000101100010000101",
			5649 => "0000010101100010000101",
			5650 => "1111111101100010000101",
			5651 => "0001001011100100001000",
			5652 => "0001101011111100000100",
			5653 => "1111111101100010000101",
			5654 => "0000000101100010000101",
			5655 => "1111111101100010000101",
			5656 => "0010100111110100010000",
			5657 => "0000101100111000001100",
			5658 => "0001111100101000001000",
			5659 => "0010000000001000000100",
			5660 => "1111111101100010000101",
			5661 => "0000001101100010000101",
			5662 => "1111111101100010000101",
			5663 => "0000011101100010000101",
			5664 => "1111111101100010000101",
			5665 => "0000101110101001010100",
			5666 => "0000011001111001001100",
			5667 => "0011101000111100111000",
			5668 => "0001011110001100100000",
			5669 => "0011100000110000010000",
			5670 => "0011010101101100001000",
			5671 => "0011111010001100000100",
			5672 => "0000000101101000000001",
			5673 => "1111111101101000000001",
			5674 => "0000111000111100000100",
			5675 => "0000000101101000000001",
			5676 => "1111111101101000000001",
			5677 => "0010001001101000001000",
			5678 => "0001100001111000000100",
			5679 => "0000000101101000000001",
			5680 => "1111111101101000000001",
			5681 => "0001110000101000000100",
			5682 => "0000001101101000000001",
			5683 => "0000001101101000000001",
			5684 => "0011111111011100001100",
			5685 => "0001001010110100001000",
			5686 => "0000100000110100000100",
			5687 => "1111111101101000000001",
			5688 => "0000001101101000000001",
			5689 => "1111111101101000000001",
			5690 => "0001011110001100000100",
			5691 => "1111111101101000000001",
			5692 => "0011011101111000000100",
			5693 => "0000000101101000000001",
			5694 => "1111111101101000000001",
			5695 => "0010100011101000001100",
			5696 => "0001000110111100001000",
			5697 => "0000011100110100000100",
			5698 => "0000000101101000000001",
			5699 => "0000000101101000000001",
			5700 => "1111111101101000000001",
			5701 => "0011110010001000000100",
			5702 => "0000001101101000000001",
			5703 => "0000000101101000000001",
			5704 => "0011111001010100000100",
			5705 => "1111111101101000000001",
			5706 => "0000000101101000000001",
			5707 => "0000101110101000010100",
			5708 => "0001110000101000001100",
			5709 => "0011100000110000001000",
			5710 => "0001111110111100000100",
			5711 => "0000001101101000000001",
			5712 => "1111111101101000000001",
			5713 => "0000000101101000000001",
			5714 => "0001010011100000000100",
			5715 => "1111111101101000000001",
			5716 => "0000000101101000000001",
			5717 => "0000110100010100101000",
			5718 => "0001001011100000001100",
			5719 => "0001100001111000001000",
			5720 => "0000010110000000000100",
			5721 => "0000001101101000000001",
			5722 => "1111111101101000000001",
			5723 => "1111111101101000000001",
			5724 => "0001110100010100010000",
			5725 => "0000100101110000001000",
			5726 => "0000111110111100000100",
			5727 => "0000000101101000000001",
			5728 => "0000001101101000000001",
			5729 => "0011111111011100000100",
			5730 => "0000000101101000000001",
			5731 => "1111111101101000000001",
			5732 => "0000100101110000000100",
			5733 => "1111111101101000000001",
			5734 => "0011100111000000000100",
			5735 => "0000000101101000000001",
			5736 => "0000000101101000000001",
			5737 => "0011010011011100010100",
			5738 => "0001110100010100010000",
			5739 => "0011110100010000001000",
			5740 => "0001001010110100000100",
			5741 => "0000000101101000000001",
			5742 => "0000001101101000000001",
			5743 => "0000100011001000000100",
			5744 => "1111111101101000000001",
			5745 => "0000000101101000000001",
			5746 => "1111111101101000000001",
			5747 => "0011111010011100001100",
			5748 => "0011111010011100001000",
			5749 => "0011010110000100000100",
			5750 => "1111111101101000000001",
			5751 => "0000001101101000000001",
			5752 => "0000001101101000000001",
			5753 => "0000110011011100001000",
			5754 => "0011110110110100000100",
			5755 => "0000000101101000000001",
			5756 => "0000000101101000000001",
			5757 => "0010010110101000000100",
			5758 => "0000000101101000000001",
			5759 => "0000000101101000000001",
			5760 => "0011000011011101101000",
			5761 => "0001000011111001100100",
			5762 => "0001111001110001000000",
			5763 => "0011101000111000100000",
			5764 => "0011110010001000010000",
			5765 => "0011010000001100001000",
			5766 => "0000111101100000000100",
			5767 => "0000000101101100100101",
			5768 => "0000001101101100100101",
			5769 => "0000010010001100000100",
			5770 => "1111111101101100100101",
			5771 => "0000001101101100100101",
			5772 => "0010101001000100001000",
			5773 => "0001011101111000000100",
			5774 => "1111111101101100100101",
			5775 => "0000000101101100100101",
			5776 => "0000000011111100000100",
			5777 => "0000001101101100100101",
			5778 => "0000000101101100100101",
			5779 => "0010011101101000010000",
			5780 => "0001111100001000001000",
			5781 => "0001111100001000000100",
			5782 => "0000000101101100100101",
			5783 => "0000000101101100100101",
			5784 => "0001001111100000000100",
			5785 => "0000001101101100100101",
			5786 => "0000000101101100100101",
			5787 => "0011100110000100001000",
			5788 => "0000010010001100000100",
			5789 => "1111111101101100100101",
			5790 => "0000000101101100100101",
			5791 => "0001001101001000000100",
			5792 => "0000000101101100100101",
			5793 => "0000000101101100100101",
			5794 => "0001011100101000000100",
			5795 => "0000001101101100100101",
			5796 => "0000110100011000010000",
			5797 => "0001010111001000001000",
			5798 => "0011111110101100000100",
			5799 => "1111111101101100100101",
			5800 => "0000000101101100100101",
			5801 => "0000110111001000000100",
			5802 => "0000001101101100100101",
			5803 => "1111111101101100100101",
			5804 => "0001101011001100001000",
			5805 => "0011111001010000000100",
			5806 => "0000000101101100100101",
			5807 => "0000001101101100100101",
			5808 => "0010100110011000000100",
			5809 => "0000001101101100100101",
			5810 => "1111111101101100100101",
			5811 => "1111111101101100100101",
			5812 => "0011000110000100011000",
			5813 => "0010111000000000010100",
			5814 => "0010011101011100000100",
			5815 => "1111111101101100100101",
			5816 => "0010011101011100000100",
			5817 => "0000001101101100100101",
			5818 => "0010111010111100001000",
			5819 => "0011010111010000000100",
			5820 => "0000000101101100100101",
			5821 => "0000001101101100100101",
			5822 => "1111111101101100100101",
			5823 => "0000001101101100100101",
			5824 => "0011001010111100010000",
			5825 => "0010100111110100001100",
			5826 => "0010100111110100000100",
			5827 => "1111111101101100100101",
			5828 => "0011000000001100000100",
			5829 => "0000000101101100100101",
			5830 => "0000001101101100100101",
			5831 => "1111111101101100100101",
			5832 => "1111111101101100100101",
			5833 => "0011101000000010001100",
			5834 => "0010011111001101010100",
			5835 => "0010110101101101000000",
			5836 => "0000011110100000100000",
			5837 => "0010010010001100010000",
			5838 => "0000111100001000001000",
			5839 => "0011110001011000000100",
			5840 => "0000000101110011101001",
			5841 => "0000000101110011101001",
			5842 => "0001011100110000000100",
			5843 => "0000001101110011101001",
			5844 => "1111111101110011101001",
			5845 => "0001011100110000001000",
			5846 => "0010101010110000000100",
			5847 => "1111111101110011101001",
			5848 => "0000000101110011101001",
			5849 => "0011100000110000000100",
			5850 => "0000000101110011101001",
			5851 => "0000001101110011101001",
			5852 => "0011111111011100010000",
			5853 => "0011111010011100001000",
			5854 => "0010111011000100000100",
			5855 => "0000001101110011101001",
			5856 => "0000000101110011101001",
			5857 => "0010110000101000000100",
			5858 => "0000000101110011101001",
			5859 => "0000001101110011101001",
			5860 => "0001010011011100001000",
			5861 => "0011000111111000000100",
			5862 => "0000000101110011101001",
			5863 => "0000001101110011101001",
			5864 => "0010111011000100000100",
			5865 => "0000000101110011101001",
			5866 => "0000000101110011101001",
			5867 => "0001011110110000001100",
			5868 => "0001010111001000000100",
			5869 => "0000000101110011101001",
			5870 => "0000110011100000000100",
			5871 => "0000000101110011101001",
			5872 => "0000010101110011101001",
			5873 => "0010011111001100000100",
			5874 => "1111111101110011101001",
			5875 => "0000001101110011101001",
			5876 => "0000000000110000100000",
			5877 => "0000011001111000000100",
			5878 => "1111111101110011101001",
			5879 => "0001111000111000001100",
			5880 => "0010100110011000001000",
			5881 => "0000111001001000000100",
			5882 => "1111111101110011101001",
			5883 => "0000000101110011101001",
			5884 => "0000000101110011101001",
			5885 => "0010011101011100001000",
			5886 => "0011001001110000000100",
			5887 => "0000001101110011101001",
			5888 => "1111111101110011101001",
			5889 => "0010100001010000000100",
			5890 => "0000000101110011101001",
			5891 => "1111111101110011101001",
			5892 => "0010011001011000010000",
			5893 => "0001101001100100000100",
			5894 => "1111111101110011101001",
			5895 => "0001010100011000000100",
			5896 => "1111111101110011101001",
			5897 => "0000011001111000000100",
			5898 => "0000001101110011101001",
			5899 => "0000000101110011101001",
			5900 => "0010110000001100000100",
			5901 => "0000001101110011101001",
			5902 => "0000000101110011101001",
			5903 => "0001101001100101000100",
			5904 => "0010101100011100110000",
			5905 => "0011000100000000011000",
			5906 => "0001101011001100001100",
			5907 => "0000110110100100000100",
			5908 => "0000000101110011101001",
			5909 => "0011000000101000000100",
			5910 => "0000000101110011101001",
			5911 => "0000001101110011101001",
			5912 => "0000010111100100001000",
			5913 => "0000000011111100000100",
			5914 => "0000000101110011101001",
			5915 => "1111111101110011101001",
			5916 => "0000001101110011101001",
			5917 => "0000011001111000001000",
			5918 => "0000011001111000000100",
			5919 => "0000000101110011101001",
			5920 => "1111111101110011101001",
			5921 => "0001101001100100001000",
			5922 => "0011101010001100000100",
			5923 => "0000000101110011101001",
			5924 => "0000000101110011101001",
			5925 => "0001011000000000000100",
			5926 => "0000000101110011101001",
			5927 => "0000001101110011101001",
			5928 => "0011110100101000001000",
			5929 => "0011000100000000000100",
			5930 => "0000001101110011101001",
			5931 => "1111111101110011101001",
			5932 => "0011110010000000001000",
			5933 => "0011000011011100000100",
			5934 => "0000001101110011101001",
			5935 => "0000000101110011101001",
			5936 => "1111111101110011101001",
			5937 => "0000010110101000001000",
			5938 => "0010110110000100000100",
			5939 => "0000001101110011101001",
			5940 => "1111111101110011101001",
			5941 => "0001100100111100000100",
			5942 => "1111111101110011101001",
			5943 => "0011110010000000000100",
			5944 => "0000001101110011101001",
			5945 => "1111111101110011101001",
			5946 => "0001111101100010011000",
			5947 => "0000101110101001001000",
			5948 => "0000010110000000011100",
			5949 => "0001010011011100011000",
			5950 => "0001011001110000001100",
			5951 => "0001011000111000001000",
			5952 => "0000110011111100000100",
			5953 => "0000000101111010010101",
			5954 => "0000001101111010010101",
			5955 => "1111111101111010010101",
			5956 => "0000110000111000000100",
			5957 => "1111111101111010010101",
			5958 => "0000000000111000000100",
			5959 => "0000000101111010010101",
			5960 => "0000010101111010010101",
			5961 => "1111111101111010010101",
			5962 => "0010010010001100010000",
			5963 => "0001110100010100001000",
			5964 => "0000111110111100000100",
			5965 => "0000000101111010010101",
			5966 => "0000010101111010010101",
			5967 => "0001010011011100000100",
			5968 => "0000010101111010010101",
			5969 => "0000011101111010010101",
			5970 => "0001100111101000010000",
			5971 => "0011100000110000001000",
			5972 => "0001000110111000000100",
			5973 => "0000001101111010010101",
			5974 => "1111111101111010010101",
			5975 => "0010100111110100000100",
			5976 => "0000000101111010010101",
			5977 => "0000001101111010010101",
			5978 => "0000111110111100000100",
			5979 => "1111111101111010010101",
			5980 => "0001110000101000000100",
			5981 => "0000001101111010010101",
			5982 => "0000000101111010010101",
			5983 => "0011111001011100111000",
			5984 => "0010011101011100100000",
			5985 => "0010101000010100010000",
			5986 => "0001001110000000001000",
			5987 => "0000101001010000000100",
			5988 => "0000000101111010010101",
			5989 => "0000000101111010010101",
			5990 => "0010111100001000000100",
			5991 => "0000000101111010010101",
			5992 => "1111111101111010010101",
			5993 => "0001001110100100001000",
			5994 => "0000001111000100000100",
			5995 => "0000000101111010010101",
			5996 => "0000001101111010010101",
			5997 => "0010100110011000000100",
			5998 => "0000000101111010010101",
			5999 => "0000000101111010010101",
			6000 => "0000000011111100001100",
			6001 => "0011111110101100000100",
			6002 => "1111111101111010010101",
			6003 => "0001101101011000000100",
			6004 => "0000001101111010010101",
			6005 => "0000000101111010010101",
			6006 => "0010100001010000000100",
			6007 => "1111110101111010010101",
			6008 => "0011101011000000000100",
			6009 => "1111111101111010010101",
			6010 => "0000000101111010010101",
			6011 => "0000111001010100010100",
			6012 => "0010011011111100010000",
			6013 => "0010000111000100001000",
			6014 => "0001000010110000000100",
			6015 => "0000001101111010010101",
			6016 => "1111111101111010010101",
			6017 => "0001000100001100000100",
			6018 => "0000010101111010010101",
			6019 => "0000000101111010010101",
			6020 => "0000011101111010010101",
			6021 => "1111111101111010010101",
			6022 => "0000111010011100010000",
			6023 => "0011110010011100001100",
			6024 => "0010111100101100000100",
			6025 => "1111111101111010010101",
			6026 => "0010111100101100000100",
			6027 => "0000000101111010010101",
			6028 => "1111111101111010010101",
			6029 => "0000001101111010010101",
			6030 => "0010010101011100011000",
			6031 => "0000011001111000000100",
			6032 => "1111111101111010010101",
			6033 => "0000100010000100001000",
			6034 => "0000100110010000000100",
			6035 => "0000001101111010010101",
			6036 => "1111111101111010010101",
			6037 => "0011111110010000001000",
			6038 => "0001101001100100000100",
			6039 => "0000010101111010010101",
			6040 => "0000000101111010010101",
			6041 => "1111111101111010010101",
			6042 => "0001110110100100010100",
			6043 => "0001010001000000010000",
			6044 => "0010110100001000001000",
			6045 => "0001001100111000000100",
			6046 => "0000000101111010010101",
			6047 => "1111111101111010010101",
			6048 => "0001110110000100000100",
			6049 => "0000001101111010010101",
			6050 => "0000000101111010010101",
			6051 => "0000001101111010010101",
			6052 => "1111111101111010010101",
			6053 => "0011000110000101111000",
			6054 => "0001000011111001110100",
			6055 => "0011000000101000111100",
			6056 => "0011000100010100011100",
			6057 => "0011000100010100010000",
			6058 => "0010100001010000001000",
			6059 => "0000100101110000000100",
			6060 => "0000000101111111010001",
			6061 => "0000000101111111010001",
			6062 => "0001001001001100000100",
			6063 => "0000001101111111010001",
			6064 => "0000000101111111010001",
			6065 => "0001000001101100001000",
			6066 => "0001000011000000000100",
			6067 => "1111110101111111010001",
			6068 => "0000000101111111010001",
			6069 => "0000010101111111010001",
			6070 => "0011000100010100010000",
			6071 => "0000110011011100001000",
			6072 => "0011010110000100000100",
			6073 => "0000001101111111010001",
			6074 => "1111111101111111010001",
			6075 => "0011011101111000000100",
			6076 => "0000001101111111010001",
			6077 => "0000001101111111010001",
			6078 => "0001000100001100001000",
			6079 => "0010000001110100000100",
			6080 => "0000000101111111010001",
			6081 => "0000001101111111010001",
			6082 => "0000011110100000000100",
			6083 => "0000000101111111010001",
			6084 => "1111111101111111010001",
			6085 => "0011000000101000011000",
			6086 => "0011011010111100010000",
			6087 => "0010001011010100001000",
			6088 => "0000101100100100000100",
			6089 => "0000000101111111010001",
			6090 => "1111111101111111010001",
			6091 => "0001011100101000000100",
			6092 => "0000000101111111010001",
			6093 => "0000001101111111010001",
			6094 => "0011010111001000000100",
			6095 => "1111111101111111010001",
			6096 => "1111111101111111010001",
			6097 => "0011101001110000010000",
			6098 => "0011110111010000001000",
			6099 => "0011100000111000000100",
			6100 => "0000000101111111010001",
			6101 => "0000001101111111010001",
			6102 => "0001010101101100000100",
			6103 => "0000001101111111010001",
			6104 => "0000000101111111010001",
			6105 => "0010011101101000001000",
			6106 => "0011001000111100000100",
			6107 => "0000001101111111010001",
			6108 => "1111111101111111010001",
			6109 => "0001001001001100000100",
			6110 => "0000000101111111010001",
			6111 => "0000000101111111010001",
			6112 => "1111111101111111010001",
			6113 => "0011001010111100100100",
			6114 => "0001111011000000011000",
			6115 => "0001110100011000010000",
			6116 => "0001111101111000001100",
			6117 => "0001111110001100000100",
			6118 => "1111111101111111010001",
			6119 => "0011000110000100000100",
			6120 => "0000000101111111010001",
			6121 => "0000000101111111010001",
			6122 => "1111111101111111010001",
			6123 => "0011000100001000000100",
			6124 => "0000001101111111010001",
			6125 => "1111111101111111010001",
			6126 => "0001111000000000000100",
			6127 => "0000011101111111010001",
			6128 => "0001001011110000000100",
			6129 => "0000000101111111010001",
			6130 => "0000001101111111010001",
			6131 => "1111111101111111010001",
			6132 => "0011001000111010011100",
			6133 => "0001000100001101011100",
			6134 => "0000110100000000101100",
			6135 => "0010110100010100010100",
			6136 => "0001001110000000000100",
			6137 => "0000011110000101110101",
			6138 => "0000111010000000001000",
			6139 => "0010110100010100000100",
			6140 => "1111111110000101110101",
			6141 => "0000000110000101110101",
			6142 => "0010011100110100000100",
			6143 => "0000011110000101110101",
			6144 => "0000000110000101110101",
			6145 => "0011100000111000001100",
			6146 => "0011001010000000000100",
			6147 => "0000001110000101110101",
			6148 => "0000001010000000000100",
			6149 => "0000000110000101110101",
			6150 => "1111111110000101110101",
			6151 => "0010101000010100000100",
			6152 => "1111111110000101110101",
			6153 => "0011111111011100000100",
			6154 => "0000011110000101110101",
			6155 => "0000000110000101110101",
			6156 => "0000110001011000011100",
			6157 => "0010100111110100001100",
			6158 => "0001101101111100001000",
			6159 => "0001101011111100000100",
			6160 => "1111111110000101110101",
			6161 => "0000000110000101110101",
			6162 => "0000010110000101110101",
			6163 => "0001000110001100001000",
			6164 => "0000111101100000000100",
			6165 => "0000001110000101110101",
			6166 => "0000010110000101110101",
			6167 => "0010001001101000000100",
			6168 => "0000000110000101110101",
			6169 => "0000001110000101110101",
			6170 => "0000001000101100000100",
			6171 => "0000010110000101110101",
			6172 => "0000000000110000001000",
			6173 => "0010110000001100000100",
			6174 => "1111111110000101110101",
			6175 => "0000001110000101110101",
			6176 => "0000010111100100000100",
			6177 => "0000001110000101110101",
			6178 => "1111111110000101110101",
			6179 => "0010010110000000000100",
			6180 => "1111111110000101110101",
			6181 => "0000101100010100011100",
			6182 => "0010110111111000001100",
			6183 => "0001100001111000000100",
			6184 => "1111111110000101110101",
			6185 => "0000101101000100000100",
			6186 => "0000000110000101110101",
			6187 => "0000010110000101110101",
			6188 => "0000001011000100001000",
			6189 => "0010001010101100000100",
			6190 => "0000000110000101110101",
			6191 => "0000010110000101110101",
			6192 => "0001000011011000000100",
			6193 => "0000000110000101110101",
			6194 => "0000001110000101110101",
			6195 => "0001000011101100010000",
			6196 => "0010101100011100001000",
			6197 => "0011000111111000000100",
			6198 => "0000001110000101110101",
			6199 => "1111111110000101110101",
			6200 => "0010011101011100000100",
			6201 => "0000001110000101110101",
			6202 => "1111111110000101110101",
			6203 => "0011101110001100001000",
			6204 => "0010101011010100000100",
			6205 => "1111111110000101110101",
			6206 => "0000000110000101110101",
			6207 => "0000110011100000000100",
			6208 => "0000001110000101110101",
			6209 => "1111111110000101110101",
			6210 => "0011001100110000101100",
			6211 => "0011111101000100001100",
			6212 => "0000110111001000001000",
			6213 => "0001011010111000000100",
			6214 => "0000000110000101110101",
			6215 => "1111111110000101110101",
			6216 => "1111111110000101110101",
			6217 => "0000101000001100011000",
			6218 => "0010110100001000010000",
			6219 => "0000010110101000001000",
			6220 => "0010111101111000000100",
			6221 => "0000000110000101110101",
			6222 => "0000010110000101110101",
			6223 => "0010111101111000000100",
			6224 => "0000000110000101110101",
			6225 => "1111111110000101110101",
			6226 => "0001011010001100000100",
			6227 => "0000010110000101110101",
			6228 => "0000000110000101110101",
			6229 => "0010100001010000000100",
			6230 => "0000001110000101110101",
			6231 => "1111111110000101110101",
			6232 => "0011000100001000001000",
			6233 => "0011000000001100000100",
			6234 => "1111111110000101110101",
			6235 => "0000000110000101110101",
			6236 => "1111111110000101110101",
			6237 => "0001110110000110001000",
			6238 => "0000010000011000001000",
			6239 => "0001100100110100000100",
			6240 => "1111111110001011011001",
			6241 => "0000001110001011011001",
			6242 => "0010011001111001000000",
			6243 => "0000110100000000100000",
			6244 => "0010011001111000010000",
			6245 => "0000110100010100001000",
			6246 => "0010100111110100000100",
			6247 => "0000010110001011011001",
			6248 => "0000000110001011011001",
			6249 => "0010010010001100000100",
			6250 => "0000001110001011011001",
			6251 => "0000000110001011011001",
			6252 => "0000011110100000001000",
			6253 => "0001010011011100000100",
			6254 => "0000000110001011011001",
			6255 => "1111111110001011011001",
			6256 => "0000011110100000000100",
			6257 => "0000010110001011011001",
			6258 => "0000000110001011011001",
			6259 => "0011110110110100010000",
			6260 => "0010001100000100001000",
			6261 => "0010111011000100000100",
			6262 => "1111111110001011011001",
			6263 => "0000000110001011011001",
			6264 => "0010101010110000000100",
			6265 => "0000001110001011011001",
			6266 => "0000011110001011011001",
			6267 => "0000111000111000001000",
			6268 => "0010010010001100000100",
			6269 => "0000001110001011011001",
			6270 => "1111111110001011011001",
			6271 => "0001110100010100000100",
			6272 => "0000001110001011011001",
			6273 => "0000000110001011011001",
			6274 => "0011101000111100100000",
			6275 => "0010010110101000010000",
			6276 => "0000110011011100001000",
			6277 => "0011110110110100000100",
			6278 => "0000000110001011011001",
			6279 => "1111111110001011011001",
			6280 => "0010110100000000000100",
			6281 => "0000000110001011011001",
			6282 => "0000010110001011011001",
			6283 => "0011111010010100001000",
			6284 => "0001010110000100000100",
			6285 => "0000001110001011011001",
			6286 => "0000000110001011011001",
			6287 => "0001000011010100000100",
			6288 => "1111111110001011011001",
			6289 => "0000000110001011011001",
			6290 => "0010011101101000010000",
			6291 => "0000100010000000001000",
			6292 => "0010101100011100000100",
			6293 => "0000000110001011011001",
			6294 => "0000001110001011011001",
			6295 => "0010000001110100000100",
			6296 => "0000000110001011011001",
			6297 => "0000000110001011011001",
			6298 => "0011101101111000001000",
			6299 => "0000100100101000000100",
			6300 => "0000000110001011011001",
			6301 => "0000000110001011011001",
			6302 => "0010011111001100000100",
			6303 => "0000000110001011011001",
			6304 => "0000000110001011011001",
			6305 => "0001111100101000011000",
			6306 => "0010110001111100000100",
			6307 => "1111111110001011011001",
			6308 => "0000100111010100010000",
			6309 => "0000100010000000000100",
			6310 => "1111111110001011011001",
			6311 => "0001001000110100000100",
			6312 => "0000000110001011011001",
			6313 => "0000110001001000000100",
			6314 => "0000000110001011011001",
			6315 => "0000010110001011011001",
			6316 => "1111111110001011011001",
			6317 => "0010100111110100010000",
			6318 => "0000100001011100001100",
			6319 => "0001110001111100001000",
			6320 => "0011110001011000000100",
			6321 => "0000000110001011011001",
			6322 => "0000000110001011011001",
			6323 => "1111111110001011011001",
			6324 => "0000010110001011011001",
			6325 => "1111111110001011011001",
			6326 => "0000001100001010100100",
			6327 => "0000100010110101000000",
			6328 => "0000100001001000011100",
			6329 => "0000001000110000010100",
			6330 => "0010111011000100000100",
			6331 => "0000001110010010110101",
			6332 => "0011001011000100001000",
			6333 => "0000001011010100000100",
			6334 => "0000000110010010110101",
			6335 => "1111111110010010110101",
			6336 => "0001101011111100000100",
			6337 => "0000000110010010110101",
			6338 => "0000001110010010110101",
			6339 => "0011001010000000000100",
			6340 => "0000000110010010110101",
			6341 => "1111111110010010110101",
			6342 => "0010110100010100010000",
			6343 => "0011010011011100001100",
			6344 => "0011111001110100001000",
			6345 => "0011111011000000000100",
			6346 => "0000001110010010110101",
			6347 => "1111111110010010110101",
			6348 => "0000001110010010110101",
			6349 => "1111111110010010110101",
			6350 => "0000001110111100010000",
			6351 => "0010101000010100001000",
			6352 => "0000001000110000000100",
			6353 => "0000000110010010110101",
			6354 => "0000001110010010110101",
			6355 => "0010101001000100000100",
			6356 => "1111111110010010110101",
			6357 => "0000000110010010110101",
			6358 => "0000001110010010110101",
			6359 => "0010101100011100110100",
			6360 => "0001011001110100100000",
			6361 => "0000101001100000010000",
			6362 => "0011110110100000001000",
			6363 => "0011110010110100000100",
			6364 => "0000000110010010110101",
			6365 => "0000000110010010110101",
			6366 => "0011100001111100000100",
			6367 => "0000001110010010110101",
			6368 => "0000000110010010110101",
			6369 => "0001011010111100001000",
			6370 => "0001010101101100000100",
			6371 => "0000001110010010110101",
			6372 => "0000000110010010110101",
			6373 => "0010011101011100000100",
			6374 => "0000000110010010110101",
			6375 => "1111111110010010110101",
			6376 => "0010010101011100000100",
			6377 => "0000001110010010110101",
			6378 => "0010111110001100001000",
			6379 => "0001111001110000000100",
			6380 => "0000000110010010110101",
			6381 => "0000001110010010110101",
			6382 => "0010011011111100000100",
			6383 => "1111111110010010110101",
			6384 => "0000000110010010110101",
			6385 => "0001011100110000010100",
			6386 => "0001101100011000001000",
			6387 => "0000001011000100000100",
			6388 => "0000001110010010110101",
			6389 => "1111111110010010110101",
			6390 => "0001010011011100000100",
			6391 => "0000000110010010110101",
			6392 => "0010011001111000000100",
			6393 => "0000001110010010110101",
			6394 => "0000000110010010110101",
			6395 => "0011000100010100001100",
			6396 => "0001001111100000001000",
			6397 => "0011101100001000000100",
			6398 => "1111111110010010110101",
			6399 => "0000001110010010110101",
			6400 => "1111111110010010110101",
			6401 => "0010010111100100001000",
			6402 => "0000111101111000000100",
			6403 => "0000000110010010110101",
			6404 => "0000001110010010110101",
			6405 => "0001101101011000000100",
			6406 => "0000000110010010110101",
			6407 => "0000000110010010110101",
			6408 => "0000100010000000101100",
			6409 => "0011100000101000101000",
			6410 => "0011000100010100011000",
			6411 => "0000110100000000010000",
			6412 => "0000111011000100001000",
			6413 => "0010100110011100000100",
			6414 => "1111111110010010110101",
			6415 => "0000000110010010110101",
			6416 => "0010100110011100000100",
			6417 => "0000001110010010110101",
			6418 => "0000000110010010110101",
			6419 => "0010100101000100000100",
			6420 => "1111111110010010110101",
			6421 => "0000000110010010110101",
			6422 => "0000101010001000000100",
			6423 => "1111111110010010110101",
			6424 => "0000101010001000001000",
			6425 => "0001101010011000000100",
			6426 => "0000000110010010110101",
			6427 => "0000001110010010110101",
			6428 => "1111111110010010110101",
			6429 => "0000001110010010110101",
			6430 => "0001011110001100000100",
			6431 => "1111111110010010110101",
			6432 => "0010010110101000001100",
			6433 => "0000100010000100000100",
			6434 => "0000000110010010110101",
			6435 => "0000000001101000000100",
			6436 => "0000001110010010110101",
			6437 => "0000000110010010110101",
			6438 => "0011001001110000001000",
			6439 => "0011101001001000000100",
			6440 => "1111111110010010110101",
			6441 => "0000000110010010110101",
			6442 => "0000111010111000000100",
			6443 => "0000001110010010110101",
			6444 => "0000000110010010110101",
			6445 => "0010010110101010001000",
			6446 => "0010010110101001100000",
			6447 => "0000000000110000100100",
			6448 => "0010010110101000010100",
			6449 => "0011111010010100010000",
			6450 => "0001001010110100001000",
			6451 => "0000000000111000000100",
			6452 => "0000000110011010100001",
			6453 => "0000000110011010100001",
			6454 => "0011110101110100000100",
			6455 => "0000001110011010100001",
			6456 => "1111111110011010100001",
			6457 => "1111111110011010100001",
			6458 => "0000000000111000001100",
			6459 => "0000101001010000001000",
			6460 => "0001100001111000000100",
			6461 => "1111111110011010100001",
			6462 => "0000000110011010100001",
			6463 => "1111111110011010100001",
			6464 => "0000000110011010100001",
			6465 => "0000111100110000100000",
			6466 => "0011110110110100010000",
			6467 => "0000110100000000001000",
			6468 => "0010001111001000000100",
			6469 => "0000000110011010100001",
			6470 => "0000000110011010100001",
			6471 => "0011110000011100000100",
			6472 => "0000001110011010100001",
			6473 => "0000000110011010100001",
			6474 => "0001111011000100001000",
			6475 => "0000100100101000000100",
			6476 => "1111111110011010100001",
			6477 => "0000000110011010100001",
			6478 => "0011000111111000000100",
			6479 => "0000000110011010100001",
			6480 => "1111111110011010100001",
			6481 => "0011000100010100001100",
			6482 => "0010101100011100001000",
			6483 => "0010011001111000000100",
			6484 => "0000001110011010100001",
			6485 => "0000000110011010100001",
			6486 => "1111111110011010100001",
			6487 => "0000011110100000001000",
			6488 => "0011000000101000000100",
			6489 => "0000000110011010100001",
			6490 => "1111111110011010100001",
			6491 => "0011000100010100000100",
			6492 => "0000001110011010100001",
			6493 => "0000000110011010100001",
			6494 => "0001101100011000011100",
			6495 => "0000101110000100001000",
			6496 => "0010001100000100000100",
			6497 => "0000001110011010100001",
			6498 => "1111111110011010100001",
			6499 => "0000111101100000001000",
			6500 => "0000001010000000000100",
			6501 => "0000001110011010100001",
			6502 => "0000010110011010100001",
			6503 => "0011011100101100001000",
			6504 => "0000110101101100000100",
			6505 => "0000001110011010100001",
			6506 => "0000000110011010100001",
			6507 => "0000000110011010100001",
			6508 => "0000100101110000000100",
			6509 => "0000001110011010100001",
			6510 => "0000100011001000000100",
			6511 => "1111111110011010100001",
			6512 => "0000000110011010100001",
			6513 => "0000011110100000001100",
			6514 => "0011000111111000000100",
			6515 => "0000000110011010100001",
			6516 => "0000000000110000000100",
			6517 => "1111111110011010100001",
			6518 => "1111111110011010100001",
			6519 => "0000110101101100111000",
			6520 => "0011000000101000011100",
			6521 => "0000001010000000010000",
			6522 => "0001001000000100001000",
			6523 => "0001001011110000000100",
			6524 => "0000000110011010100001",
			6525 => "1111111110011010100001",
			6526 => "0000011100110100000100",
			6527 => "0000000110011010100001",
			6528 => "0000000110011010100001",
			6529 => "0011010110000100000100",
			6530 => "0000000110011010100001",
			6531 => "0001110100000000000100",
			6532 => "1111111110011010100001",
			6533 => "0000000110011010100001",
			6534 => "0011110101100100001100",
			6535 => "0011000000101000000100",
			6536 => "1111111110011010100001",
			6537 => "0011000100000000000100",
			6538 => "0000000110011010100001",
			6539 => "1111111110011010100001",
			6540 => "0011110101110100001000",
			6541 => "0000110101101100000100",
			6542 => "1111111110011010100001",
			6543 => "1111111110011010100001",
			6544 => "0001101100011000000100",
			6545 => "0000000110011010100001",
			6546 => "1111111110011010100001",
			6547 => "0000110110000100010000",
			6548 => "0000100100101000001000",
			6549 => "0000100101001000000100",
			6550 => "0000001110011010100001",
			6551 => "1111111110011010100001",
			6552 => "0010101010110000000100",
			6553 => "0000001110011010100001",
			6554 => "0000000110011010100001",
			6555 => "0000110110000100001100",
			6556 => "0001001010110100000100",
			6557 => "1111111110011010100001",
			6558 => "0011101011000100000100",
			6559 => "1111111110011010100001",
			6560 => "0000000110011010100001",
			6561 => "0011000111111000001000",
			6562 => "0011110111110000000100",
			6563 => "0000000110011010100001",
			6564 => "1111111110011010100001",
			6565 => "0000011110100000000100",
			6566 => "0000000110011010100001",
			6567 => "0000000110011010100001",
			6568 => "0011000011011101110000",
			6569 => "0001001011100101101100",
			6570 => "0000000100010100111100",
			6571 => "0001111011000100011100",
			6572 => "0001011100110000010000",
			6573 => "0011000111111000001000",
			6574 => "0010011110100000000100",
			6575 => "1111111110100000001101",
			6576 => "0000001110100000001101",
			6577 => "0001001111100000000100",
			6578 => "0000000110100000001101",
			6579 => "0000010110100000001101",
			6580 => "0000100000110100000100",
			6581 => "1111111110100000001101",
			6582 => "0010011001111000000100",
			6583 => "0000010110100000001101",
			6584 => "0000001110100000001101",
			6585 => "0001100111101000010000",
			6586 => "0010110100000000001000",
			6587 => "0001001000011100000100",
			6588 => "0000001110100000001101",
			6589 => "1111111110100000001101",
			6590 => "0010010001000100000100",
			6591 => "1111111110100000001101",
			6592 => "0000001110100000001101",
			6593 => "0001000011001100001000",
			6594 => "0001101101111100000100",
			6595 => "0000000110100000001101",
			6596 => "0000001110100000001101",
			6597 => "0010100110011000000100",
			6598 => "0000000110100000001101",
			6599 => "0000000110100000001101",
			6600 => "0001101010011000010100",
			6601 => "0001101010011000010000",
			6602 => "0000001000111100001000",
			6603 => "0000110100010100000100",
			6604 => "0000000110100000001101",
			6605 => "0000000110100000001101",
			6606 => "0011110111010000000100",
			6607 => "0000001110100000001101",
			6608 => "0000000110100000001101",
			6609 => "0000010110100000001101",
			6610 => "0000101100010000010000",
			6611 => "0000001011000100001000",
			6612 => "0000011100110100000100",
			6613 => "0000001110100000001101",
			6614 => "1111111110100000001101",
			6615 => "0011011010111000000100",
			6616 => "1111111110100000001101",
			6617 => "0000000110100000001101",
			6618 => "0001000011101100000100",
			6619 => "0000010110100000001101",
			6620 => "0011110001000000000100",
			6621 => "1111111110100000001101",
			6622 => "0000000110100000001101",
			6623 => "1111111110100000001101",
			6624 => "0011000110000100101000",
			6625 => "0000110110100100000100",
			6626 => "1111111110100000001101",
			6627 => "0000100111011000010100",
			6628 => "0001000010110000010000",
			6629 => "0010011011111100001000",
			6630 => "0011001100110000000100",
			6631 => "1111111110100000001101",
			6632 => "0000000110100000001101",
			6633 => "0010111010111100000100",
			6634 => "0000001110100000001101",
			6635 => "1111111110100000001101",
			6636 => "0000001110100000001101",
			6637 => "0011011001010100001100",
			6638 => "0001101001100100000100",
			6639 => "1111111110100000001101",
			6640 => "0000010111100100000100",
			6641 => "0000000110100000001101",
			6642 => "1111111110100000001101",
			6643 => "0000001110100000001101",
			6644 => "0011001010111100011100",
			6645 => "0001110110100100011000",
			6646 => "0001111101111000001100",
			6647 => "0000000011010000001000",
			6648 => "0001111110001100000100",
			6649 => "1111111110100000001101",
			6650 => "0000001110100000001101",
			6651 => "1111111110100000001101",
			6652 => "0001110100011000000100",
			6653 => "1111111110100000001101",
			6654 => "0001110100011000000100",
			6655 => "0000000110100000001101",
			6656 => "1111111110100000001101",
			6657 => "0000001110100000001101",
			6658 => "1111111110100000001101",
			6659 => "0011000110000110101100",
			6660 => "0010010110101001100100",
			6661 => "0011000100010100111100",
			6662 => "0000101110101000011100",
			6663 => "0011100000110000010000",
			6664 => "0001110000101000001000",
			6665 => "0000110010111100000100",
			6666 => "0000000110100101111001",
			6667 => "0000000110100101111001",
			6668 => "0010100001010000000100",
			6669 => "1111111110100101111001",
			6670 => "0000001110100101111001",
			6671 => "0000000011111100001000",
			6672 => "0010110000101000000100",
			6673 => "0000000110100101111001",
			6674 => "0000001110100101111001",
			6675 => "0000010110100101111001",
			6676 => "0010100110011000010000",
			6677 => "0000100101110000001000",
			6678 => "0010001011010100000100",
			6679 => "0000000110100101111001",
			6680 => "0000000110100101111001",
			6681 => "0000000000111000000100",
			6682 => "1111111110100101111001",
			6683 => "0000001110100101111001",
			6684 => "0001000010111000001000",
			6685 => "0000100101110000000100",
			6686 => "0000001110100101111001",
			6687 => "0000000110100101111001",
			6688 => "0011011110001100000100",
			6689 => "0000000110100101111001",
			6690 => "0000001110100101111001",
			6691 => "0000011100110100100000",
			6692 => "0011101110111100010000",
			6693 => "0011010101101100001000",
			6694 => "0010111011000100000100",
			6695 => "0000000110100101111001",
			6696 => "0000010110100101111001",
			6697 => "0000101001010000000100",
			6698 => "0000000110100101111001",
			6699 => "1111111110100101111001",
			6700 => "0000101110010000001000",
			6701 => "0010100110011100000100",
			6702 => "0000001110100101111001",
			6703 => "0000011110100101111001",
			6704 => "0001110000101000000100",
			6705 => "0000000110100101111001",
			6706 => "1111111110100101111001",
			6707 => "0011000000101000000100",
			6708 => "0000001110100101111001",
			6709 => "0000011110100101111001",
			6710 => "0000011110100000001100",
			6711 => "0000100011001000001000",
			6712 => "0001111011000100000100",
			6713 => "1111111110100101111001",
			6714 => "1111110110100101111001",
			6715 => "0000000110100101111001",
			6716 => "0000111101111000011100",
			6717 => "0010011101101000010000",
			6718 => "0001111100001000001000",
			6719 => "0001111011000100000100",
			6720 => "0000000110100101111001",
			6721 => "0000000110100101111001",
			6722 => "0000110011011100000100",
			6723 => "1111111110100101111001",
			6724 => "0000000110100101111001",
			6725 => "0011101100110000001000",
			6726 => "0010110100000000000100",
			6727 => "1111111110100101111001",
			6728 => "0000000110100101111001",
			6729 => "1111110110100101111001",
			6730 => "0010010111100100010000",
			6731 => "0011000000101000001000",
			6732 => "0000100110010000000100",
			6733 => "0000001110100101111001",
			6734 => "0000000110100101111001",
			6735 => "0000011100110100000100",
			6736 => "0000001110100101111001",
			6737 => "0000010110100101111001",
			6738 => "0000110000001100001000",
			6739 => "0010011101101000000100",
			6740 => "0000001110100101111001",
			6741 => "1111111110100101111001",
			6742 => "0011101101100000000100",
			6743 => "0000000110100101111001",
			6744 => "0000000110100101111001",
			6745 => "0011001010111100001000",
			6746 => "0001011110101000000100",
			6747 => "1111111110100101111001",
			6748 => "0000001110100101111001",
			6749 => "1111111110100101111001",
			6750 => "0011000110000110111100",
			6751 => "0010011101101001011100",
			6752 => "0001110000101000110100",
			6753 => "0001110000101000011000",
			6754 => "0011000000101000010000",
			6755 => "0000100001000000001000",
			6756 => "0000000100010100000100",
			6757 => "0000000110101100000101",
			6758 => "0000000110101100000101",
			6759 => "0010101001000100000100",
			6760 => "1111111110101100000101",
			6761 => "0000000110101100000101",
			6762 => "0001001110111000000100",
			6763 => "0000000110101100000101",
			6764 => "0000010110101100000101",
			6765 => "0010101010110000010000",
			6766 => "0011000100010100001000",
			6767 => "0011111011011100000100",
			6768 => "1111111110101100000101",
			6769 => "1111111110101100000101",
			6770 => "0000101100100100000100",
			6771 => "1111111110101100000101",
			6772 => "0000000110101100000101",
			6773 => "0011000111111000000100",
			6774 => "1111111110101100000101",
			6775 => "0001010110000100000100",
			6776 => "0000001110101100000101",
			6777 => "0000000110101100000101",
			6778 => "0010100111110100001100",
			6779 => "0000011100110100001000",
			6780 => "0001111100001000000100",
			6781 => "1111111110101100000101",
			6782 => "1111111110101100000101",
			6783 => "0000001110101100000101",
			6784 => "0001000011001100010000",
			6785 => "0011000111111000001000",
			6786 => "0011100100000000000100",
			6787 => "1111111110101100000101",
			6788 => "0000000110101100000101",
			6789 => "0010010111100100000100",
			6790 => "0000001110101100000101",
			6791 => "0000000110101100000101",
			6792 => "0011011101100000000100",
			6793 => "0000010110101100000101",
			6794 => "0011101100001000000100",
			6795 => "0000000110101100000101",
			6796 => "0000000110101100000101",
			6797 => "0011100110000100110000",
			6798 => "0000011100110100010000",
			6799 => "0001001100001100000100",
			6800 => "1111110110101100000101",
			6801 => "0000100100101000000100",
			6802 => "0000001110101100000101",
			6803 => "0001001010110100000100",
			6804 => "1111110110101100000101",
			6805 => "1111111110101100000101",
			6806 => "0011011101010100010000",
			6807 => "0011110001001000001000",
			6808 => "0011101101100000000100",
			6809 => "0000000110101100000101",
			6810 => "0000000110101100000101",
			6811 => "0010000110001000000100",
			6812 => "1111111110101100000101",
			6813 => "0000000110101100000101",
			6814 => "0011001000111000001000",
			6815 => "0011111110101100000100",
			6816 => "1111111110101100000101",
			6817 => "0000000110101100000101",
			6818 => "0010000111000100000100",
			6819 => "1111111110101100000101",
			6820 => "0000010110101100000101",
			6821 => "0010011101101000011000",
			6822 => "0000101001100000001100",
			6823 => "0011110110100000001000",
			6824 => "0011000000101000000100",
			6825 => "0000001110101100000101",
			6826 => "0000000110101100000101",
			6827 => "0000001110101100000101",
			6828 => "0010000001110100000100",
			6829 => "1111111110101100000101",
			6830 => "0010111000111000000100",
			6831 => "0000000110101100000101",
			6832 => "0000001110101100000101",
			6833 => "0011111011110100001100",
			6834 => "0011000000101000000100",
			6835 => "0000000110101100000101",
			6836 => "0011110101110100000100",
			6837 => "1111111110101100000101",
			6838 => "1111110110101100000101",
			6839 => "0011110111110000000100",
			6840 => "0000001110101100000101",
			6841 => "0011101101111000000100",
			6842 => "0000000110101100000101",
			6843 => "0000000110101100000101",
			6844 => "0010100111110100001000",
			6845 => "0000100001011100000100",
			6846 => "1111111110101100000101",
			6847 => "0000001110101100000101",
			6848 => "1111111110101100000101",
			6849 => "0011000110000111000000",
			6850 => "0011111011011101010000",
			6851 => "0000111100110000101000",
			6852 => "0010010110101000011000",
			6853 => "0000011100110100010000",
			6854 => "0010010110101000001000",
			6855 => "0000110100000000000100",
			6856 => "0000000110110010011001",
			6857 => "0000000110110010011001",
			6858 => "0011011100101100000100",
			6859 => "0000000110110010011001",
			6860 => "0000000110110010011001",
			6861 => "0011000100010100000100",
			6862 => "0000010110110010011001",
			6863 => "0000000110110010011001",
			6864 => "0011100111111000000100",
			6865 => "1111111110110010011001",
			6866 => "0000101110000100001000",
			6867 => "0011011101111000000100",
			6868 => "0000001110110010011001",
			6869 => "1111111110110010011001",
			6870 => "1111111110110010011001",
			6871 => "0011010001111100011100",
			6872 => "0001000010111000001100",
			6873 => "0010001011010100001000",
			6874 => "0011110111010000000100",
			6875 => "0000001110110010011001",
			6876 => "0000000110110010011001",
			6877 => "1111111110110010011001",
			6878 => "0000101111010000001000",
			6879 => "0011110101100100000100",
			6880 => "0000010110110010011001",
			6881 => "0000001110110010011001",
			6882 => "0011100100010100000100",
			6883 => "0000000110110010011001",
			6884 => "0000010110110010011001",
			6885 => "0011101100110000000100",
			6886 => "1111111110110010011001",
			6887 => "0001100101011100000100",
			6888 => "0000000110110010011001",
			6889 => "0000001110110010011001",
			6890 => "0001100100110101000000",
			6891 => "0000111010111100100000",
			6892 => "0011101101100000010000",
			6893 => "0010001001101000001000",
			6894 => "0000110101101100000100",
			6895 => "1111111110110010011001",
			6896 => "0000000110110010011001",
			6897 => "0011101001110000000100",
			6898 => "0000000110110010011001",
			6899 => "1111111110110010011001",
			6900 => "0011010001111100001000",
			6901 => "0010001001101000000100",
			6902 => "0000001110110010011001",
			6903 => "0000000110110010011001",
			6904 => "0011110111110000000100",
			6905 => "1111111110110010011001",
			6906 => "0000000110110010011001",
			6907 => "0011101100101000010000",
			6908 => "0000100010011100001000",
			6909 => "0000100101001000000100",
			6910 => "1111111110110010011001",
			6911 => "0000000110110010011001",
			6912 => "0010011101101000000100",
			6913 => "0000000110110010011001",
			6914 => "1111111110110010011001",
			6915 => "0010100111110100001000",
			6916 => "0001001011101100000100",
			6917 => "0000000110110010011001",
			6918 => "1111111110110010011001",
			6919 => "0000101110010000000100",
			6920 => "0000001110110010011001",
			6921 => "0000000110110010011001",
			6922 => "0011001010000000010100",
			6923 => "0001100100110100001000",
			6924 => "0000100111111100000100",
			6925 => "1111111110110010011001",
			6926 => "0000000110110010011001",
			6927 => "0000101010001000000100",
			6928 => "0000000110110010011001",
			6929 => "0011010110000100000100",
			6930 => "1111111110110010011001",
			6931 => "1111110110110010011001",
			6932 => "0011001110111100001100",
			6933 => "0000101100010100001000",
			6934 => "0010101010110000000100",
			6935 => "0000001110110010011001",
			6936 => "0000000110110010011001",
			6937 => "0000001110110010011001",
			6938 => "0010000001110000001000",
			6939 => "0000101100010100000100",
			6940 => "0000001110110010011001",
			6941 => "0000000110110010011001",
			6942 => "0000001000110000000100",
			6943 => "1111111110110010011001",
			6944 => "0000000110110010011001",
			6945 => "0010100111110100001000",
			6946 => "0000100001011100000100",
			6947 => "1111111110110010011001",
			6948 => "0000001110110010011001",
			6949 => "1111111110110010011001",
			6950 => "0010000111000010011100",
			6951 => "0010100110011101111000",
			6952 => "0010011001111000111100",
			6953 => "0001011101100000100000",
			6954 => "0000000000110000010000",
			6955 => "0001110111111000001000",
			6956 => "0001011000111100000100",
			6957 => "0000001110111001010101",
			6958 => "1111111110111001010101",
			6959 => "0010100110011000000100",
			6960 => "0000000110111001010101",
			6961 => "0000001110111001010101",
			6962 => "0000000000110000001000",
			6963 => "0011000111111000000100",
			6964 => "1111111110111001010101",
			6965 => "0000000110111001010101",
			6966 => "0011100010011000000100",
			6967 => "0000000110111001010101",
			6968 => "0000000110111001010101",
			6969 => "0010100110011000010000",
			6970 => "0010010010001100001000",
			6971 => "0010010010001100000100",
			6972 => "1111111110111001010101",
			6973 => "0000001110111001010101",
			6974 => "0011100000110000000100",
			6975 => "1111111110111001010101",
			6976 => "0000000110111001010101",
			6977 => "0000010110000000000100",
			6978 => "0000000110111001010101",
			6979 => "0000001110111100000100",
			6980 => "0000001110111001010101",
			6981 => "0000001110111001010101",
			6982 => "0000011110100000011100",
			6983 => "0001011100110000010000",
			6984 => "0001010011011100001000",
			6985 => "0001100100110100000100",
			6986 => "0000000110111001010101",
			6987 => "0000001110111001010101",
			6988 => "0011110100010000000100",
			6989 => "0000000110111001010101",
			6990 => "1111111110111001010101",
			6991 => "0001110100010100000100",
			6992 => "0000001110111001010101",
			6993 => "0011100000110000000100",
			6994 => "1111111110111001010101",
			6995 => "0000000110111001010101",
			6996 => "0010010110101000010000",
			6997 => "0001110100010100001000",
			6998 => "0010010110101000000100",
			6999 => "0000000110111001010101",
			7000 => "1111111110111001010101",
			7001 => "0010010110101000000100",
			7002 => "0000000110111001010101",
			7003 => "0000001110111001010101",
			7004 => "0011100000101000001000",
			7005 => "0001100001111000000100",
			7006 => "0000000110111001010101",
			7007 => "0000000110111001010101",
			7008 => "0010100110011100000100",
			7009 => "0000000110111001010101",
			7010 => "0000000110111001010101",
			7011 => "0010010110101000000100",
			7012 => "0000010110111001010101",
			7013 => "0010111000111100001000",
			7014 => "0000000000101000000100",
			7015 => "0000000110111001010101",
			7016 => "1111111110111001010101",
			7017 => "0001010100001000001000",
			7018 => "0011101101100000000100",
			7019 => "0000000110111001010101",
			7020 => "0000001110111001010101",
			7021 => "0011111001010000001000",
			7022 => "0001101001100100000100",
			7023 => "1111111110111001010101",
			7024 => "0000000110111001010101",
			7025 => "0000011001111000000100",
			7026 => "0000001110111001010101",
			7027 => "1111111110111001010101",
			7028 => "0000101100000001000000",
			7029 => "0000101001100000101100",
			7030 => "0011111111011100011000",
			7031 => "0011101000110000010000",
			7032 => "0011001010000000001000",
			7033 => "0000101110101000000100",
			7034 => "0000000110111001010101",
			7035 => "0000001110111001010101",
			7036 => "0001100100110100000100",
			7037 => "0000000110111001010101",
			7038 => "1111111110111001010101",
			7039 => "0000011110100000000100",
			7040 => "0000001110111001010101",
			7041 => "1111111110111001010101",
			7042 => "0001111011000100001000",
			7043 => "0000101010001000000100",
			7044 => "1111111110111001010101",
			7045 => "0000000110111001010101",
			7046 => "0010111100001000001000",
			7047 => "0011010110000100000100",
			7048 => "1111111110111001010101",
			7049 => "0000000110111001010101",
			7050 => "1111111110111001010101",
			7051 => "0001011110001100000100",
			7052 => "1111111110111001010101",
			7053 => "0001101010011000001000",
			7054 => "0001111010111100000100",
			7055 => "0000010110111001010101",
			7056 => "0000000110111001010101",
			7057 => "0001101011001100000100",
			7058 => "0000000110111001010101",
			7059 => "0000001110111001010101",
			7060 => "1111111110111001010101",
			7061 => "0011000011011111001000",
			7062 => "0000101110101001011000",
			7063 => "0000010110000000101100",
			7064 => "0011000111111000011100",
			7065 => "0001111110111100001100",
			7066 => "0010111010000000001000",
			7067 => "0000011110011100000100",
			7068 => "1111111111000000100001",
			7069 => "0000000111000000100001",
			7070 => "1111111111000000100001",
			7071 => "0001110111111000001000",
			7072 => "0010110111111000000100",
			7073 => "0000001111000000100001",
			7074 => "0000000111000000100001",
			7075 => "0011000111111000000100",
			7076 => "0000000111000000100001",
			7077 => "0000010111000000100001",
			7078 => "0001111011000100001000",
			7079 => "0001111110111100000100",
			7080 => "0000000111000000100001",
			7081 => "1111111111000000100001",
			7082 => "0010110100010100000100",
			7083 => "0000001111000000100001",
			7084 => "1111111111000000100001",
			7085 => "0010010010001100010000",
			7086 => "0001110100010100001000",
			7087 => "0000001110111100000100",
			7088 => "0000001111000000100001",
			7089 => "0000000111000000100001",
			7090 => "0001010011011100000100",
			7091 => "0000001111000000100001",
			7092 => "0000010111000000100001",
			7093 => "0001100111101000010000",
			7094 => "0011011100101100001000",
			7095 => "0011110000011100000100",
			7096 => "0000000111000000100001",
			7097 => "0000001111000000100001",
			7098 => "0001001111100100000100",
			7099 => "0000000111000000100001",
			7100 => "1111111111000000100001",
			7101 => "0000010010001100001000",
			7102 => "0011011100101000000100",
			7103 => "0000000111000000100001",
			7104 => "1111111111000000100001",
			7105 => "0000001111000000100001",
			7106 => "0011111001010001000000",
			7107 => "0011010111001000100000",
			7108 => "0011000100010100010000",
			7109 => "0011000100010100001000",
			7110 => "0001111100001000000100",
			7111 => "0000000111000000100001",
			7112 => "0000000111000000100001",
			7113 => "0011010001111100000100",
			7114 => "0000000111000000100001",
			7115 => "1111111111000000100001",
			7116 => "0010111100001000001000",
			7117 => "0001100001111000000100",
			7118 => "0000000111000000100001",
			7119 => "0000001111000000100001",
			7120 => "0010111100001000000100",
			7121 => "0000000111000000100001",
			7122 => "0000000111000000100001",
			7123 => "0001001000011100010000",
			7124 => "0000001101010000001000",
			7125 => "0001000000010000000100",
			7126 => "0000001111000000100001",
			7127 => "0000000111000000100001",
			7128 => "0010100110011000000100",
			7129 => "0000001111000000100001",
			7130 => "0000000111000000100001",
			7131 => "0000000010011000001000",
			7132 => "0000100011001000000100",
			7133 => "1111110111000000100001",
			7134 => "1111111111000000100001",
			7135 => "0010011101011100000100",
			7136 => "0000000111000000100001",
			7137 => "1111111111000000100001",
			7138 => "0010001111001000011100",
			7139 => "0000000010011000010000",
			7140 => "0011000100000000001000",
			7141 => "0011000100000000000100",
			7142 => "0000001111000000100001",
			7143 => "0000100111000000100001",
			7144 => "0010110100001000000100",
			7145 => "1111111111000000100001",
			7146 => "0000001111000000100001",
			7147 => "0011001001110000001000",
			7148 => "0001001100001100000100",
			7149 => "1111111111000000100001",
			7150 => "0000000111000000100001",
			7151 => "0000001111000000100001",
			7152 => "0001001001000000010000",
			7153 => "0001101101011000001000",
			7154 => "0001101101011000000100",
			7155 => "0000000111000000100001",
			7156 => "0000001111000000100001",
			7157 => "0011110111111100000100",
			7158 => "0000000111000000100001",
			7159 => "0000001111000000100001",
			7160 => "1111111111000000100001",
			7161 => "0011001010111100011100",
			7162 => "0001011110101000011000",
			7163 => "0011000110000100010100",
			7164 => "0000100111011000001100",
			7165 => "0000101001100000001000",
			7166 => "0011001100110000000100",
			7167 => "1111111111000000100001",
			7168 => "0000000111000000100001",
			7169 => "0000000111000000100001",
			7170 => "0010110011100000000100",
			7171 => "1111111111000000100001",
			7172 => "0000000111000000100001",
			7173 => "1111111111000000100001",
			7174 => "0000001111000000100001",
			7175 => "1111111111000000100001",
			7176 => "0011001000111011010100",
			7177 => "0011000111111001101000",
			7178 => "0010010110101000111100",
			7179 => "0000111001110000100000",
			7180 => "0001111011000100010000",
			7181 => "0000000010111100001000",
			7182 => "0001010011011100000100",
			7183 => "0000001111001001000101",
			7184 => "0000000111001001000101",
			7185 => "0000111011000100000100",
			7186 => "0000000111001001000101",
			7187 => "0000000111001001000101",
			7188 => "0011111010011100001000",
			7189 => "0000110100010100000100",
			7190 => "1111111111001001000101",
			7191 => "0000001111001001000101",
			7192 => "0000110100000000000100",
			7193 => "1111111111001001000101",
			7194 => "0000000111001001000101",
			7195 => "0011110010001000001100",
			7196 => "0010011001111000000100",
			7197 => "0000000111001001000101",
			7198 => "0011111011011100000100",
			7199 => "0000001111001001000101",
			7200 => "0000001111001001000101",
			7201 => "0001011101100000001000",
			7202 => "0000100011001000000100",
			7203 => "0000000111001001000101",
			7204 => "0000001111001001000101",
			7205 => "0010101010110000000100",
			7206 => "0000000111001001000101",
			7207 => "0000000111001001000101",
			7208 => "0001011100110000010000",
			7209 => "0010110000101000001100",
			7210 => "0011101000111100001000",
			7211 => "0011110101110100000100",
			7212 => "0000000111001001000101",
			7213 => "1111111111001001000101",
			7214 => "0000000111001001000101",
			7215 => "1111110111001001000101",
			7216 => "0011001110111100001100",
			7217 => "0010101001000100000100",
			7218 => "1111111111001001000101",
			7219 => "0011001010000000000100",
			7220 => "0000000111001001000101",
			7221 => "0000001111001001000101",
			7222 => "0001111100001000001000",
			7223 => "0011101001110000000100",
			7224 => "0000000111001001000101",
			7225 => "0000000111001001000101",
			7226 => "0001011110001100000100",
			7227 => "0000001111001001000101",
			7228 => "0000000111001001000101",
			7229 => "0011000100010100101100",
			7230 => "0010101001000100010100",
			7231 => "0001110100010100000100",
			7232 => "0000001111001001000101",
			7233 => "0011000111111000001000",
			7234 => "0011111011011100000100",
			7235 => "1111111111001001000101",
			7236 => "1111111111001001000101",
			7237 => "0010010110101000000100",
			7238 => "0000000111001001000101",
			7239 => "0000001111001001000101",
			7240 => "0000100011001000010000",
			7241 => "0001110100010100001000",
			7242 => "0010111110111100000100",
			7243 => "1111111111001001000101",
			7244 => "0000000111001001000101",
			7245 => "0010011100110100000100",
			7246 => "1111111111001001000101",
			7247 => "0000001111001001000101",
			7248 => "0001101100011000000100",
			7249 => "0000000111001001000101",
			7250 => "0000001111001001000101",
			7251 => "0000111100110000100000",
			7252 => "0010010110101000010000",
			7253 => "0011000100010100001000",
			7254 => "0011000100010100000100",
			7255 => "0000000111001001000101",
			7256 => "0000000111001001000101",
			7257 => "0011110101100100000100",
			7258 => "0000000111001001000101",
			7259 => "0000000111001001000101",
			7260 => "0010001011010100001000",
			7261 => "0011011101111000000100",
			7262 => "0000000111001001000101",
			7263 => "1111111111001001000101",
			7264 => "0011110110110100000100",
			7265 => "1111111111001001000101",
			7266 => "0000000111001001000101",
			7267 => "0010010111100100010000",
			7268 => "0000111101111000001000",
			7269 => "0011111010010100000100",
			7270 => "0000000111001001000101",
			7271 => "0000000111001001000101",
			7272 => "0011000100010100000100",
			7273 => "0000000111001001000101",
			7274 => "0000001111001001000101",
			7275 => "0010111100001000001000",
			7276 => "0011000000101000000100",
			7277 => "0000000111001001000101",
			7278 => "0000000111001001000101",
			7279 => "0000110101101100000100",
			7280 => "1111111111001001000101",
			7281 => "0000000111001001000101",
			7282 => "0011111101000100011000",
			7283 => "0001011000000000001100",
			7284 => "0011100110000100001000",
			7285 => "0000000000111000000100",
			7286 => "0000001111001001000101",
			7287 => "1111111111001001000101",
			7288 => "1111111111001001000101",
			7289 => "0001011000000000001000",
			7290 => "0000100010011100000100",
			7291 => "0000000111001001000101",
			7292 => "0000010111001001000101",
			7293 => "1111111111001001000101",
			7294 => "0010011111001100001000",
			7295 => "0001101101011000000100",
			7296 => "0000001111001001000101",
			7297 => "1111111111001001000101",
			7298 => "0010111101111000000100",
			7299 => "1111111111001001000101",
			7300 => "0011111110010000010000",
			7301 => "0000101001100000001000",
			7302 => "0011010111010000000100",
			7303 => "1111111111001001000101",
			7304 => "0000001111001001000101",
			7305 => "0010010101011100000100",
			7306 => "0000001111001001000101",
			7307 => "0000000111001001000101",
			7308 => "0010100111110100001000",
			7309 => "0001111101010100000100",
			7310 => "0000001111001001000101",
			7311 => "0000000111001001000101",
			7312 => "1111111111001001000101",
			7313 => "0000100000010011000100",
			7314 => "0010101010110001101000",
			7315 => "0000000111111001000000",
			7316 => "0000101110101000100000",
			7317 => "0001100111101000010000",
			7318 => "0011000111111000001000",
			7319 => "0000001111000100000100",
			7320 => "0000001111001111100001",
			7321 => "0000000111001111100001",
			7322 => "0000111001110000000100",
			7323 => "1111111111001111100001",
			7324 => "0000000111001111100001",
			7325 => "0011000111111000001000",
			7326 => "0000110111111000000100",
			7327 => "1111111111001111100001",
			7328 => "0000000111001111100001",
			7329 => "0011110001101000000100",
			7330 => "0000001111001111100001",
			7331 => "0000000111001111100001",
			7332 => "0000010110000000010000",
			7333 => "0011011101100000001000",
			7334 => "0010110100010100000100",
			7335 => "0000000111001111100001",
			7336 => "0000000111001111100001",
			7337 => "0001110100010100000100",
			7338 => "0000001111001111100001",
			7339 => "1111111111001111100001",
			7340 => "0000111000111000001000",
			7341 => "0010110100010100000100",
			7342 => "0000000111001111100001",
			7343 => "0000000111001111100001",
			7344 => "0011110101110100000100",
			7345 => "0000000111001111100001",
			7346 => "0000000111001111100001",
			7347 => "0010111011000100100000",
			7348 => "0001101101111100010000",
			7349 => "0001000011110100001000",
			7350 => "0011011100110000000100",
			7351 => "1111111111001111100001",
			7352 => "0000000111001111100001",
			7353 => "0010000001110100000100",
			7354 => "1111111111001111100001",
			7355 => "0000001111001111100001",
			7356 => "0001100100110100001000",
			7357 => "0001000011010100000100",
			7358 => "0000000111001111100001",
			7359 => "0000001111001111100001",
			7360 => "0000100100101000000100",
			7361 => "0000000111001111100001",
			7362 => "1111111111001111100001",
			7363 => "0001000010100100000100",
			7364 => "1111111111001111100001",
			7365 => "0000000111001111100001",
			7366 => "0001001001001100100100",
			7367 => "0000101100000000011100",
			7368 => "0010111001110000010000",
			7369 => "0011110111110000001000",
			7370 => "0001000101010100000100",
			7371 => "1111111111001111100001",
			7372 => "0000000111001111100001",
			7373 => "0011000000101000000100",
			7374 => "0000001111001111100001",
			7375 => "0000000111001111100001",
			7376 => "0000000000111000000100",
			7377 => "0000000111001111100001",
			7378 => "0011111110000100000100",
			7379 => "1111111111001111100001",
			7380 => "0000000111001111100001",
			7381 => "0011011001001000000100",
			7382 => "0000001111001111100001",
			7383 => "1111111111001111100001",
			7384 => "0000000100010100011100",
			7385 => "0011110110110100001100",
			7386 => "0001000000010100000100",
			7387 => "0000000111001111100001",
			7388 => "0010110000101000000100",
			7389 => "0000001111001111100001",
			7390 => "0000010111001111100001",
			7391 => "0001000000010100001000",
			7392 => "0001000000010100000100",
			7393 => "0000000111001111100001",
			7394 => "0000001111001111100001",
			7395 => "0001111101100000000100",
			7396 => "0000000111001111100001",
			7397 => "0000001111001111100001",
			7398 => "0001000011010100001100",
			7399 => "0010000010101000000100",
			7400 => "1111111111001111100001",
			7401 => "0000001011000100000100",
			7402 => "0000001111001111100001",
			7403 => "1111111111001111100001",
			7404 => "0001110000101000001000",
			7405 => "0001000010100100000100",
			7406 => "0000000111001111100001",
			7407 => "0000000111001111100001",
			7408 => "0011011100110000000100",
			7409 => "0000010111001111100001",
			7410 => "0000000111001111100001",
			7411 => "0010100111110100001000",
			7412 => "0011001101010100000100",
			7413 => "0000001111001111100001",
			7414 => "0000000111001111100001",
			7415 => "1111111111001111100001",
			7416 => "0000100010110101010100",
			7417 => "0001100100110101001100",
			7418 => "0001100001111000100100",
			7419 => "0010001100000100010100",
			7420 => "0000101110101100010000",
			7421 => "0001011100110000001000",
			7422 => "0000001111000100000100",
			7423 => "0000001111010111111101",
			7424 => "0000000111010111111101",
			7425 => "0011110000011100000100",
			7426 => "0000000111010111111101",
			7427 => "0000001111010111111101",
			7428 => "0000001111010111111101",
			7429 => "0010110100010100001100",
			7430 => "0001110100010100001000",
			7431 => "0010111110111100000100",
			7432 => "0000001111010111111101",
			7433 => "1111111111010111111101",
			7434 => "0000001111010111111101",
			7435 => "1111111111010111111101",
			7436 => "0010110111111000010000",
			7437 => "0001101101111100001100",
			7438 => "0011110011100000001000",
			7439 => "0011001010000000000100",
			7440 => "0000000111010111111101",
			7441 => "0000001111010111111101",
			7442 => "1111111111010111111101",
			7443 => "1111111111010111111101",
			7444 => "0011000111111000001000",
			7445 => "0010000111000100000100",
			7446 => "0000000111010111111101",
			7447 => "0000001111010111111101",
			7448 => "0001010110000100001000",
			7449 => "0000010110000000000100",
			7450 => "0000000111010111111101",
			7451 => "0000001111010111111101",
			7452 => "0011000000101000000100",
			7453 => "0000000111010111111101",
			7454 => "0000001111010111111101",
			7455 => "0011111010111000000100",
			7456 => "0000000111010111111101",
			7457 => "1111111111010111111101",
			7458 => "0010011001111001101100",
			7459 => "0000111100001000111100",
			7460 => "0011110000011100011100",
			7461 => "0001000010111000001100",
			7462 => "0010011001111000001000",
			7463 => "0010001011010100000100",
			7464 => "0000000111010111111101",
			7465 => "1111111111010111111101",
			7466 => "1111111111010111111101",
			7467 => "0011100011111100001000",
			7468 => "0010000110001000000100",
			7469 => "0000001111010111111101",
			7470 => "0000000111010111111101",
			7471 => "0010000001110100000100",
			7472 => "0000000111010111111101",
			7473 => "0000001111010111111101",
			7474 => "0010110100010100010000",
			7475 => "0010110111111000001000",
			7476 => "0000010110000000000100",
			7477 => "0000000111010111111101",
			7478 => "1111111111010111111101",
			7479 => "0001110111111000000100",
			7480 => "0000001111010111111101",
			7481 => "0000000111010111111101",
			7482 => "0010010010001100001000",
			7483 => "0001101101111100000100",
			7484 => "0000000111010111111101",
			7485 => "0000001111010111111101",
			7486 => "0000000100010100000100",
			7487 => "1111111111010111111101",
			7488 => "1111111111010111111101",
			7489 => "0011110010001000011000",
			7490 => "0010001100000100001000",
			7491 => "0000111000111000000100",
			7492 => "1111111111010111111101",
			7493 => "0000000111010111111101",
			7494 => "0001001001000000001000",
			7495 => "0001000011101100000100",
			7496 => "0000000111010111111101",
			7497 => "0000001111010111111101",
			7498 => "0000110100000000000100",
			7499 => "0000000111010111111101",
			7500 => "1111111111010111111101",
			7501 => "0010000010101000010000",
			7502 => "0010000001110100001000",
			7503 => "0001001010110100000100",
			7504 => "0000001111010111111101",
			7505 => "0000000111010111111101",
			7506 => "0001110100010100000100",
			7507 => "0000001111010111111101",
			7508 => "0000000111010111111101",
			7509 => "0001110000101000000100",
			7510 => "1111111111010111111101",
			7511 => "0000000111010111111101",
			7512 => "0000011110100000101100",
			7513 => "0001010011011100001100",
			7514 => "0011000111111000000100",
			7515 => "0000000111010111111101",
			7516 => "0010011001111000000100",
			7517 => "0000001111010111111101",
			7518 => "0000000111010111111101",
			7519 => "0011000111111000010000",
			7520 => "0000100001000000001000",
			7521 => "0001000110001100000100",
			7522 => "0000000111010111111101",
			7523 => "0000001111010111111101",
			7524 => "0000111001110000000100",
			7525 => "1111111111010111111101",
			7526 => "0000000111010111111101",
			7527 => "0011000100010100001000",
			7528 => "0000000100000000000100",
			7529 => "0000000111010111111101",
			7530 => "0000000111010111111101",
			7531 => "0011000000101000000100",
			7532 => "0000000111010111111101",
			7533 => "0000000111010111111101",
			7534 => "0000111100001000000100",
			7535 => "0000001111010111111101",
			7536 => "0011000111111000010000",
			7537 => "0001010101101100001000",
			7538 => "0001011101100000000100",
			7539 => "0000000111010111111101",
			7540 => "1111111111010111111101",
			7541 => "0010001100000100000100",
			7542 => "1111111111010111111101",
			7543 => "0000000111010111111101",
			7544 => "0010111100001000001000",
			7545 => "0001111100001000000100",
			7546 => "0000000111010111111101",
			7547 => "0000001111010111111101",
			7548 => "0000111001110000000100",
			7549 => "1111111111010111111101",
			7550 => "0000000111010111111101",
			7551 => "0010000111000011001000",
			7552 => "0001101101011001110100",
			7553 => "0011000000101000111000",
			7554 => "0011000100010100100000",
			7555 => "0011000100010100010000",
			7556 => "0001111100001000001000",
			7557 => "0001111100001000000100",
			7558 => "0000000111100000011001",
			7559 => "1111111111100000011001",
			7560 => "0000101100010100000100",
			7561 => "0000001111100000011001",
			7562 => "0000000111100000011001",
			7563 => "0011000100010100001000",
			7564 => "0001001011110000000100",
			7565 => "1111111111100000011001",
			7566 => "0000000111100000011001",
			7567 => "0011011100101100000100",
			7568 => "0000000111100000011001",
			7569 => "0000000111100000011001",
			7570 => "0001110000101000001100",
			7571 => "0001001001001100001000",
			7572 => "0001110000101000000100",
			7573 => "0000000111100000011001",
			7574 => "0000001111100000011001",
			7575 => "0000001111100000011001",
			7576 => "0011101100101100001000",
			7577 => "0000100101110000000100",
			7578 => "0000000111100000011001",
			7579 => "0000000111100000011001",
			7580 => "0000001111100000011001",
			7581 => "0011000000101000011100",
			7582 => "0000101110000100001100",
			7583 => "0000011100110100001000",
			7584 => "0001111100001000000100",
			7585 => "0000000111100000011001",
			7586 => "1111111111100000011001",
			7587 => "0000001111100000011001",
			7588 => "0010101000010100001000",
			7589 => "0000010010001100000100",
			7590 => "1111110111100000011001",
			7591 => "1111111111100000011001",
			7592 => "0001000011001100000100",
			7593 => "0000000111100000011001",
			7594 => "1111111111100000011001",
			7595 => "0011000000101000010000",
			7596 => "0011101101111000001000",
			7597 => "0011011100101000000100",
			7598 => "0000000111100000011001",
			7599 => "0000000111100000011001",
			7600 => "0011010001111100000100",
			7601 => "0000000111100000011001",
			7602 => "0000001111100000011001",
			7603 => "0011000000101000001000",
			7604 => "0001100001111000000100",
			7605 => "1111111111100000011001",
			7606 => "0000000111100000011001",
			7607 => "0011000000101000000100",
			7608 => "0000000111100000011001",
			7609 => "0000000111100000011001",
			7610 => "0001111000111000100000",
			7611 => "0011011100101000001100",
			7612 => "0001000100001100001000",
			7613 => "0000110100001000000100",
			7614 => "0000000111100000011001",
			7615 => "0000001111100000011001",
			7616 => "1111111111100000011001",
			7617 => "0010011101101000001000",
			7618 => "0010111000111100000100",
			7619 => "0000000111100000011001",
			7620 => "0000001111100000011001",
			7621 => "0000010010001100000100",
			7622 => "1111111111100000011001",
			7623 => "0011101010111100000100",
			7624 => "0000000111100000011001",
			7625 => "0000001111100000011001",
			7626 => "0000100010000000010100",
			7627 => "0000000000111000001100",
			7628 => "0000111010011100000100",
			7629 => "0000001111100000011001",
			7630 => "0000110000011100000100",
			7631 => "1111111111100000011001",
			7632 => "0000000111100000011001",
			7633 => "0000101100010100000100",
			7634 => "1111111111100000011001",
			7635 => "1111111111100000011001",
			7636 => "0001101011001100010000",
			7637 => "0011001000111000001000",
			7638 => "0010111101100000000100",
			7639 => "0000000111100000011001",
			7640 => "0000001111100000011001",
			7641 => "0011100110100100000100",
			7642 => "1111111111100000011001",
			7643 => "0000000111100000011001",
			7644 => "0000111111011100001000",
			7645 => "0000001011000100000100",
			7646 => "1111111111100000011001",
			7647 => "0000000111100000011001",
			7648 => "0000110100000100000100",
			7649 => "0000001111100000011001",
			7650 => "0000000111100000011001",
			7651 => "0000101100000001000100",
			7652 => "0000101001100000110100",
			7653 => "0011000111111000011000",
			7654 => "0010110100010100010000",
			7655 => "0010011100110100001000",
			7656 => "0000111000110000000100",
			7657 => "1111111111100000011001",
			7658 => "0000001111100000011001",
			7659 => "0011101000110000000100",
			7660 => "0000000111100000011001",
			7661 => "1111111111100000011001",
			7662 => "0011010011011100000100",
			7663 => "1111111111100000011001",
			7664 => "0000010111100000011001",
			7665 => "0001111011000100010000",
			7666 => "0001000010010000001000",
			7667 => "0011011001110000000100",
			7668 => "0000000111100000011001",
			7669 => "1111111111100000011001",
			7670 => "0001100100110100000100",
			7671 => "0000000111100000011001",
			7672 => "0000000111100000011001",
			7673 => "0001111100001000001000",
			7674 => "0010001000110000000100",
			7675 => "0000000111100000011001",
			7676 => "0000000111100000011001",
			7677 => "1111111111100000011001",
			7678 => "0010100101000100000100",
			7679 => "1111111111100000011001",
			7680 => "0011101100001000001000",
			7681 => "0000101100000000000100",
			7682 => "0000000111100000011001",
			7683 => "0000000111100000011001",
			7684 => "0000001111100000011001",
			7685 => "1111111111100000011001",
			7686 => "0011100101101111001000",
			7687 => "0011000100010101011100",
			7688 => "0011000100010101000000",
			7689 => "0001001101001000100000",
			7690 => "0000000011010000010000",
			7691 => "0001001000001000001000",
			7692 => "0000100101110000000100",
			7693 => "0000000111101010100101",
			7694 => "1111111111101010100101",
			7695 => "0011100100010100000100",
			7696 => "0000001111101010100101",
			7697 => "0000000111101010100101",
			7698 => "0011101011000100001000",
			7699 => "0010001011010100000100",
			7700 => "1111111111101010100101",
			7701 => "0000000111101010100101",
			7702 => "0010100001010000000100",
			7703 => "1111111111101010100101",
			7704 => "0000000111101010100101",
			7705 => "0000100010000000010000",
			7706 => "0000000100010100001000",
			7707 => "0010000001110100000100",
			7708 => "0000000111101010100101",
			7709 => "0000001111101010100101",
			7710 => "0010101010110000000100",
			7711 => "1111111111101010100101",
			7712 => "0000000111101010100101",
			7713 => "0011001110111100001000",
			7714 => "0001001011100000000100",
			7715 => "0000001111101010100101",
			7716 => "1111111111101010100101",
			7717 => "0001011100101100000100",
			7718 => "1111111111101010100101",
			7719 => "0000000111101010100101",
			7720 => "0010111011000100001000",
			7721 => "0000000111111000000100",
			7722 => "1111111111101010100101",
			7723 => "0000000111101010100101",
			7724 => "0010001100000100000100",
			7725 => "0000010111101010100101",
			7726 => "0001100100110100001000",
			7727 => "0001010101101100000100",
			7728 => "0000001111101010100101",
			7729 => "0000000111101010100101",
			7730 => "0001101100011000000100",
			7731 => "0000010111101010100101",
			7732 => "0000000111101010100101",
			7733 => "0011000100010100101100",
			7734 => "0010100110011100011100",
			7735 => "0000101110000100010000",
			7736 => "0011100000101000001000",
			7737 => "0010101001000100000100",
			7738 => "1111111111101010100101",
			7739 => "0000000111101010100101",
			7740 => "0010000001110000000100",
			7741 => "0000000111101010100101",
			7742 => "0000001111101010100101",
			7743 => "0011011101100000000100",
			7744 => "0000000111101010100101",
			7745 => "0000111101111000000100",
			7746 => "1111111111101010100101",
			7747 => "0000000111101010100101",
			7748 => "0001111100001000001100",
			7749 => "0010111100001000001000",
			7750 => "0010100101000100000100",
			7751 => "0000001111101010100101",
			7752 => "0000000111101010100101",
			7753 => "1111111111101010100101",
			7754 => "0000001111101010100101",
			7755 => "0010111100001000100000",
			7756 => "0010110000101000010000",
			7757 => "0001010101101100001000",
			7758 => "0000011110100000000100",
			7759 => "0000000111101010100101",
			7760 => "0000000111101010100101",
			7761 => "0011100000101000000100",
			7762 => "1111111111101010100101",
			7763 => "0000000111101010100101",
			7764 => "0011000100010100001000",
			7765 => "0001110000101000000100",
			7766 => "0000001111101010100101",
			7767 => "0000010111101010100101",
			7768 => "0000111101100000000100",
			7769 => "0000000111101010100101",
			7770 => "0000001111101010100101",
			7771 => "0010111100001000010000",
			7772 => "0001010110000100001000",
			7773 => "0001101101111100000100",
			7774 => "0000001111101010100101",
			7775 => "1111111111101010100101",
			7776 => "0011000000101000000100",
			7777 => "1111111111101010100101",
			7778 => "0000000111101010100101",
			7779 => "0000100101110000001000",
			7780 => "0011010001111100000100",
			7781 => "0000000111101010100101",
			7782 => "1111111111101010100101",
			7783 => "0010001011010100000100",
			7784 => "1111111111101010100101",
			7785 => "0000000111101010100101",
			7786 => "0000001111000101001000",
			7787 => "0001001000000100101100",
			7788 => "0000001101010000011000",
			7789 => "0001001011110000010000",
			7790 => "0001101010011000001000",
			7791 => "0010100111110100000100",
			7792 => "0000000111101010100101",
			7793 => "0000000111101010100101",
			7794 => "0001001000101000000100",
			7795 => "1111111111101010100101",
			7796 => "0000000111101010100101",
			7797 => "0000000111000100000100",
			7798 => "0000000111101010100101",
			7799 => "1111111111101010100101",
			7800 => "0011000000101000001000",
			7801 => "0010101000010100000100",
			7802 => "0000001111101010100101",
			7803 => "1111111111101010100101",
			7804 => "0010111110001100001000",
			7805 => "0000010111100100000100",
			7806 => "0000001111101010100101",
			7807 => "0000000111101010100101",
			7808 => "0000000111101010100101",
			7809 => "0000101100010100001100",
			7810 => "0000100100101000000100",
			7811 => "0000000111101010100101",
			7812 => "0010001100000100000100",
			7813 => "1111111111101010100101",
			7814 => "1111110111101010100101",
			7815 => "0001000110001100001100",
			7816 => "0010001001101000001000",
			7817 => "0000001101010000000100",
			7818 => "0000000111101010100101",
			7819 => "0000001111101010100101",
			7820 => "1111111111101010100101",
			7821 => "1111111111101010100101",
			7822 => "0010001001101000010100",
			7823 => "0001000110001100001100",
			7824 => "0000010010001100001000",
			7825 => "0010101000010100000100",
			7826 => "0000000111101010100101",
			7827 => "0000001111101010100101",
			7828 => "0000001111101010100101",
			7829 => "0000000010111100000100",
			7830 => "1111111111101010100101",
			7831 => "0000001111101010100101",
			7832 => "0000110000001100000100",
			7833 => "1111111111101010100101",
			7834 => "0000101110010000010000",
			7835 => "0001101010011000001000",
			7836 => "0011010001111100000100",
			7837 => "0000000111101010100101",
			7838 => "0000001111101010100101",
			7839 => "0011000100000000000100",
			7840 => "0000000111101010100101",
			7841 => "1111111111101010100101",
			7842 => "0001101100011000001000",
			7843 => "0001011100101100000100",
			7844 => "0000000111101010100101",
			7845 => "0000000111101010100101",
			7846 => "0001010100001000000100",
			7847 => "0000000111101010100101",
			7848 => "0000000111101010100101",
			7849 => "0011000100001010111000",
			7850 => "0011110010001001011000",
			7851 => "0000110100000000100000",
			7852 => "0001111100001000011100",
			7853 => "0000011110100000010000",
			7854 => "0010010010001100001000",
			7855 => "0000110100010100000100",
			7856 => "0000000111110000011001",
			7857 => "0000000111110000011001",
			7858 => "0000101110101000000100",
			7859 => "0000000111110000011001",
			7860 => "0000000111110000011001",
			7861 => "0000110000101000000100",
			7862 => "0000011111110000011001",
			7863 => "0010010110101000000100",
			7864 => "1111111111110000011001",
			7865 => "0000000111110000011001",
			7866 => "1111111111110000011001",
			7867 => "0010010110101000011100",
			7868 => "0000111101100000010000",
			7869 => "0011110001011000001000",
			7870 => "0000111000111000000100",
			7871 => "0000000111110000011001",
			7872 => "0000001111110000011001",
			7873 => "0000101001010000000100",
			7874 => "0000000111110000011001",
			7875 => "0000000111110000011001",
			7876 => "0000011110100000000100",
			7877 => "1111110111110000011001",
			7878 => "0010010110101000000100",
			7879 => "0000001111110000011001",
			7880 => "0000001111110000011001",
			7881 => "0000011110100000001100",
			7882 => "0011111011011100001000",
			7883 => "0011110000011100000100",
			7884 => "1111111111110000011001",
			7885 => "1111111111110000011001",
			7886 => "0000000111110000011001",
			7887 => "0001100001111000001000",
			7888 => "0001011110001100000100",
			7889 => "0000000111110000011001",
			7890 => "1111111111110000011001",
			7891 => "0000001011000100000100",
			7892 => "0000000111110000011001",
			7893 => "1111111111110000011001",
			7894 => "0000110101101100100000",
			7895 => "0000110101101100011000",
			7896 => "0000111100110000010000",
			7897 => "0001111011000100001000",
			7898 => "0010100110011000000100",
			7899 => "1111111111110000011001",
			7900 => "0000000111110000011001",
			7901 => "0011000111111000000100",
			7902 => "1111111111110000011001",
			7903 => "0000000111110000011001",
			7904 => "0011000100010100000100",
			7905 => "0000001111110000011001",
			7906 => "0000000111110000011001",
			7907 => "0011110101110100000100",
			7908 => "1111111111110000011001",
			7909 => "1111111111110000011001",
			7910 => "0010000010101000100000",
			7911 => "0010010110101000010000",
			7912 => "0011110111110000001000",
			7913 => "0001110100010100000100",
			7914 => "0000000111110000011001",
			7915 => "0000010111110000011001",
			7916 => "0001100100110100000100",
			7917 => "1111111111110000011001",
			7918 => "0000001111110000011001",
			7919 => "0000111100101100001000",
			7920 => "0010010111100100000100",
			7921 => "0000000111110000011001",
			7922 => "1111111111110000011001",
			7923 => "0010010111100100000100",
			7924 => "0000000111110000011001",
			7925 => "0000000111110000011001",
			7926 => "0010100110011100010000",
			7927 => "0011000000101000001000",
			7928 => "0011110001001000000100",
			7929 => "0000011111110000011001",
			7930 => "0000001111110000011001",
			7931 => "0001000011101100000100",
			7932 => "0000001111110000011001",
			7933 => "1111111111110000011001",
			7934 => "0000001011000100001000",
			7935 => "0001000010100100000100",
			7936 => "0000001111110000011001",
			7937 => "1111111111110000011001",
			7938 => "0001110000101000000100",
			7939 => "0000001111110000011001",
			7940 => "0000000111110000011001",
			7941 => "1111111111110000011001",
			7942 => "0000101100010110110100",
			7943 => "0001101101011010000000",
			7944 => "0001101100011001000000",
			7945 => "0000100111111100100000",
			7946 => "0000100111111100010000",
			7947 => "0000100100101000001000",
			7948 => "0001101101111100000100",
			7949 => "0000000111111100000111",
			7950 => "0000000111111100000111",
			7951 => "0011110010001000000100",
			7952 => "0000001111111100000111",
			7953 => "1111111111111100000111",
			7954 => "0000011100110100001000",
			7955 => "0011011100110000000100",
			7956 => "0000010111111100000111",
			7957 => "1111111111111100000111",
			7958 => "0000011100110100000100",
			7959 => "0000001111111100000111",
			7960 => "0000000111111100000111",
			7961 => "0001010000001100010000",
			7962 => "0000101100010100001000",
			7963 => "0011101011000100000100",
			7964 => "0000000111111100000111",
			7965 => "0000000111111100000111",
			7966 => "0010101010110000000100",
			7967 => "0000000111111100000111",
			7968 => "0000001111111100000111",
			7969 => "0011100101101100001000",
			7970 => "0010010111100100000100",
			7971 => "0000001111111100000111",
			7972 => "1111111111111100000111",
			7973 => "0000100011001000000100",
			7974 => "0000000111111100000111",
			7975 => "1111111111111100000111",
			7976 => "0001101100011000100000",
			7977 => "0011101001110000010000",
			7978 => "0010000001110100001000",
			7979 => "0000000111111000000100",
			7980 => "0000000111111100000111",
			7981 => "1111111111111100000111",
			7982 => "0000000100010100000100",
			7983 => "0000010111111100000111",
			7984 => "0000000111111100000111",
			7985 => "0010011011101000001000",
			7986 => "0010100001010000000100",
			7987 => "0000001111111100000111",
			7988 => "0000001111111100000111",
			7989 => "0011110010110100000100",
			7990 => "0000000111111100000111",
			7991 => "0000001111111100000111",
			7992 => "0011000100000000010000",
			7993 => "0011101110001100001000",
			7994 => "0010010111100100000100",
			7995 => "0000000111111100000111",
			7996 => "0000000111111100000111",
			7997 => "0001101010011000000100",
			7998 => "0000001111111100000111",
			7999 => "0000000111111100000111",
			8000 => "0011001001110000001000",
			8001 => "0011110000110100000100",
			8002 => "1111111111111100000111",
			8003 => "0000000111111100000111",
			8004 => "0010111100101100000100",
			8005 => "0000010111111100000111",
			8006 => "0000000111111100000111",
			8007 => "0001010011100000100000",
			8008 => "0001101101011000010000",
			8009 => "0000101100010100001100",
			8010 => "0000100010011100000100",
			8011 => "0000000111111100000111",
			8012 => "0011100110000100000100",
			8013 => "1111111111111100000111",
			8014 => "1111111111111100000111",
			8015 => "0000000111111100000111",
			8016 => "0000000011111100000100",
			8017 => "1111111111111100000111",
			8018 => "0000001110111100000100",
			8019 => "0000001111111100000111",
			8020 => "0010111001110000000100",
			8021 => "0000000111111100000111",
			8022 => "1111111111111100000111",
			8023 => "0011010110100100001000",
			8024 => "0011000110000100000100",
			8025 => "0000010111111100000111",
			8026 => "0000000111111100000111",
			8027 => "0011011000011000000100",
			8028 => "0000000111111100000111",
			8029 => "0001011000011000000100",
			8030 => "0000001111111100000111",
			8031 => "0000000111111100000111",
			8032 => "0001101100011001011000",
			8033 => "0011000111111000100100",
			8034 => "0010101010110000010000",
			8035 => "0000100110010000001000",
			8036 => "0010001111001000000100",
			8037 => "0000000111111100000111",
			8038 => "0000001111111100000111",
			8039 => "0001000011010100000100",
			8040 => "0000001111111100000111",
			8041 => "1111111111111100000111",
			8042 => "0000101110110100001100",
			8043 => "0010110100010100001000",
			8044 => "0000100010000000000100",
			8045 => "0000001111111100000111",
			8046 => "1111111111111100000111",
			8047 => "1111111111111100000111",
			8048 => "0011001010000000000100",
			8049 => "0000000111111100000111",
			8050 => "0000001111111100000111",
			8051 => "0001010100001000011000",
			8052 => "0010011101101000010000",
			8053 => "0010010111100100001000",
			8054 => "0001011110001100000100",
			8055 => "0000000111111100000111",
			8056 => "0000001111111100000111",
			8057 => "0011101110001100000100",
			8058 => "1111111111111100000111",
			8059 => "0000000111111100000111",
			8060 => "0001101100011000000100",
			8061 => "1111111111111100000111",
			8062 => "1111110111111100000111",
			8063 => "0001101100011000001100",
			8064 => "0000010111100100000100",
			8065 => "1111111111111100000111",
			8066 => "0011100011001000000100",
			8067 => "0000000111111100000111",
			8068 => "0000000111111100000111",
			8069 => "0011110001000000001000",
			8070 => "0001000000010100000100",
			8071 => "0000001111111100000111",
			8072 => "1111111111111100000111",
			8073 => "0000101001100000000100",
			8074 => "1111111111111100000111",
			8075 => "0000000111111100000111",
			8076 => "0010011011101001000000",
			8077 => "0001000100001100100000",
			8078 => "0001011010111100010000",
			8079 => "0010011101101000001000",
			8080 => "0001011101111000000100",
			8081 => "0000000111111100000111",
			8082 => "0000001111111100000111",
			8083 => "0000010010001100000100",
			8084 => "1111111111111100000111",
			8085 => "0000000111111100000111",
			8086 => "0011111101000100001000",
			8087 => "0011000100000000000100",
			8088 => "0000001111111100000111",
			8089 => "0000000111111100000111",
			8090 => "0011101101010100000100",
			8091 => "0000010111111100000111",
			8092 => "0000001111111100000111",
			8093 => "0010111100001000010000",
			8094 => "0010100110011100001000",
			8095 => "0011101000111000000100",
			8096 => "0000000111111100000111",
			8097 => "0000010111111100000111",
			8098 => "0011110010110100000100",
			8099 => "0000001111111100000111",
			8100 => "1111111111111100000111",
			8101 => "0010111000111100001000",
			8102 => "0010010110101000000100",
			8103 => "0000000111111100000111",
			8104 => "1111111111111100000111",
			8105 => "0001101101011000000100",
			8106 => "1111111111111100000111",
			8107 => "0000000111111100000111",
			8108 => "0011000100000000010100",
			8109 => "0001101101011000000100",
			8110 => "1111111111111100000111",
			8111 => "0001001110111000001000",
			8112 => "0010011111001100000100",
			8113 => "0000001111111100000111",
			8114 => "1111111111111100000111",
			8115 => "0010100101000100000100",
			8116 => "1111111111111100000111",
			8117 => "0000000111111100000111",
			8118 => "0011000100000000001000",
			8119 => "0001101111000000000100",
			8120 => "0000001111111100000111",
			8121 => "1111111111111100000111",
			8122 => "0011111101000100001000",
			8123 => "0001101001100100000100",
			8124 => "1111111111111100000111",
			8125 => "0000001111111100000111",
			8126 => "0001101011001100000100",
			8127 => "0000000111111100000111",
			8128 => "0000000111111100000111",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(2792, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(5598, initial_addr_3'length));
	end generate gen_rom_14;

	gen_rom_15: if SELECT_ROM = 15 generate
		bank <= (
			0 => "0000000000000000000101",
			1 => "0000000000000000001001",
			2 => "0000000000000000001101",
			3 => "0000000000000000010001",
			4 => "0000000000000000010101",
			5 => "0000000000000000011001",
			6 => "0000000000000000011101",
			7 => "0000000000000000100001",
			8 => "0000000000000000100101",
			9 => "0000000000000000101001",
			10 => "0000000000000000101101",
			11 => "0000000000000000110001",
			12 => "0000000000000000110101",
			13 => "0000000000000000111001",
			14 => "0000000000000000111101",
			15 => "0000000000000001000001",
			16 => "0000000000000001000101",
			17 => "0000000000000001001001",
			18 => "0000000000000001001101",
			19 => "0010111101010100000100",
			20 => "0000000000000001011001",
			21 => "0000000000000001011001",
			22 => "0001111110001100000100",
			23 => "0000000000000001100101",
			24 => "0000000000000001100101",
			25 => "0011001010000000000100",
			26 => "0000000000000001110001",
			27 => "0000000000000001110001",
			28 => "0011001010000000000100",
			29 => "0000000000000010000101",
			30 => "0010100000001000000100",
			31 => "0000000000000010000101",
			32 => "0000000000000010000101",
			33 => "0001111110001100001000",
			34 => "0010110000111000000100",
			35 => "0000000000000010011001",
			36 => "0000000000000010011001",
			37 => "0000000000000010011001",
			38 => "0001100001000100000100",
			39 => "0000000000000010101101",
			40 => "0001101010011000000100",
			41 => "0000000000000010101101",
			42 => "0000000000000010101101",
			43 => "0001101101111100001000",
			44 => "0001101101011100000100",
			45 => "0000000000000011000001",
			46 => "0000000000000011000001",
			47 => "0000000000000011000001",
			48 => "0000011110100000001000",
			49 => "0010011100100000000100",
			50 => "0000000000000011010101",
			51 => "0000000000000011010101",
			52 => "0000000000000011010101",
			53 => "0001101110010100000100",
			54 => "0000000000000011101001",
			55 => "0001101111000000000100",
			56 => "0000000000000011101001",
			57 => "0000000000000011101001",
			58 => "0001100001111000000100",
			59 => "0000000000000100000101",
			60 => "0001101010011000001000",
			61 => "0001001101000000000100",
			62 => "0000000000000100000101",
			63 => "0000000000000100000101",
			64 => "0000000000000100000101",
			65 => "0001111110001100001100",
			66 => "0011111001001000000100",
			67 => "0000000000000100100001",
			68 => "0011001100110000000100",
			69 => "0000000000000100100001",
			70 => "0000000000000100100001",
			71 => "0000000000000100100001",
			72 => "0001100001111000001100",
			73 => "0001101101011100000100",
			74 => "0000000000000100111101",
			75 => "0001101011111100000100",
			76 => "0000000000000100111101",
			77 => "0000000000000100111101",
			78 => "0000000000000100111101",
			79 => "0001111110001100001100",
			80 => "0011110100011000000100",
			81 => "0000000000000101011001",
			82 => "0000011011101000000100",
			83 => "0000000000000101011001",
			84 => "0000000000000101011001",
			85 => "0000000000000101011001",
			86 => "0001101101111100001100",
			87 => "0010101001100100000100",
			88 => "0000000000000101111101",
			89 => "0010100011101000000100",
			90 => "0000000000000101111101",
			91 => "0000000000000101111101",
			92 => "0001101001100100000100",
			93 => "0000000000000101111101",
			94 => "0000000000000101111101",
			95 => "0000010110000000001100",
			96 => "0000011110011100000100",
			97 => "0000000000000110100001",
			98 => "0000101010010100000100",
			99 => "0000000000000110100001",
			100 => "0000000000000110100001",
			101 => "0000101100010100000100",
			102 => "0000000000000110100001",
			103 => "0000000000000110100001",
			104 => "0000010000011000001100",
			105 => "0011000111111000001000",
			106 => "0011111010111100000100",
			107 => "0000000000000111001101",
			108 => "0000000000000111001101",
			109 => "0000000000000111001101",
			110 => "0000001001101000000100",
			111 => "0000000000000111001101",
			112 => "0001101011111100000100",
			113 => "0000000000000111001101",
			114 => "0000000000000111001101",
			115 => "0001111110001100010000",
			116 => "0010101000100100001100",
			117 => "0011010100000000000100",
			118 => "0000000000000111110001",
			119 => "0010000000001000000100",
			120 => "0000000000000111110001",
			121 => "0000000000000111110001",
			122 => "0000000000000111110001",
			123 => "0000000000000111110001",
			124 => "0001100001000100000100",
			125 => "0000000000001000010101",
			126 => "0011000000110000000100",
			127 => "0000000000001000010101",
			128 => "0011001110001100001000",
			129 => "0001101101111100000100",
			130 => "0000000000001000010101",
			131 => "0000000000001000010101",
			132 => "0000000000001000010101",
			133 => "0010111010111000010000",
			134 => "0011111110110000000100",
			135 => "0000000000001000111001",
			136 => "0011001100110000001000",
			137 => "0001111110001100000100",
			138 => "0000000000001000111001",
			139 => "0000000000001000111001",
			140 => "0000000000001000111001",
			141 => "0000000000001000111001",
			142 => "0001111110001100010000",
			143 => "0011111010111100000100",
			144 => "0000000000001001011101",
			145 => "0010101001100100000100",
			146 => "0000000000001001011101",
			147 => "0011001100110000000100",
			148 => "0000000000001001011101",
			149 => "0000000000001001011101",
			150 => "0000000000001001011101",
			151 => "0011111010111100000100",
			152 => "0000000000001010000001",
			153 => "0011000100001000001100",
			154 => "0011111100111000001000",
			155 => "0001111110110000000100",
			156 => "0000000000001010000001",
			157 => "0000000000001010000001",
			158 => "0000000000001010000001",
			159 => "0000000000001010000001",
			160 => "0001110110000100010000",
			161 => "0001101101111100001100",
			162 => "0001101001011000000100",
			163 => "0000000000001010101101",
			164 => "0010110000111000000100",
			165 => "0000000000001010101101",
			166 => "0000000000001010101101",
			167 => "0000000000001010101101",
			168 => "0010111001110100000100",
			169 => "0000000000001010101101",
			170 => "0000000000001010101101",
			171 => "0000101110010000001100",
			172 => "0000010000011000000100",
			173 => "0000000000001011100001",
			174 => "0011000000111000000100",
			175 => "0000000000001011100001",
			176 => "0000000000001011100001",
			177 => "0001111110001100001100",
			178 => "0000011011101000001000",
			179 => "0011000011011100000100",
			180 => "0000000000001011100001",
			181 => "0000000000001011100001",
			182 => "0000000000001011100001",
			183 => "0000000000001011100001",
			184 => "0000011110100000010000",
			185 => "0010011100100000000100",
			186 => "0000000000001100010101",
			187 => "0001010100000000000100",
			188 => "0000000000001100010101",
			189 => "0001110000101000000100",
			190 => "0000000000001100010101",
			191 => "0000000000001100010101",
			192 => "0001101010011000001000",
			193 => "0000011110100000000100",
			194 => "0000000000001100010101",
			195 => "0000000000001100010101",
			196 => "0000000000001100010101",
			197 => "0001111110001100011000",
			198 => "0011110101100100001100",
			199 => "0001100001000100000100",
			200 => "0000000000001101010001",
			201 => "0000011100100000000100",
			202 => "0000000000001101010001",
			203 => "0000000000001101010001",
			204 => "0000011011101000001000",
			205 => "0010101000100100000100",
			206 => "0000000000001101010001",
			207 => "0000000000001101010001",
			208 => "0000000000001101010001",
			209 => "0001101001100100000100",
			210 => "0000000000001101010001",
			211 => "0000000000001101010001",
			212 => "0001111110001100010100",
			213 => "0011111010111100000100",
			214 => "0000000000001101111101",
			215 => "0010101001100100000100",
			216 => "0000000000001101111101",
			217 => "0011001100110000001000",
			218 => "0010110000111000000100",
			219 => "0000000000001101111101",
			220 => "0000000000001101111101",
			221 => "0000000000001101111101",
			222 => "0000000000001101111101",
			223 => "0011001010000000000100",
			224 => "0000000000001110101001",
			225 => "0001100101011100000100",
			226 => "0000000000001110101001",
			227 => "0001101001100100001100",
			228 => "0001111010000000000100",
			229 => "0000000000001110101001",
			230 => "0001101011111100000100",
			231 => "0000000000001110101001",
			232 => "0000000000001110101001",
			233 => "0000000000001110101001",
			234 => "0011001010000000010100",
			235 => "0000100001001000000100",
			236 => "0000000000001111100101",
			237 => "0000011110100000001100",
			238 => "0010011100100000000100",
			239 => "0000000000001111100101",
			240 => "0010110000111000000100",
			241 => "0000000000001111100101",
			242 => "0000000000001111100101",
			243 => "0000000000001111100101",
			244 => "0001101010011000001000",
			245 => "0001100001111000000100",
			246 => "0000000000001111100101",
			247 => "0000000000001111100101",
			248 => "0000000000001111100101",
			249 => "0011001010000000010100",
			250 => "0000011110100000010000",
			251 => "0011010000101000000100",
			252 => "0000000000010000100001",
			253 => "0010011100100000000100",
			254 => "0000000000010000100001",
			255 => "0001110100010100000100",
			256 => "0000000000010000100001",
			257 => "0000000000010000100001",
			258 => "0000000000010000100001",
			259 => "0001110111001000001000",
			260 => "0000011110100000000100",
			261 => "0000000000010000100001",
			262 => "0000000000010000100001",
			263 => "0000000000010000100001",
			264 => "0000010110000000010000",
			265 => "0011000100000000001100",
			266 => "0010011100100000000100",
			267 => "0000000000010001100101",
			268 => "0000011110011100000100",
			269 => "0000000000010001100101",
			270 => "0000000000010001100101",
			271 => "0000000000010001100101",
			272 => "0011001100110000010000",
			273 => "0001101010011000001100",
			274 => "0011001010000000000100",
			275 => "0000000000010001100101",
			276 => "0001101001011000000100",
			277 => "0000000000010001100101",
			278 => "0000000000010001100101",
			279 => "0000000000010001100101",
			280 => "0000000000010001100101",
			281 => "0010010010001100001100",
			282 => "0000111010101100000100",
			283 => "0000000000010010110001",
			284 => "0001111100001000000100",
			285 => "0000000000010010110001",
			286 => "0000000000010010110001",
			287 => "0011100101001000010000",
			288 => "0010100000001000000100",
			289 => "0000000000010010110001",
			290 => "0011000000111000000100",
			291 => "0000000000010010110001",
			292 => "0001101011111100000100",
			293 => "0000000000010010110001",
			294 => "0000000000010010110001",
			295 => "0011101001010000000100",
			296 => "0000000000010010110001",
			297 => "0000101100111000000100",
			298 => "0000000000010010110001",
			299 => "0000000000010010110001",
			300 => "0011001010000000010100",
			301 => "0000101010010100000100",
			302 => "0000000000010011111101",
			303 => "0010111011000100001100",
			304 => "0010110000111000000100",
			305 => "0000000000010011111101",
			306 => "0001110100010100000100",
			307 => "0000000000010011111101",
			308 => "0000000000010011111101",
			309 => "0000000000010011111101",
			310 => "0000101100010100001000",
			311 => "0001111010000000000100",
			312 => "0000000000010011111101",
			313 => "0000000000010011111101",
			314 => "0001111110001100001000",
			315 => "0001110101101100000100",
			316 => "0000000000010011111101",
			317 => "0000000000010011111101",
			318 => "0000000000010011111101",
			319 => "0010000101000100011000",
			320 => "0011100010111100000100",
			321 => "0000000000010101001001",
			322 => "0011101001010000001100",
			323 => "0010100011101000001000",
			324 => "0000001010110000000100",
			325 => "0000000000010101001001",
			326 => "0000000000010101001001",
			327 => "0000000000010101001001",
			328 => "0010001010110000000100",
			329 => "0000000000010101001001",
			330 => "0000000000010101001001",
			331 => "0011100111010100001100",
			332 => "0011101000110000000100",
			333 => "0000000000010101001001",
			334 => "0010100111110100000100",
			335 => "0000000000010101001001",
			336 => "0000000000010101001001",
			337 => "0000000000010101001001",
			338 => "0000011110100000011000",
			339 => "0000100100101000010000",
			340 => "0001100001000100001000",
			341 => "0000110000111000000100",
			342 => "0000000000010110100101",
			343 => "0000000000010110100101",
			344 => "0011101110111100000100",
			345 => "0000000000010110100101",
			346 => "0000000000010110100101",
			347 => "0011000100010100000100",
			348 => "0000000000010110100101",
			349 => "0000000000010110100101",
			350 => "0011010010001000001000",
			351 => "0010100111101100000100",
			352 => "0000000000010110100101",
			353 => "1111111000010110100101",
			354 => "0010011011001100001100",
			355 => "0011000100001000001000",
			356 => "0011011110101100000100",
			357 => "0000000000010110100101",
			358 => "0000000000010110100101",
			359 => "0000000000010110100101",
			360 => "0000000000010110100101",
			361 => "0000010000011000010100",
			362 => "0011000111111000010000",
			363 => "0010011100100000000100",
			364 => "0000000000010111110001",
			365 => "0010110000111000000100",
			366 => "0000000000010111110001",
			367 => "0000011110011100000100",
			368 => "0000000000010111110001",
			369 => "0000000000010111110001",
			370 => "0000000000010111110001",
			371 => "0000101011111000010000",
			372 => "0011001100110000001100",
			373 => "0010001001000100000100",
			374 => "0000000000010111110001",
			375 => "0011000000111000000100",
			376 => "0000000000010111110001",
			377 => "0000000000010111110001",
			378 => "0000000000010111110001",
			379 => "0000000000010111110001",
			380 => "0001101101111100100000",
			381 => "0011110010001000010100",
			382 => "0001100001000100001100",
			383 => "0000010110000000001000",
			384 => "0000011110011100000100",
			385 => "0000000000011001001101",
			386 => "0000000000011001001101",
			387 => "0000000000011001001101",
			388 => "0000011100100000000100",
			389 => "0000000000011001001101",
			390 => "0000000000011001001101",
			391 => "0010111101010100001000",
			392 => "0010100011101000000100",
			393 => "0000000000011001001101",
			394 => "0000000000011001001101",
			395 => "0000000000011001001101",
			396 => "0010101000110000001100",
			397 => "0011111000001100001000",
			398 => "0001000110111100000100",
			399 => "0000000000011001001101",
			400 => "0000000000011001001101",
			401 => "0000000000011001001101",
			402 => "0000000000011001001101",
			403 => "0011000100001000011000",
			404 => "0011111110110000000100",
			405 => "0000000000011010000001",
			406 => "0010101000100100010000",
			407 => "0000110010000000001100",
			408 => "0010101001100100000100",
			409 => "0000000000011010000001",
			410 => "0011011110101100000100",
			411 => "0000000000011010000001",
			412 => "0000000000011010000001",
			413 => "0000000000011010000001",
			414 => "0000000000011010000001",
			415 => "0000000000011010000001",
			416 => "0001101110010100010100",
			417 => "0010011001111000001000",
			418 => "0000100101110100000100",
			419 => "1101010000011011100101",
			420 => "1111100000011011100101",
			421 => "0000011110100000001000",
			422 => "0011100000110000000100",
			423 => "1100100000011011100101",
			424 => "1110000000011011100101",
			425 => "1100100000011011100101",
			426 => "0001100111101000001000",
			427 => "0000101110010000000100",
			428 => "1100100000011011100101",
			429 => "1111011000011011100101",
			430 => "0011000000110000001000",
			431 => "0000101100010100000100",
			432 => "1100100000011011100101",
			433 => "1111010000011011100101",
			434 => "0001111110111100001100",
			435 => "0011011000111100000100",
			436 => "1100100000011011100101",
			437 => "0010111110111100000100",
			438 => "1101010000011011100101",
			439 => "1100100000011011100101",
			440 => "1100100000011011100101",
			441 => "0000101100010100010100",
			442 => "0001100001111000010000",
			443 => "0000100001101000000100",
			444 => "0000000000011100111001",
			445 => "0001101011111100001000",
			446 => "0000011110100000000100",
			447 => "0000000000011100111001",
			448 => "0000000000011100111001",
			449 => "0000000000011100111001",
			450 => "0000000000011100111001",
			451 => "0000011101011100010100",
			452 => "0011000100001000010000",
			453 => "0010011100100000000100",
			454 => "0000000000011100111001",
			455 => "0001001101001100001000",
			456 => "0000100011000000000100",
			457 => "0000000000011100111001",
			458 => "0000000000011100111001",
			459 => "0000000000011100111001",
			460 => "0000000000011100111001",
			461 => "0000000000011100111001",
			462 => "0000010110000000010000",
			463 => "0011111110110000001000",
			464 => "0001110000110000000100",
			465 => "0000000000011110010101",
			466 => "0000000000011110010101",
			467 => "0001111100001000000100",
			468 => "0000000000011110010101",
			469 => "0000000000011110010101",
			470 => "0001111101100000001000",
			471 => "0000011110100000000100",
			472 => "0000000000011110010101",
			473 => "1111111000011110010101",
			474 => "0001110111001000010100",
			475 => "0010000001110000010000",
			476 => "0000011001011000001100",
			477 => "0011111010010100000100",
			478 => "0000000000011110010101",
			479 => "0010000111110100000100",
			480 => "0000000000011110010101",
			481 => "0000000000011110010101",
			482 => "0000000000011110010101",
			483 => "0000000000011110010101",
			484 => "0000000000011110010101",
			485 => "0010000101000100100000",
			486 => "0000110010000000011100",
			487 => "0000101100010100010100",
			488 => "0000011110100000001100",
			489 => "0011100010111100000100",
			490 => "0000000000100000000001",
			491 => "0010001100011100000100",
			492 => "0000000000100000000001",
			493 => "0000000000100000000001",
			494 => "0010000111110100000100",
			495 => "0000000000100000000001",
			496 => "0000000000100000000001",
			497 => "0000011011111100000100",
			498 => "0000000000100000000001",
			499 => "0000000000100000000001",
			500 => "0000000000100000000001",
			501 => "0010011100110100001100",
			502 => "0011001010000000001000",
			503 => "0011010000101000000100",
			504 => "0000000000100000000001",
			505 => "0000000000100000000001",
			506 => "0000000000100000000001",
			507 => "0000101100010000001000",
			508 => "0001011000111100000100",
			509 => "0000000000100000000001",
			510 => "1111111000100000000001",
			511 => "0000000000100000000001",
			512 => "0000010000011000010100",
			513 => "0011111011000000001000",
			514 => "0011000000110000000100",
			515 => "0000000000100001101101",
			516 => "0000000000100001101101",
			517 => "0011010001111100001000",
			518 => "0010011100110100000100",
			519 => "0000001000100001101101",
			520 => "0000000000100001101101",
			521 => "0000000000100001101101",
			522 => "0000000111000000011100",
			523 => "0000011101011100011000",
			524 => "0011110011001000001100",
			525 => "0000011110100000001000",
			526 => "0011100000101000000100",
			527 => "0000000000100001101101",
			528 => "0000000000100001101101",
			529 => "0000000000100001101101",
			530 => "0010011011001100001000",
			531 => "0001010001001000000100",
			532 => "0000001000100001101101",
			533 => "0000000000100001101101",
			534 => "0000000000100001101101",
			535 => "0000000000100001101101",
			536 => "0001101011111100000100",
			537 => "0000000000100001101101",
			538 => "1111111000100001101101",
			539 => "0000010110000000011000",
			540 => "0011111110110000000100",
			541 => "0000000000100011011001",
			542 => "0011010001111100010000",
			543 => "0011010100000000000100",
			544 => "0000000000100011011001",
			545 => "0011000100010100001000",
			546 => "0011000011111100000100",
			547 => "0000000000100011011001",
			548 => "0000000000100011011001",
			549 => "0000000000100011011001",
			550 => "0000000000100011011001",
			551 => "0010011100011000001100",
			552 => "0001110111111000000100",
			553 => "0000000000100011011001",
			554 => "0001101001011000000100",
			555 => "0000000000100011011001",
			556 => "1111111000100011011001",
			557 => "0000011101011100010000",
			558 => "0001111110110000001100",
			559 => "0011001000111000000100",
			560 => "0000000000100011011001",
			561 => "0001011001010100000100",
			562 => "0000000000100011011001",
			563 => "0000000000100011011001",
			564 => "0000000000100011011001",
			565 => "0000000000100011011001",
			566 => "0000010110000000011000",
			567 => "0011111011000000001100",
			568 => "0011000000110000000100",
			569 => "0000000000100101010101",
			570 => "0011101100011100000100",
			571 => "0000000000100101010101",
			572 => "0000000000100101010101",
			573 => "0011010001111100001000",
			574 => "0000010000011000000100",
			575 => "0000001000100101010101",
			576 => "0000000000100101010101",
			577 => "0000000000100101010101",
			578 => "0000000111000000011100",
			579 => "0000011101011100011000",
			580 => "0011110011001000001100",
			581 => "0000011110100000001000",
			582 => "0000110110000100000100",
			583 => "0000000000100101010101",
			584 => "0000000000100101010101",
			585 => "0000000000100101010101",
			586 => "0010011011001100001000",
			587 => "0001010001001000000100",
			588 => "0000001000100101010101",
			589 => "0000000000100101010101",
			590 => "0000000000100101010101",
			591 => "0000000000100101010101",
			592 => "0010010010001100000100",
			593 => "0000000000100101010101",
			594 => "0010111110111100000100",
			595 => "0000000000100101010101",
			596 => "1111111000100101010101",
			597 => "0010101000100100100000",
			598 => "0010011011001100011100",
			599 => "0011111011011100001000",
			600 => "0000010110000000000100",
			601 => "0000000000100111000001",
			602 => "0000000000100111000001",
			603 => "0011000100001000010000",
			604 => "0010000011101000000100",
			605 => "0000000000100111000001",
			606 => "0001011010010100001000",
			607 => "0010000101000100000100",
			608 => "0000000000100111000001",
			609 => "0000000000100111000001",
			610 => "0000000000100111000001",
			611 => "0000000000100111000001",
			612 => "0000000000100111000001",
			613 => "0001100001111000010000",
			614 => "0001001111100000000100",
			615 => "0000000000100111000001",
			616 => "0001110100010100001000",
			617 => "0000110001110100000100",
			618 => "0000000000100111000001",
			619 => "0000000000100111000001",
			620 => "0000000000100111000001",
			621 => "0011000000111000000100",
			622 => "0000000000100111000001",
			623 => "1111111000100111000001",
			624 => "0001100001111000100100",
			625 => "0000100101001000011100",
			626 => "0010100011101000010100",
			627 => "0011111110110000000100",
			628 => "0000000000101001000101",
			629 => "0001110110000100001100",
			630 => "0000000011101000000100",
			631 => "0000000000101001000101",
			632 => "0010100010101100000100",
			633 => "0000001000101001000101",
			634 => "0000000000101001000101",
			635 => "0000000000101001000101",
			636 => "0001101011111100000100",
			637 => "0000000000101001000101",
			638 => "1111111000101001000101",
			639 => "0001110000101000000100",
			640 => "0000001000101001000101",
			641 => "0000000000101001000101",
			642 => "0000000111000000010100",
			643 => "0001010110110100001000",
			644 => "0011110011001000000100",
			645 => "0000000000101001000101",
			646 => "0000000000101001000101",
			647 => "0010000001110000000100",
			648 => "1111111000101001000101",
			649 => "0000110010010100000100",
			650 => "0000000000101001000101",
			651 => "0000000000101001000101",
			652 => "0011000000111000000100",
			653 => "0000000000101001000101",
			654 => "0001111110111100000100",
			655 => "0000000000101001000101",
			656 => "1111111000101001000101",
			657 => "0011001010000000010000",
			658 => "0000100100101000001000",
			659 => "0001101110010100000100",
			660 => "0000001000101010111001",
			661 => "0000000000101010111001",
			662 => "0000011110100000000100",
			663 => "0000001000101010111001",
			664 => "0000000000101010111001",
			665 => "0010000001110000100000",
			666 => "0011000000001100011100",
			667 => "0010101000100100010100",
			668 => "0010011001111000001000",
			669 => "0011100011111100000100",
			670 => "0000000000101010111001",
			671 => "0000000000101010111001",
			672 => "0000001001101000001000",
			673 => "0000100101110000000100",
			674 => "0000000000101010111001",
			675 => "0000000000101010111001",
			676 => "1111111000101010111001",
			677 => "0011100100101000000100",
			678 => "0000000000101010111001",
			679 => "0000001000101010111001",
			680 => "1111111000101010111001",
			681 => "0001101011111100000100",
			682 => "0000000000101010111001",
			683 => "0001111010000000000100",
			684 => "0000000000101010111001",
			685 => "1111111000101010111001",
			686 => "0001100111101000101000",
			687 => "0000010110000000010100",
			688 => "0011111010111100000100",
			689 => "1111111000101101001101",
			690 => "0001101110010100000100",
			691 => "0000001000101101001101",
			692 => "0011000000110000000100",
			693 => "0000001000101101001101",
			694 => "0001100111101000000100",
			695 => "0000000000101101001101",
			696 => "0000001000101101001101",
			697 => "0011111011011100001100",
			698 => "0001101001011000001000",
			699 => "0011111110110000000100",
			700 => "0000000000101101001101",
			701 => "0000001000101101001101",
			702 => "1111111000101101001101",
			703 => "0000011100110100000100",
			704 => "0000001000101101001101",
			705 => "1111111000101101001101",
			706 => "0011001010000000010000",
			707 => "0000100110010000001100",
			708 => "0000100011001000000100",
			709 => "1111111000101101001101",
			710 => "0011110010001000000100",
			711 => "0000001000101101001101",
			712 => "1111111000101101001101",
			713 => "0000001000101101001101",
			714 => "0000000111000000010000",
			715 => "0011000000001100001100",
			716 => "0000100010000100000100",
			717 => "1111111000101101001101",
			718 => "0010000110011100000100",
			719 => "0000000000101101001101",
			720 => "0000010000101101001101",
			721 => "1111111000101101001101",
			722 => "1111111000101101001101",
			723 => "0001101110010100010000",
			724 => "0011110111001000001000",
			725 => "0000000001110100000100",
			726 => "0000000000101111010001",
			727 => "0000000000101111010001",
			728 => "0010010110101000000100",
			729 => "0000001000101111010001",
			730 => "0000000000101111010001",
			731 => "0000000111000000011000",
			732 => "0001110111001000010100",
			733 => "0001110101101100000100",
			734 => "0000000000101111010001",
			735 => "0001111110001100000100",
			736 => "0000001000101111010001",
			737 => "0001110111001000000100",
			738 => "1111111000101111010001",
			739 => "0000011001011000000100",
			740 => "0000001000101111010001",
			741 => "0000000000101111010001",
			742 => "1111111000101111010001",
			743 => "0010111110111100001100",
			744 => "0000101110010000000100",
			745 => "1111111000101111010001",
			746 => "0001000010010000000100",
			747 => "0000000000101111010001",
			748 => "0000001000101111010001",
			749 => "0010000101000100000100",
			750 => "0000000000101111010001",
			751 => "0001010100000000000100",
			752 => "0000000000101111010001",
			753 => "0011100001010100000100",
			754 => "0000000000101111010001",
			755 => "1111111000101111010001",
			756 => "0001101110010100010100",
			757 => "0011110111001000001000",
			758 => "0011001010000000000100",
			759 => "0000000000110001011101",
			760 => "0000000000110001011101",
			761 => "0010010110101000001000",
			762 => "0000011110100000000100",
			763 => "0000001000110001011101",
			764 => "0000000000110001011101",
			765 => "0000000000110001011101",
			766 => "0000000111000000011000",
			767 => "0011000000001100010100",
			768 => "0011001000111000000100",
			769 => "1111111000110001011101",
			770 => "0001111110001100000100",
			771 => "0000001000110001011101",
			772 => "0001110111001000000100",
			773 => "1111111000110001011101",
			774 => "0000010000111100000100",
			775 => "0000001000110001011101",
			776 => "0000000000110001011101",
			777 => "1111111000110001011101",
			778 => "0001111110111100010000",
			779 => "0000100010000000001100",
			780 => "0001100111101000000100",
			781 => "0000000000110001011101",
			782 => "0010001011000100000100",
			783 => "1111111000110001011101",
			784 => "0000000000110001011101",
			785 => "0000001000110001011101",
			786 => "0010000101000100000100",
			787 => "0000000000110001011101",
			788 => "0011000000111000000100",
			789 => "0000000000110001011101",
			790 => "1111111000110001011101",
			791 => "0001100111101000011100",
			792 => "0010011001111000011000",
			793 => "0000001001101000001000",
			794 => "0011011100110000000100",
			795 => "0000010000110011011001",
			796 => "0000010000110011011001",
			797 => "0000100001001000000100",
			798 => "1111111000110011011001",
			799 => "0011000111111000001000",
			800 => "0000110001110100000100",
			801 => "0000000000110011011001",
			802 => "0000001000110011011001",
			803 => "0000000000110011011001",
			804 => "1111111000110011011001",
			805 => "0011000000110000001000",
			806 => "0000101100010100000100",
			807 => "1111111000110011011001",
			808 => "0000001000110011011001",
			809 => "0001000101110000000100",
			810 => "0000010000110011011001",
			811 => "0001110000110000001000",
			812 => "0011001010000000000100",
			813 => "1111111000110011011001",
			814 => "0000010000110011011001",
			815 => "0001001000110100001100",
			816 => "0011011101000100001000",
			817 => "0011010101100100000100",
			818 => "1111111000110011011001",
			819 => "0000000000110011011001",
			820 => "1111111000110011011001",
			821 => "1111111000110011011001",
			822 => "0000010000011000010000",
			823 => "0011111110110000000100",
			824 => "0000000000110101011101",
			825 => "0001111100001000001000",
			826 => "0011010100000000000100",
			827 => "0000000000110101011101",
			828 => "0000001000110101011101",
			829 => "0000000000110101011101",
			830 => "0000001000110000101000",
			831 => "0001000110111000011100",
			832 => "0001001010000100010000",
			833 => "0011111011000000000100",
			834 => "0000000000110101011101",
			835 => "0001110110000100001000",
			836 => "0010000000001000000100",
			837 => "0000000000110101011101",
			838 => "0000000000110101011101",
			839 => "0000000000110101011101",
			840 => "0010111001110100001000",
			841 => "0000011110100000000100",
			842 => "0000000000110101011101",
			843 => "1111111000110101011101",
			844 => "0000000000110101011101",
			845 => "0011001110001100001000",
			846 => "0000001000101100000100",
			847 => "0000000000110101011101",
			848 => "0000000000110101011101",
			849 => "0000000000110101011101",
			850 => "0010101000100100000100",
			851 => "0000000000110101011101",
			852 => "0011000000111000000100",
			853 => "0000000000110101011101",
			854 => "1111111000110101011101",
			855 => "0001100111101000101100",
			856 => "0000010110000000011100",
			857 => "0001101110010100001100",
			858 => "0001001111011000001000",
			859 => "0011111110110000000100",
			860 => "0000000000111000010001",
			861 => "0000001000111000010001",
			862 => "0000000000111000010001",
			863 => "0001111110111100001000",
			864 => "0000101110010000000100",
			865 => "0000000000111000010001",
			866 => "0000001000111000010001",
			867 => "0000110000111000000100",
			868 => "0000000000111000010001",
			869 => "1111111000111000010001",
			870 => "0011110100010000001000",
			871 => "0011111011011100000100",
			872 => "1111111000111000010001",
			873 => "0000000000111000010001",
			874 => "0000011100110100000100",
			875 => "0000001000111000010001",
			876 => "0000000000111000010001",
			877 => "0011001010000000010000",
			878 => "0010100111000100001100",
			879 => "0000100011001000000100",
			880 => "1111111000111000010001",
			881 => "0000010000011000000100",
			882 => "0000001000111000010001",
			883 => "1111111000111000010001",
			884 => "0000100000111000010001",
			885 => "0001000110101100010000",
			886 => "0010000110011000000100",
			887 => "1111111000111000010001",
			888 => "0011101110101000000100",
			889 => "0000000000111000010001",
			890 => "0000011011111100000100",
			891 => "0000001000111000010001",
			892 => "0000000000111000010001",
			893 => "0000000111000000001100",
			894 => "0010010100111100001000",
			895 => "0011111010000100000100",
			896 => "1111111000111000010001",
			897 => "0000001000111000010001",
			898 => "1111111000111000010001",
			899 => "1111111000111000010001",
			900 => "0001101110010100010000",
			901 => "0011110111001000001000",
			902 => "0010111110111100000100",
			903 => "0000000000111010011101",
			904 => "1111111000111010011101",
			905 => "0010010110101000000100",
			906 => "0000001000111010011101",
			907 => "0000000000111010011101",
			908 => "0000000111000000011000",
			909 => "0011000000001100010100",
			910 => "0011001000111000000100",
			911 => "1111111000111010011101",
			912 => "0001111110001100000100",
			913 => "0000001000111010011101",
			914 => "0001110111001000000100",
			915 => "1111111000111010011101",
			916 => "0000010000111100000100",
			917 => "0000001000111010011101",
			918 => "0000000000111010011101",
			919 => "1111111000111010011101",
			920 => "0001111110111100010000",
			921 => "0000110001110100000100",
			922 => "0000000000111010011101",
			923 => "0001000001100100001000",
			924 => "0010001011010100000100",
			925 => "0000000000111010011101",
			926 => "0000000000111010011101",
			927 => "0000001000111010011101",
			928 => "0011000000111000000100",
			929 => "0000000000111010011101",
			930 => "0010000101000100000100",
			931 => "0000000000111010011101",
			932 => "0010110000110000000100",
			933 => "0000000000111010011101",
			934 => "1111111000111010011101",
			935 => "0001100111101000100100",
			936 => "0000011110100000011000",
			937 => "0011111101010100001000",
			938 => "0000101110101100000100",
			939 => "1111111000111100111001",
			940 => "0000000000111100111001",
			941 => "0010001000010100000100",
			942 => "0000011000111100111001",
			943 => "0000100001001000000100",
			944 => "0000000000111100111001",
			945 => "0000100010110100000100",
			946 => "0000001000111100111001",
			947 => "0000010000111100111001",
			948 => "0000011110100000001000",
			949 => "0011000100010100000100",
			950 => "1111111000111100111001",
			951 => "0000011000111100111001",
			952 => "1111111000111100111001",
			953 => "0011000000110000001000",
			954 => "0000101100010100000100",
			955 => "1111111000111100111001",
			956 => "0000010000111100111001",
			957 => "0001111110111100001100",
			958 => "0000111000101100000100",
			959 => "1111111000111100111001",
			960 => "0001001101110100000100",
			961 => "1111111000111100111001",
			962 => "0000110000111100111001",
			963 => "0001000110111000010100",
			964 => "0010000110011000000100",
			965 => "1111111000111100111001",
			966 => "0001000110101100001000",
			967 => "0001000111010100000100",
			968 => "0000001000111100111001",
			969 => "0000000000111100111001",
			970 => "0001000110111000000100",
			971 => "1111111000111100111001",
			972 => "0000000000111100111001",
			973 => "1111111000111100111001",
			974 => "0000010000011000011000",
			975 => "0010011100100000001000",
			976 => "0001001111101100000100",
			977 => "0000000000111111000101",
			978 => "0000000000111111000101",
			979 => "0001111100001000001100",
			980 => "0011111010111100000100",
			981 => "0000000000111111000101",
			982 => "0011010100000000000100",
			983 => "0000000000111111000101",
			984 => "0000001000111111000101",
			985 => "0000000000111111000101",
			986 => "0010000001110000101000",
			987 => "0011000100001000100100",
			988 => "0011111010010100010100",
			989 => "0001100001000100001100",
			990 => "0011111001001000000100",
			991 => "0000000000111111000101",
			992 => "0000011001111000000100",
			993 => "0000000000111111000101",
			994 => "0000000000111111000101",
			995 => "0010101010100000000100",
			996 => "0000000000111111000101",
			997 => "0000000000111111000101",
			998 => "0000011101011100001100",
			999 => "0001011001010100001000",
			1000 => "0001111010111100000100",
			1001 => "0000000000111111000101",
			1002 => "0000001000111111000101",
			1003 => "0000000000111111000101",
			1004 => "0000000000111111000101",
			1005 => "0000000000111111000101",
			1006 => "0001101110010100000100",
			1007 => "0000000000111111000101",
			1008 => "1111111000111111000101",
			1009 => "0001100001111000101000",
			1010 => "0000101111010000100000",
			1011 => "0010100011101000011000",
			1012 => "0011111110110000000100",
			1013 => "0000000001000001010001",
			1014 => "0000010111100100010000",
			1015 => "0010101010100100001000",
			1016 => "0010000000001000000100",
			1017 => "0000000001000001010001",
			1018 => "0000001001000001010001",
			1019 => "0001110100010100000100",
			1020 => "0000000001000001010001",
			1021 => "0000000001000001010001",
			1022 => "0000000001000001010001",
			1023 => "0001101011111100000100",
			1024 => "0000000001000001010001",
			1025 => "1111111001000001010001",
			1026 => "0001110000101000000100",
			1027 => "0000001001000001010001",
			1028 => "0000000001000001010001",
			1029 => "0000101110110100000100",
			1030 => "1111111001000001010001",
			1031 => "0011000100001000011000",
			1032 => "0000000111000000010000",
			1033 => "0010111001110100001000",
			1034 => "0011110010000100000100",
			1035 => "0000000001000001010001",
			1036 => "0000000001000001010001",
			1037 => "0010110001101000000100",
			1038 => "0000001001000001010001",
			1039 => "0000000001000001010001",
			1040 => "0010111011000100000100",
			1041 => "0000000001000001010001",
			1042 => "1111111001000001010001",
			1043 => "1111111001000001010001",
			1044 => "0001100111101000011100",
			1045 => "0010010110101000011000",
			1046 => "0001101011111100001100",
			1047 => "0011110111001000000100",
			1048 => "0000000001000011101101",
			1049 => "0010000111110100000100",
			1050 => "0000001001000011101101",
			1051 => "0000001001000011101101",
			1052 => "0000101010001000000100",
			1053 => "1111111001000011101101",
			1054 => "0001011000111000000100",
			1055 => "0000001001000011101101",
			1056 => "0000000001000011101101",
			1057 => "1111111001000011101101",
			1058 => "0011001010000000010000",
			1059 => "0000100011001000000100",
			1060 => "1111111001000011101101",
			1061 => "0000010000011000001000",
			1062 => "0011000000111000000100",
			1063 => "0000001001000011101101",
			1064 => "0000001001000011101101",
			1065 => "1111111001000011101101",
			1066 => "0001001000110100100000",
			1067 => "0001001000000100010100",
			1068 => "0001011001010100010000",
			1069 => "0010111000011000001000",
			1070 => "0011110110010000000100",
			1071 => "1111111001000011101101",
			1072 => "0000000001000011101101",
			1073 => "0000101010000100000100",
			1074 => "0000000001000011101101",
			1075 => "0000010001000011101101",
			1076 => "1111111001000011101101",
			1077 => "0010101001000100000100",
			1078 => "1111111001000011101101",
			1079 => "0000010111100100000100",
			1080 => "0000000001000011101101",
			1081 => "0000010001000011101101",
			1082 => "1111111001000011101101",
			1083 => "0001100111101000100000",
			1084 => "0000011110100000011100",
			1085 => "0000100010110100001100",
			1086 => "0001101011111100001000",
			1087 => "0011010011011100000100",
			1088 => "0000000001000110001001",
			1089 => "0000001001000110001001",
			1090 => "1111111001000110001001",
			1091 => "0001101110010100001000",
			1092 => "0001000100100100000100",
			1093 => "0000001001000110001001",
			1094 => "0000000001000110001001",
			1095 => "0000010000011000000100",
			1096 => "0000001001000110001001",
			1097 => "0000000001000110001001",
			1098 => "1111111001000110001001",
			1099 => "0001000101110000000100",
			1100 => "0000010001000110001001",
			1101 => "0000000111000000010000",
			1102 => "0001111110110000001100",
			1103 => "0011110011001000000100",
			1104 => "1111111001000110001001",
			1105 => "0000011001011000000100",
			1106 => "0000001001000110001001",
			1107 => "1111111001000110001001",
			1108 => "1111111001000110001001",
			1109 => "0001111110111100001100",
			1110 => "0000100011001000000100",
			1111 => "1111111001000110001001",
			1112 => "0001100001111000000100",
			1113 => "0000001001000110001001",
			1114 => "0000000001000110001001",
			1115 => "0011000000110000001100",
			1116 => "0011100001110100001000",
			1117 => "0001010100000000000100",
			1118 => "0000000001000110001001",
			1119 => "0000000001000110001001",
			1120 => "0000000001000110001001",
			1121 => "1111111001000110001001",
			1122 => "0010011100110100010000",
			1123 => "0011111010111100000100",
			1124 => "0000000001001000001101",
			1125 => "0001011100101000001000",
			1126 => "0010011100110100000100",
			1127 => "0000001001001000001101",
			1128 => "0000000001001000001101",
			1129 => "0000000001001000001101",
			1130 => "0010000001110000101100",
			1131 => "0011000100001000101000",
			1132 => "0011111010010100010100",
			1133 => "0001100001000100001100",
			1134 => "0011111001001000000100",
			1135 => "0000000001001000001101",
			1136 => "0000100001101000000100",
			1137 => "0000000001001000001101",
			1138 => "0000000001001000001101",
			1139 => "0010101010100000000100",
			1140 => "0000000001001000001101",
			1141 => "0000000001001000001101",
			1142 => "0010010100111100010000",
			1143 => "0001110111001000001000",
			1144 => "0001110110000100000100",
			1145 => "0000000001001000001101",
			1146 => "0000000001001000001101",
			1147 => "0001010000110100000100",
			1148 => "0000001001001000001101",
			1149 => "0000000001001000001101",
			1150 => "0000000001001000001101",
			1151 => "0000000001001000001101",
			1152 => "0001101110010100000100",
			1153 => "0000000001001000001101",
			1154 => "1111111001001000001101",
			1155 => "0001101110010100010000",
			1156 => "0001011101010100001100",
			1157 => "0000101101000100001000",
			1158 => "0001100001000100000100",
			1159 => "0000001001001010100011",
			1160 => "1111111001001010100011",
			1161 => "0000001001001010100011",
			1162 => "1111111001001010100011",
			1163 => "0001000101110000000100",
			1164 => "0000001001001010100011",
			1165 => "0010011110100000011100",
			1166 => "0011110100000100010000",
			1167 => "0001100111101000001000",
			1168 => "0000101110010000000100",
			1169 => "0000000001001010100011",
			1170 => "0000000001001010100011",
			1171 => "0011111111011100000100",
			1172 => "1111111001001010100011",
			1173 => "0000000001001010100011",
			1174 => "0001101010011000001000",
			1175 => "0001011010111000000100",
			1176 => "0000001001001010100011",
			1177 => "0000000001001010100011",
			1178 => "0000010001001010100011",
			1179 => "0001000001011100010000",
			1180 => "0000001011010100000100",
			1181 => "1111111001001010100011",
			1182 => "0011101110101000000100",
			1183 => "1111111001001010100011",
			1184 => "0000110010000000000100",
			1185 => "0000001001001010100011",
			1186 => "1111111001001010100011",
			1187 => "0001100111101000001000",
			1188 => "0010000001010100000100",
			1189 => "0000000001001010100011",
			1190 => "0000000001001010100011",
			1191 => "1111111001001010100011",
			1192 => "0000000001001010100101",
			1193 => "0000000001001010101001",
			1194 => "0000000001001010101101",
			1195 => "0000000001001010110001",
			1196 => "0000000001001010110101",
			1197 => "0000000001001010111001",
			1198 => "0000000001001010111101",
			1199 => "0000000001001011000001",
			1200 => "0000000001001011000101",
			1201 => "0000000001001011001001",
			1202 => "0000000001001011001101",
			1203 => "0000000001001011010001",
			1204 => "0000000001001011010101",
			1205 => "0000000001001011011001",
			1206 => "0000000001001011011101",
			1207 => "0000000001001011100001",
			1208 => "0000000001001011100101",
			1209 => "0000000001001011101001",
			1210 => "0000000001001011101101",
			1211 => "0001111110001100000100",
			1212 => "0000000001001011111001",
			1213 => "0000000001001011111001",
			1214 => "0001110100010100000100",
			1215 => "0000000001001100000101",
			1216 => "0000000001001100000101",
			1217 => "0000010110000000001000",
			1218 => "0000011110011100000100",
			1219 => "0000000001001100011001",
			1220 => "0000000001001100011001",
			1221 => "0000000001001100011001",
			1222 => "0001100001111000001000",
			1223 => "0001101101011100000100",
			1224 => "0000000001001100101101",
			1225 => "0000000001001100101101",
			1226 => "0000000001001100101101",
			1227 => "0000010110000000001000",
			1228 => "0000011110011100000100",
			1229 => "0000000001001101000001",
			1230 => "0000000001001101000001",
			1231 => "0000000001001101000001",
			1232 => "0001110111111000000100",
			1233 => "0000000001001101010101",
			1234 => "0001110111001000000100",
			1235 => "0000000001001101010101",
			1236 => "0000000001001101010101",
			1237 => "0001111110001100001000",
			1238 => "0010011100100000000100",
			1239 => "0000000001001101101001",
			1240 => "0000000001001101101001",
			1241 => "0000000001001101101001",
			1242 => "0001101110010100000100",
			1243 => "0000000001001101111101",
			1244 => "0001101111000000000100",
			1245 => "0000000001001101111101",
			1246 => "0000000001001101111101",
			1247 => "0000011110100000001100",
			1248 => "0000011110011100000100",
			1249 => "0000000001001110011001",
			1250 => "0000010110000000000100",
			1251 => "0000000001001110011001",
			1252 => "0000000001001110011001",
			1253 => "0000000001001110011001",
			1254 => "0011111001001000000100",
			1255 => "0000000001001110110101",
			1256 => "0010111010111000001000",
			1257 => "0011001100110000000100",
			1258 => "0000000001001110110101",
			1259 => "0000000001001110110101",
			1260 => "0000000001001110110101",
			1261 => "0010111010111000001100",
			1262 => "0011111110110000000100",
			1263 => "0000000001001111010001",
			1264 => "0001111110001100000100",
			1265 => "0000000001001111010001",
			1266 => "0000000001001111010001",
			1267 => "0000000001001111010001",
			1268 => "0001100001111000001100",
			1269 => "0001101101011100000100",
			1270 => "0000000001001111101101",
			1271 => "0001101011111100000100",
			1272 => "0000000001001111101101",
			1273 => "0000000001001111101101",
			1274 => "0000000001001111101101",
			1275 => "0001101110010100000100",
			1276 => "0000000001010000001001",
			1277 => "0001101010011000001000",
			1278 => "0001101110010100000100",
			1279 => "0000000001010000001001",
			1280 => "0000000001010000001001",
			1281 => "0000000001010000001001",
			1282 => "0001101101111100001100",
			1283 => "0010101001100100000100",
			1284 => "0000000001010000101101",
			1285 => "0010101111001000000100",
			1286 => "0000000001010000101101",
			1287 => "0000000001010000101101",
			1288 => "0001101001100100000100",
			1289 => "0000000001010000101101",
			1290 => "0000000001010000101101",
			1291 => "0001101011111100001000",
			1292 => "0001101101011100000100",
			1293 => "0000000001010001010001",
			1294 => "0000000001010001010001",
			1295 => "0011000000110000000100",
			1296 => "0000000001010001010001",
			1297 => "0010110000110000000100",
			1298 => "0000000001010001010001",
			1299 => "0000000001010001010001",
			1300 => "0001101101111100001100",
			1301 => "0010000000001000000100",
			1302 => "0000000001010001111101",
			1303 => "0010100011101000000100",
			1304 => "0000000001010001111101",
			1305 => "0000000001010001111101",
			1306 => "0001101001100100001000",
			1307 => "0001000110101100000100",
			1308 => "0000000001010001111101",
			1309 => "0000000001010001111101",
			1310 => "0000000001010001111101",
			1311 => "0001110111001000010000",
			1312 => "0011110101100100000100",
			1313 => "0000000001010010100001",
			1314 => "0010000011101000000100",
			1315 => "0000000001010010100001",
			1316 => "0000011101011100000100",
			1317 => "0000000001010010100001",
			1318 => "0000000001010010100001",
			1319 => "0000000001010010100001",
			1320 => "0001110110000100010000",
			1321 => "0011010100000000000100",
			1322 => "0000000001010011000101",
			1323 => "0001101101111100001000",
			1324 => "0001101001011000000100",
			1325 => "0000000001010011000101",
			1326 => "0000000001010011000101",
			1327 => "0000000001010011000101",
			1328 => "0000000001010011000101",
			1329 => "0001111110001100010000",
			1330 => "0011110100011000000100",
			1331 => "0000000001010011101001",
			1332 => "0000011011101000001000",
			1333 => "0011001100110000000100",
			1334 => "0000000001010011101001",
			1335 => "0000000001010011101001",
			1336 => "0000000001010011101001",
			1337 => "0000000001010011101001",
			1338 => "0001111110001100010000",
			1339 => "0011111010111100000100",
			1340 => "0000000001010100001101",
			1341 => "0011001100110000001000",
			1342 => "0010110000111000000100",
			1343 => "0000000001010100001101",
			1344 => "0000000001010100001101",
			1345 => "0000000001010100001101",
			1346 => "0000000001010100001101",
			1347 => "0000010110000000010000",
			1348 => "0011111110110000000100",
			1349 => "0000000001010100111001",
			1350 => "0001011100101000001000",
			1351 => "0011000100010100000100",
			1352 => "0000000001010100111001",
			1353 => "0000000001010100111001",
			1354 => "0000000001010100111001",
			1355 => "0000001001101000000100",
			1356 => "0000000001010100111001",
			1357 => "0000000001010100111001",
			1358 => "0001111110001100010100",
			1359 => "0010110100001000001100",
			1360 => "0001101110010100001000",
			1361 => "0001101101011100000100",
			1362 => "0000000001010101100101",
			1363 => "0000000001010101100101",
			1364 => "0000000001010101100101",
			1365 => "0001100111101000000100",
			1366 => "0000000001010101100101",
			1367 => "0000000001010101100101",
			1368 => "0000000001010101100101",
			1369 => "0001101101111100010000",
			1370 => "0011111001001000000100",
			1371 => "0000000001010110011001",
			1372 => "0001110110000100001000",
			1373 => "0010100111110100000100",
			1374 => "0000000001010110011001",
			1375 => "0000000001010110011001",
			1376 => "0000000001010110011001",
			1377 => "0001000110111100000100",
			1378 => "0000000001010110011001",
			1379 => "0001101001100100000100",
			1380 => "0000000001010110011001",
			1381 => "0000000001010110011001",
			1382 => "0000011110100000010000",
			1383 => "0001011010111000001100",
			1384 => "0011010011011100000100",
			1385 => "0000000001010111010101",
			1386 => "0001011000111000000100",
			1387 => "0000000001010111010101",
			1388 => "0000000001010111010101",
			1389 => "0000000001010111010101",
			1390 => "0011010010001000001000",
			1391 => "0001101001011000000100",
			1392 => "0000000001010111010101",
			1393 => "0000000001010111010101",
			1394 => "0010011011001100000100",
			1395 => "0000000001010111010101",
			1396 => "0000000001010111010101",
			1397 => "0011001010000000010000",
			1398 => "0010111011000100001100",
			1399 => "0010011100100000000100",
			1400 => "0000000001011000010001",
			1401 => "0000011110100000000100",
			1402 => "0000000001011000010001",
			1403 => "0000000001011000010001",
			1404 => "0000000001011000010001",
			1405 => "0001101010011000001100",
			1406 => "0001101011111100000100",
			1407 => "0000000001011000010001",
			1408 => "0001111010000000000100",
			1409 => "0000000001011000010001",
			1410 => "0000000001011000010001",
			1411 => "0000000001011000010001",
			1412 => "0001111110110000010100",
			1413 => "0011111110110000000100",
			1414 => "0000000001011000111101",
			1415 => "0000011110011100000100",
			1416 => "0000000001011000111101",
			1417 => "0000011101011100001000",
			1418 => "0001011001010100000100",
			1419 => "0000000001011000111101",
			1420 => "0000000001011000111101",
			1421 => "0000000001011000111101",
			1422 => "0000000001011000111101",
			1423 => "0000101100010100011000",
			1424 => "0001101011111100001100",
			1425 => "0010010110101000001000",
			1426 => "0001101001011000000100",
			1427 => "0000000001011010000001",
			1428 => "0000000001011010000001",
			1429 => "0000000001011010000001",
			1430 => "0010100111101100000100",
			1431 => "0000000001011010000001",
			1432 => "0010010000011000000100",
			1433 => "0000000001011010000001",
			1434 => "0000000001011010000001",
			1435 => "0001111110001100001000",
			1436 => "0000011011101000000100",
			1437 => "0000000001011010000001",
			1438 => "0000000001011010000001",
			1439 => "0000000001011010000001",
			1440 => "0000101100010100001100",
			1441 => "0001100001000100000100",
			1442 => "0000000001011010111101",
			1443 => "0010100111101100000100",
			1444 => "0000000001011010111101",
			1445 => "0000000001011010111101",
			1446 => "0001111110110000010000",
			1447 => "0000011101011100001100",
			1448 => "0001001101001100001000",
			1449 => "0000100011000000000100",
			1450 => "0000000001011010111101",
			1451 => "0000000001011010111101",
			1452 => "0000000001011010111101",
			1453 => "0000000001011010111101",
			1454 => "0000000001011010111101",
			1455 => "0011001010000000010100",
			1456 => "0000101010010100000100",
			1457 => "0000000001011100000001",
			1458 => "0000011110100000001100",
			1459 => "0000011110011100000100",
			1460 => "0000000001011100000001",
			1461 => "0001110100010100000100",
			1462 => "0000000001011100000001",
			1463 => "0000000001011100000001",
			1464 => "0000000001011100000001",
			1465 => "0000100111010100001100",
			1466 => "0010111001110100001000",
			1467 => "0001111010000000000100",
			1468 => "0000000001011100000001",
			1469 => "0000000001011100000001",
			1470 => "0000000001011100000001",
			1471 => "0000000001011100000001",
			1472 => "0000011110100000010000",
			1473 => "0011111011000000000100",
			1474 => "0000000001011101001101",
			1475 => "0011000100010100001000",
			1476 => "0001101110010100000100",
			1477 => "0000000001011101001101",
			1478 => "0000000001011101001101",
			1479 => "0000000001011101001101",
			1480 => "0011111100010000001000",
			1481 => "0010100100101100000100",
			1482 => "0000000001011101001101",
			1483 => "0000000001011101001101",
			1484 => "0010011111000000001100",
			1485 => "0010110001101000001000",
			1486 => "0010011100011000000100",
			1487 => "0000000001011101001101",
			1488 => "0000000001011101001101",
			1489 => "0000000001011101001101",
			1490 => "0000000001011101001101",
			1491 => "0010010010001100001100",
			1492 => "0000111010101100000100",
			1493 => "0000000001011110011001",
			1494 => "0001111100001000000100",
			1495 => "0000000001011110011001",
			1496 => "0000000001011110011001",
			1497 => "0001101101011000010000",
			1498 => "0000001001101000000100",
			1499 => "0000000001011110011001",
			1500 => "0001101011111100000100",
			1501 => "0000000001011110011001",
			1502 => "0011000000111000000100",
			1503 => "0000000001011110011001",
			1504 => "0000000001011110011001",
			1505 => "0000011101011100001000",
			1506 => "0000011101011100000100",
			1507 => "0000000001011110011001",
			1508 => "0000000001011110011001",
			1509 => "0000000001011110011001",
			1510 => "0001101101111100011100",
			1511 => "0011110010001000010100",
			1512 => "0001100001000100001100",
			1513 => "0000010110000000001000",
			1514 => "0000011110011100000100",
			1515 => "0000000001011111101101",
			1516 => "0000000001011111101101",
			1517 => "0000000001011111101101",
			1518 => "0000011100100000000100",
			1519 => "0000000001011111101101",
			1520 => "0000000001011111101101",
			1521 => "0010111101010100000100",
			1522 => "0000000001011111101101",
			1523 => "0000000001011111101101",
			1524 => "0000101011111000001000",
			1525 => "0010111001110100000100",
			1526 => "0000000001011111101101",
			1527 => "0000000001011111101101",
			1528 => "0011000011011100000100",
			1529 => "0000000001011111101101",
			1530 => "0000000001011111101101",
			1531 => "0001111110001100100000",
			1532 => "0000101110010000010100",
			1533 => "0010101010100000001100",
			1534 => "0011100100000000000100",
			1535 => "0000000001100000111001",
			1536 => "0001101001011000000100",
			1537 => "0000000001100000111001",
			1538 => "0000000001100000111001",
			1539 => "0001100001000100000100",
			1540 => "0000000001100000111001",
			1541 => "0000000001100000111001",
			1542 => "0000011011101000001000",
			1543 => "0011000011011100000100",
			1544 => "0000000001100000111001",
			1545 => "0000000001100000111001",
			1546 => "0000000001100000111001",
			1547 => "0001101001100100000100",
			1548 => "0000000001100000111001",
			1549 => "0000000001100000111001",
			1550 => "0010000001110000011000",
			1551 => "0001111110110000010100",
			1552 => "0011111110110000000100",
			1553 => "0000000001100001111101",
			1554 => "0000011001011000001100",
			1555 => "0010000000001000000100",
			1556 => "0000000001100001111101",
			1557 => "0001011001010100000100",
			1558 => "0000000001100001111101",
			1559 => "0000000001100001111101",
			1560 => "0000000001100001111101",
			1561 => "0000000001100001111101",
			1562 => "0001101110010100000100",
			1563 => "0000000001100001111101",
			1564 => "0010010110000000000100",
			1565 => "0000000001100001111101",
			1566 => "0000000001100001111101",
			1567 => "0010111011000100011000",
			1568 => "0011010000101000000100",
			1569 => "0000000001100011001001",
			1570 => "0011001010000000010000",
			1571 => "0010011001111000001100",
			1572 => "0001110100010100001000",
			1573 => "0010011100100000000100",
			1574 => "0000000001100011001001",
			1575 => "0000000001100011001001",
			1576 => "0000000001100011001001",
			1577 => "0000000001100011001001",
			1578 => "0000000001100011001001",
			1579 => "0011010010001000001000",
			1580 => "0010010010001100000100",
			1581 => "0000000001100011001001",
			1582 => "0000000001100011001001",
			1583 => "0010011011001100000100",
			1584 => "0000000001100011001001",
			1585 => "0000000001100011001001",
			1586 => "0001101101111100100000",
			1587 => "0011111010010100010100",
			1588 => "0001101011111100001100",
			1589 => "0011110111001000000100",
			1590 => "0000000001100100101101",
			1591 => "0001010100011000000100",
			1592 => "0000000001100100101101",
			1593 => "0000000001100100101101",
			1594 => "0010010110000000000100",
			1595 => "0000000001100100101101",
			1596 => "0000000001100100101101",
			1597 => "0001110110000100001000",
			1598 => "0010100001010000000100",
			1599 => "0000000001100100101101",
			1600 => "0000000001100100101101",
			1601 => "0000000001100100101101",
			1602 => "0000101100111000001000",
			1603 => "0001110111001000000100",
			1604 => "1111111001100100101101",
			1605 => "0000000001100100101101",
			1606 => "0001110111001000001000",
			1607 => "0000100011000000000100",
			1608 => "0000000001100100101101",
			1609 => "0000000001100100101101",
			1610 => "0000000001100100101101",
			1611 => "0010000101000100011000",
			1612 => "0011000100001000010100",
			1613 => "0011100010111100000100",
			1614 => "0000000001100101111001",
			1615 => "0011100011001000001100",
			1616 => "0010100011101000001000",
			1617 => "0010000000001000000100",
			1618 => "0000000001100101111001",
			1619 => "0000000001100101111001",
			1620 => "0000000001100101111001",
			1621 => "0000000001100101111001",
			1622 => "0000000001100101111001",
			1623 => "0011000000110000000100",
			1624 => "0000000001100101111001",
			1625 => "0011100111010100001000",
			1626 => "0011100001010100000100",
			1627 => "0000000001100101111001",
			1628 => "0000000001100101111001",
			1629 => "0000000001100101111001",
			1630 => "0001101101111100100100",
			1631 => "0011111010010100011000",
			1632 => "0001100001000100001100",
			1633 => "0011111010111100000100",
			1634 => "0000000001100111101101",
			1635 => "0001010100011000000100",
			1636 => "0000000001100111101101",
			1637 => "0000000001100111101101",
			1638 => "0000010000011000000100",
			1639 => "0000000001100111101101",
			1640 => "0010101010100000000100",
			1641 => "0000000001100111101101",
			1642 => "0000000001100111101101",
			1643 => "0001110110000100001000",
			1644 => "0010100001010000000100",
			1645 => "0000000001100111101101",
			1646 => "0000000001100111101101",
			1647 => "0000000001100111101101",
			1648 => "0000101100111000001100",
			1649 => "0001110111001000001000",
			1650 => "0000011100100000000100",
			1651 => "0000000001100111101101",
			1652 => "1111111001100111101101",
			1653 => "0000000001100111101101",
			1654 => "0001110111001000001000",
			1655 => "0000100011000000000100",
			1656 => "0000000001100111101101",
			1657 => "0000000001100111101101",
			1658 => "0000000001100111101101",
			1659 => "0000101100010100010100",
			1660 => "0001100001111000010000",
			1661 => "0000100001101000000100",
			1662 => "0000000001101001000001",
			1663 => "0001101011111100001000",
			1664 => "0000011110100000000100",
			1665 => "0000000001101001000001",
			1666 => "0000000001101001000001",
			1667 => "0000000001101001000001",
			1668 => "0000000001101001000001",
			1669 => "0000011101011100010100",
			1670 => "0011000100001000010000",
			1671 => "0010011100100000000100",
			1672 => "0000000001101001000001",
			1673 => "0000000110110100001000",
			1674 => "0000100011000000000100",
			1675 => "0000000001101001000001",
			1676 => "0000000001101001000001",
			1677 => "0000000001101001000001",
			1678 => "0000000001101001000001",
			1679 => "0000000001101001000001",
			1680 => "0000010110000000011000",
			1681 => "0000100100101000010000",
			1682 => "0001101011111100001000",
			1683 => "0000110000111000000100",
			1684 => "0000000001101010111101",
			1685 => "0000000001101010111101",
			1686 => "0011100000110000000100",
			1687 => "0000000001101010111101",
			1688 => "0000000001101010111101",
			1689 => "0001110000101000000100",
			1690 => "0000000001101010111101",
			1691 => "0000000001101010111101",
			1692 => "0001110101101100010000",
			1693 => "0000000101000100000100",
			1694 => "0000000001101010111101",
			1695 => "0000101100010000001000",
			1696 => "0011000000111000000100",
			1697 => "0000000001101010111101",
			1698 => "1111111001101010111101",
			1699 => "0000000001101010111101",
			1700 => "0001111110001100001100",
			1701 => "0001101010011000001000",
			1702 => "0000100000110100000100",
			1703 => "0000000001101010111101",
			1704 => "0000000001101010111101",
			1705 => "0000000001101010111101",
			1706 => "0001101001100100001000",
			1707 => "0001000110111100000100",
			1708 => "0000000001101010111101",
			1709 => "0000000001101010111101",
			1710 => "0000000001101010111101",
			1711 => "0010101001000100100100",
			1712 => "0001111110110000100000",
			1713 => "0011101110101000010100",
			1714 => "0000011110100000001100",
			1715 => "0011010100000000000100",
			1716 => "0000000001101100011001",
			1717 => "0001101110010100000100",
			1718 => "0000000001101100011001",
			1719 => "0000000001101100011001",
			1720 => "0001001110010000000100",
			1721 => "0000000001101100011001",
			1722 => "0000000001101100011001",
			1723 => "0010011011001100001000",
			1724 => "0000001001101000000100",
			1725 => "0000000001101100011001",
			1726 => "0000000001101100011001",
			1727 => "0000000001101100011001",
			1728 => "0000000001101100011001",
			1729 => "0001100001111000000100",
			1730 => "0000000001101100011001",
			1731 => "0000011100100000000100",
			1732 => "0000000001101100011001",
			1733 => "0000000001101100011001",
			1734 => "0000010110000000011000",
			1735 => "0000100100101000010000",
			1736 => "0001101011111100001000",
			1737 => "0000111000101100000100",
			1738 => "0000000001101110000101",
			1739 => "0000000001101110000101",
			1740 => "0011100000110000000100",
			1741 => "0000000001101110000101",
			1742 => "0000000001101110000101",
			1743 => "0001110000101000000100",
			1744 => "0000001001101110000101",
			1745 => "0000000001101110000101",
			1746 => "0011000011011100001000",
			1747 => "0001101110010100000100",
			1748 => "0000000001101110000101",
			1749 => "1111111001101110000101",
			1750 => "0011000000001100010100",
			1751 => "0011101011011100000100",
			1752 => "0000000001101110000101",
			1753 => "0000000111000000001100",
			1754 => "0000000110011100000100",
			1755 => "0000000001101110000101",
			1756 => "0001110111001000000100",
			1757 => "0000001001101110000101",
			1758 => "0000000001101110000101",
			1759 => "0000000001101110000101",
			1760 => "0000000001101110000101",
			1761 => "0000010110000000011000",
			1762 => "0011111110110000000100",
			1763 => "0000000001101111110001",
			1764 => "0011010001111100010000",
			1765 => "0011010100000000000100",
			1766 => "0000000001101111110001",
			1767 => "0011000100010100001000",
			1768 => "0011000011111100000100",
			1769 => "0000000001101111110001",
			1770 => "0000000001101111110001",
			1771 => "0000000001101111110001",
			1772 => "0000000001101111110001",
			1773 => "0000011101101000001100",
			1774 => "0001111110111100000100",
			1775 => "0000000001101111110001",
			1776 => "0001101001011000000100",
			1777 => "0000000001101111110001",
			1778 => "0000000001101111110001",
			1779 => "0000011101011100010000",
			1780 => "0011000100001000001100",
			1781 => "0011001000111000000100",
			1782 => "0000000001101111110001",
			1783 => "0001111110110000000100",
			1784 => "0000000001101111110001",
			1785 => "0000000001101111110001",
			1786 => "0000000001101111110001",
			1787 => "0000000001101111110001",
			1788 => "0000010110000000011000",
			1789 => "0011111011000000001100",
			1790 => "0011000000110000000100",
			1791 => "0000000001110001101101",
			1792 => "0001110000110000000100",
			1793 => "0000000001110001101101",
			1794 => "0000000001110001101101",
			1795 => "0011010001111100001000",
			1796 => "0000010000011000000100",
			1797 => "0000001001110001101101",
			1798 => "0000000001110001101101",
			1799 => "0000000001110001101101",
			1800 => "0000000111000000011100",
			1801 => "0000011101011100011000",
			1802 => "0011110011001000001100",
			1803 => "0000011110100000001000",
			1804 => "0000110110000100000100",
			1805 => "0000000001110001101101",
			1806 => "0000000001110001101101",
			1807 => "0000000001110001101101",
			1808 => "0010011011001100001000",
			1809 => "0011010010110100000100",
			1810 => "0000001001110001101101",
			1811 => "0000000001110001101101",
			1812 => "0000000001110001101101",
			1813 => "0000000001110001101101",
			1814 => "0010010010001100000100",
			1815 => "0000000001110001101101",
			1816 => "0010000101000100000100",
			1817 => "0000000001110001101101",
			1818 => "1111111001110001101101",
			1819 => "0010000101000100100100",
			1820 => "0000110010000000100000",
			1821 => "0000101100010100011000",
			1822 => "0010101010100000001100",
			1823 => "0011011010011100001000",
			1824 => "0000100001101000000100",
			1825 => "0000000001110011100001",
			1826 => "0000000001110011100001",
			1827 => "0000000001110011100001",
			1828 => "0000010110000000000100",
			1829 => "0000000001110011100001",
			1830 => "0010111011000100000100",
			1831 => "0000000001110011100001",
			1832 => "0000000001110011100001",
			1833 => "0000011011111100000100",
			1834 => "0000001001110011100001",
			1835 => "0000000001110011100001",
			1836 => "0000000001110011100001",
			1837 => "0001101110010100001000",
			1838 => "0011011100110000000100",
			1839 => "0000000001110011100001",
			1840 => "0000000001110011100001",
			1841 => "0010010110000000000100",
			1842 => "0000000001110011100001",
			1843 => "0000000111000000000100",
			1844 => "0000000001110011100001",
			1845 => "0011000000111000000100",
			1846 => "0000000001110011100001",
			1847 => "1111111001110011100001",
			1848 => "0011001010000000011000",
			1849 => "0000010000011000001000",
			1850 => "0011111010111100000100",
			1851 => "0000000001110101100101",
			1852 => "0000001001110101100101",
			1853 => "0011101011000100001000",
			1854 => "0011110111110000000100",
			1855 => "0000000001110101100101",
			1856 => "0000000001110101100101",
			1857 => "0010101001000100000100",
			1858 => "0000000001110101100101",
			1859 => "0000000001110101100101",
			1860 => "0000000111000000011100",
			1861 => "0011000000001100011000",
			1862 => "0011000011011100001100",
			1863 => "0000011110100000001000",
			1864 => "0011101110111100000100",
			1865 => "0000000001110101100101",
			1866 => "0000000001110101100101",
			1867 => "0000000001110101100101",
			1868 => "0010000111110100000100",
			1869 => "0000000001110101100101",
			1870 => "0000010101011100000100",
			1871 => "0000001001110101100101",
			1872 => "0000000001110101100101",
			1873 => "0000000001110101100101",
			1874 => "0010000101000100000100",
			1875 => "0000000001110101100101",
			1876 => "0001111010000000000100",
			1877 => "0000000001110101100101",
			1878 => "0010110000110000000100",
			1879 => "0000000001110101100101",
			1880 => "1111111001110101100101",
			1881 => "0001100001111000100100",
			1882 => "0000100101001000011100",
			1883 => "0010100011101000010100",
			1884 => "0011111110110000000100",
			1885 => "0000000001110111110001",
			1886 => "0001110110000100001100",
			1887 => "0000000011101000000100",
			1888 => "0000000001110111110001",
			1889 => "0010100010101100000100",
			1890 => "0000001001110111110001",
			1891 => "0000000001110111110001",
			1892 => "0000000001110111110001",
			1893 => "0001101011111100000100",
			1894 => "0000000001110111110001",
			1895 => "1111111001110111110001",
			1896 => "0001110000101000000100",
			1897 => "0000001001110111110001",
			1898 => "0000000001110111110001",
			1899 => "0000000111000000011000",
			1900 => "0000000010101000001100",
			1901 => "0011101001010000001000",
			1902 => "0011111100010100000100",
			1903 => "0000000001110111110001",
			1904 => "0000000001110111110001",
			1905 => "1111111001110111110001",
			1906 => "0011001110001100001000",
			1907 => "0010100111110100000100",
			1908 => "0000000001110111110001",
			1909 => "0000001001110111110001",
			1910 => "0000000001110111110001",
			1911 => "0011000000111000000100",
			1912 => "0000000001110111110001",
			1913 => "0001111110111100000100",
			1914 => "0000000001110111110001",
			1915 => "1111111001110111110001",
			1916 => "0011001010000000011100",
			1917 => "0010011100110100001100",
			1918 => "0011111010111100000100",
			1919 => "0000000001111001110101",
			1920 => "0011010100000000000100",
			1921 => "0000000001111001110101",
			1922 => "0000001001111001110101",
			1923 => "0011101000111100001000",
			1924 => "0011101011000100000100",
			1925 => "0000000001111001110101",
			1926 => "0000000001111001110101",
			1927 => "0010101001000100000100",
			1928 => "0000000001111001110101",
			1929 => "0000000001111001110101",
			1930 => "0010000001110000100000",
			1931 => "0011000000001100011100",
			1932 => "0010101000100100010100",
			1933 => "0010011001111000001000",
			1934 => "0011100011111100000100",
			1935 => "0000000001111001110101",
			1936 => "0000000001111001110101",
			1937 => "0000001001101000001000",
			1938 => "0011111001011100000100",
			1939 => "0000000001111001110101",
			1940 => "0000000001111001110101",
			1941 => "1111111001111001110101",
			1942 => "0011100100101000000100",
			1943 => "0000000001111001110101",
			1944 => "0000001001111001110101",
			1945 => "1111111001111001110101",
			1946 => "0001111010000000000100",
			1947 => "0000000001111001110101",
			1948 => "1111111001111001110101",
			1949 => "0001100111101000100000",
			1950 => "0000011110100000010100",
			1951 => "0011111010111100000100",
			1952 => "1111111001111100000001",
			1953 => "0010001000010100000100",
			1954 => "0000010001111100000001",
			1955 => "0011000100010100001000",
			1956 => "0000110000001100000100",
			1957 => "0000001001111100000001",
			1958 => "0000001001111100000001",
			1959 => "0000000001111100000001",
			1960 => "0000011110100000001000",
			1961 => "0011010110000100000100",
			1962 => "1111111001111100000001",
			1963 => "0000001001111100000001",
			1964 => "1111111001111100000001",
			1965 => "0011000000110000001100",
			1966 => "0011111110110000000100",
			1967 => "1111111001111100000001",
			1968 => "0000010000011000000100",
			1969 => "0000001001111100000001",
			1970 => "1111111001111100000001",
			1971 => "0001000101110000000100",
			1972 => "0000001001111100000001",
			1973 => "0001110000110000001000",
			1974 => "0011001010000000000100",
			1975 => "1111111001111100000001",
			1976 => "0000001001111100000001",
			1977 => "0001001000110100001100",
			1978 => "0001011001010100001000",
			1979 => "0011100011001000000100",
			1980 => "1111111001111100000001",
			1981 => "0000011001111100000001",
			1982 => "1111111001111100000001",
			1983 => "1111111001111100000001",
			1984 => "0001101110010100010000",
			1985 => "0010010110101000001100",
			1986 => "0011110111001000000100",
			1987 => "0000000001111110010101",
			1988 => "0001001111011000000100",
			1989 => "0000001001111110010101",
			1990 => "0000000001111110010101",
			1991 => "1111111001111110010101",
			1992 => "0011001010000000011000",
			1993 => "0000101110010000001000",
			1994 => "0000101010001000000100",
			1995 => "1111111001111110010101",
			1996 => "0000000001111110010101",
			1997 => "0000010110000000001000",
			1998 => "0001101101111100000100",
			1999 => "0000001001111110010101",
			2000 => "0000010001111110010101",
			2001 => "0001000000010100000100",
			2002 => "0000000001111110010101",
			2003 => "1111111001111110010101",
			2004 => "0001000110101100010000",
			2005 => "0010000110011000000100",
			2006 => "1111111001111110010101",
			2007 => "0011110011001000000100",
			2008 => "0000000001111110010101",
			2009 => "0011000100001000000100",
			2010 => "0000001001111110010101",
			2011 => "0000000001111110010101",
			2012 => "0000000111000000001100",
			2013 => "0001110111001000001000",
			2014 => "0000101000001100000100",
			2015 => "1111111001111110010101",
			2016 => "0000001001111110010101",
			2017 => "1111111001111110010101",
			2018 => "0001111010000000000100",
			2019 => "0000000001111110010101",
			2020 => "1111111001111110010101",
			2021 => "0001101110010100010100",
			2022 => "0000010110000000001000",
			2023 => "0000100001001000000100",
			2024 => "0000000010000000010001",
			2025 => "0000001010000000010001",
			2026 => "0011111010011100000100",
			2027 => "1111111010000000010001",
			2028 => "0010010110101000000100",
			2029 => "0000000010000000010001",
			2030 => "0000000010000000010001",
			2031 => "0001000101110000000100",
			2032 => "0000001010000000010001",
			2033 => "0011001010000000010100",
			2034 => "0000101100010100001000",
			2035 => "0010000100010100000100",
			2036 => "1111111010000000010001",
			2037 => "0000000010000000010001",
			2038 => "0010111011000100001000",
			2039 => "0000001010011100000100",
			2040 => "0000001010000000010001",
			2041 => "0000010010000000010001",
			2042 => "0000000010000000010001",
			2043 => "0001000001011100010000",
			2044 => "0000001011010100000100",
			2045 => "1111111010000000010001",
			2046 => "0011000011011100000100",
			2047 => "1111111010000000010001",
			2048 => "0001111110110000000100",
			2049 => "0000001010000000010001",
			2050 => "0000000010000000010001",
			2051 => "1111111010000000010001",
			2052 => "0001101110010100011100",
			2053 => "0000100010110100010100",
			2054 => "0000010110000000001000",
			2055 => "0001010011011100000100",
			2056 => "0000000010000010110101",
			2057 => "0000001010000010110101",
			2058 => "0011101000111000000100",
			2059 => "1111111010000010110101",
			2060 => "0010110101101100000100",
			2061 => "0000000010000010110101",
			2062 => "0000000010000010110101",
			2063 => "0000011110100000000100",
			2064 => "0000001010000010110101",
			2065 => "0000000010000010110101",
			2066 => "0000100111010100100100",
			2067 => "0011110011001000010100",
			2068 => "0000010000011000001100",
			2069 => "0000101010001000000100",
			2070 => "0000000010000010110101",
			2071 => "0001010100011000000100",
			2072 => "0000000010000010110101",
			2073 => "0000000010000010110101",
			2074 => "0001010100000000000100",
			2075 => "0000000010000010110101",
			2076 => "1111111010000010110101",
			2077 => "0001110110000100001000",
			2078 => "0000001000110000000100",
			2079 => "0000001010000010110101",
			2080 => "0000000010000010110101",
			2081 => "0010001010110000000100",
			2082 => "1111111010000010110101",
			2083 => "0000000010000010110101",
			2084 => "0011000000001100010000",
			2085 => "0001101000010000001100",
			2086 => "0000011101011100001000",
			2087 => "0000100011000000000100",
			2088 => "0000001010000010110101",
			2089 => "0000000010000010110101",
			2090 => "0000000010000010110101",
			2091 => "0000000010000010110101",
			2092 => "1111111010000010110101",
			2093 => "0001100001111000110100",
			2094 => "0000010110000000011000",
			2095 => "0001101110010100001100",
			2096 => "0000011110011100000100",
			2097 => "0000000010000101101001",
			2098 => "0011011100001000000100",
			2099 => "0000000010000101101001",
			2100 => "0000001010000101101001",
			2101 => "0000101010001000000100",
			2102 => "1111111010000101101001",
			2103 => "0001111110111100000100",
			2104 => "0000001010000101101001",
			2105 => "0000000010000101101001",
			2106 => "0001100111101000010100",
			2107 => "0001110111111000001000",
			2108 => "0000101110101000000100",
			2109 => "0000000010000101101001",
			2110 => "0000000010000101101001",
			2111 => "0001100101011100001000",
			2112 => "0011011110110000000100",
			2113 => "0000000010000101101001",
			2114 => "0000000010000101101001",
			2115 => "1111111010000101101001",
			2116 => "0001001110010000000100",
			2117 => "0000010010000101101001",
			2118 => "0000000010000101101001",
			2119 => "0001000001011100010000",
			2120 => "0000001011010100000100",
			2121 => "1111111010000101101001",
			2122 => "0010011011001100001000",
			2123 => "0000110111100000000100",
			2124 => "0000000010000101101001",
			2125 => "0000001010000101101001",
			2126 => "1111111010000101101001",
			2127 => "0011101001101000001000",
			2128 => "0000101111010100000100",
			2129 => "1111111010000101101001",
			2130 => "0000010010000101101001",
			2131 => "0001111110111100001100",
			2132 => "0001111110111100001000",
			2133 => "0001011000111100000100",
			2134 => "0000000010000101101001",
			2135 => "0000000010000101101001",
			2136 => "0000000010000101101001",
			2137 => "1111111010000101101001",
			2138 => "0001100111101000011100",
			2139 => "0000011110100000011000",
			2140 => "0010100100101100000100",
			2141 => "0000010010000111101101",
			2142 => "0011000100010100010000",
			2143 => "0000110001110100000100",
			2144 => "0000000010000111101101",
			2145 => "0000100001001000000100",
			2146 => "0000000010000111101101",
			2147 => "0000110000001100000100",
			2148 => "0000001010000111101101",
			2149 => "0000001010000111101101",
			2150 => "1111111010000111101101",
			2151 => "1111111010000111101101",
			2152 => "0001111110111100001100",
			2153 => "0000100011001000000100",
			2154 => "1111111010000111101101",
			2155 => "0000101001100000000100",
			2156 => "0000001010000111101101",
			2157 => "0000010010000111101101",
			2158 => "0011000000111000001000",
			2159 => "0010001110111100000100",
			2160 => "0000000010000111101101",
			2161 => "0000000010000111101101",
			2162 => "0001001000110100010000",
			2163 => "0001001000000100000100",
			2164 => "1111111010000111101101",
			2165 => "0010000001110000000100",
			2166 => "1111111010000111101101",
			2167 => "0000001000110000000100",
			2168 => "0000100010000111101101",
			2169 => "1111111010000111101101",
			2170 => "1111111010000111101101",
			2171 => "0000010000011000010100",
			2172 => "0011000100010100010000",
			2173 => "0011111010111100000100",
			2174 => "0000000010001001100001",
			2175 => "0000010000011000000100",
			2176 => "0000001010001001100001",
			2177 => "0010101001000100000100",
			2178 => "0000000010001001100001",
			2179 => "0000000010001001100001",
			2180 => "0000000010001001100001",
			2181 => "0010000001110000100100",
			2182 => "0011000100001000100000",
			2183 => "0011111010010100010000",
			2184 => "0010010010001100001000",
			2185 => "0011010011011100000100",
			2186 => "0000000010001001100001",
			2187 => "0000000010001001100001",
			2188 => "0010100100111100000100",
			2189 => "0000000010001001100001",
			2190 => "1111111010001001100001",
			2191 => "0000011101011100001100",
			2192 => "0000101100010000001000",
			2193 => "0001001010000100000100",
			2194 => "0000001010001001100001",
			2195 => "0000000010001001100001",
			2196 => "0000001010001001100001",
			2197 => "0000000010001001100001",
			2198 => "1111111010001001100001",
			2199 => "1111111010001001100001",
			2200 => "0001100111101000011100",
			2201 => "0000011110100000011000",
			2202 => "0001101110010100010000",
			2203 => "0010000111110100000100",
			2204 => "0000010010001011111101",
			2205 => "0010010010001100000100",
			2206 => "0000001010001011111101",
			2207 => "0010110100010100000100",
			2208 => "0000001010001011111101",
			2209 => "0000000010001011111101",
			2210 => "0000101110010000000100",
			2211 => "1111111010001011111101",
			2212 => "0000001010001011111101",
			2213 => "1111111010001011111101",
			2214 => "0001111110111100001100",
			2215 => "0000100011001000000100",
			2216 => "1111111010001011111101",
			2217 => "0011011000111000000100",
			2218 => "0000001010001011111101",
			2219 => "0000001010001011111101",
			2220 => "0010100011101000010000",
			2221 => "0001010111110000001100",
			2222 => "0011001000111000000100",
			2223 => "1111111010001011111101",
			2224 => "0010011011001100000100",
			2225 => "0000011010001011111101",
			2226 => "0000000010001011111101",
			2227 => "1111111010001011111101",
			2228 => "0011001010000000010100",
			2229 => "0011001010000000001100",
			2230 => "0011000000110000001000",
			2231 => "0010010110000000000100",
			2232 => "0000000010001011111101",
			2233 => "1111111010001011111101",
			2234 => "1111111010001011111101",
			2235 => "0000111010000000000100",
			2236 => "0000100010001011111101",
			2237 => "0000000010001011111101",
			2238 => "1111111010001011111101",
			2239 => "0001100111101000011100",
			2240 => "0010010110101000011000",
			2241 => "0001101110010100010000",
			2242 => "0011111101010100000100",
			2243 => "0000000010001110010001",
			2244 => "0010000111110100000100",
			2245 => "0000010010001110010001",
			2246 => "0010010010001100000100",
			2247 => "0000001010001110010001",
			2248 => "0000000010001110010001",
			2249 => "0000101110010000000100",
			2250 => "1111111010001110010001",
			2251 => "0000001010001110010001",
			2252 => "1111111010001110010001",
			2253 => "0001111110111100001100",
			2254 => "0000100011001000000100",
			2255 => "1111111010001110010001",
			2256 => "0011110110110100000100",
			2257 => "0000001010001110010001",
			2258 => "0000000010001110010001",
			2259 => "0001000101110000000100",
			2260 => "0000001010001110010001",
			2261 => "0001000110101100001100",
			2262 => "0011000100001000001000",
			2263 => "0000101100010100000100",
			2264 => "1111111010001110010001",
			2265 => "0000011010001110010001",
			2266 => "1111111010001110010001",
			2267 => "0011001010000000010000",
			2268 => "0011001010000000001000",
			2269 => "0011000000110000000100",
			2270 => "0000000010001110010001",
			2271 => "1111111010001110010001",
			2272 => "0000111010000000000100",
			2273 => "0000011010001110010001",
			2274 => "0000000010001110010001",
			2275 => "1111111010001110010001",
			2276 => "0001101110010100011100",
			2277 => "0000100010110100010100",
			2278 => "0000010110000000001000",
			2279 => "0001010011011100000100",
			2280 => "0000000010010001001101",
			2281 => "0000000010010001001101",
			2282 => "0011101000111000000100",
			2283 => "0000000010010001001101",
			2284 => "0011011110110000000100",
			2285 => "0000000010010001001101",
			2286 => "0000000010010001001101",
			2287 => "0000011110100000000100",
			2288 => "0000001010010001001101",
			2289 => "0000000010010001001101",
			2290 => "0000100111010100110000",
			2291 => "0011110011001000011100",
			2292 => "0000010000011000001100",
			2293 => "0000101010001000000100",
			2294 => "0000000010010001001101",
			2295 => "0001010100011000000100",
			2296 => "0000000010010001001101",
			2297 => "0000000010010001001101",
			2298 => "0001010100000000000100",
			2299 => "0000000010010001001101",
			2300 => "0000101100010000000100",
			2301 => "1111111010010001001101",
			2302 => "0000101100010000000100",
			2303 => "0000000010010001001101",
			2304 => "0000000010010001001101",
			2305 => "0001101101111100001000",
			2306 => "0011100111111100000100",
			2307 => "0000001010010001001101",
			2308 => "0000000010010001001101",
			2309 => "0011111100010000000100",
			2310 => "1111111010010001001101",
			2311 => "0011111100000000000100",
			2312 => "0000000010010001001101",
			2313 => "0000000010010001001101",
			2314 => "0011000000001100010000",
			2315 => "0001101000010000001100",
			2316 => "0000011101011100001000",
			2317 => "0000100011000000000100",
			2318 => "0000001010010001001101",
			2319 => "0000000010010001001101",
			2320 => "0000000010010001001101",
			2321 => "0000000010010001001101",
			2322 => "1111111010010001001101",
			2323 => "0001100111101000100000",
			2324 => "0010010110101000011100",
			2325 => "0000100010110100001100",
			2326 => "0001101011111100001000",
			2327 => "0000110100000000000100",
			2328 => "0000000010010011100001",
			2329 => "0000001010010011100001",
			2330 => "1111111010010011100001",
			2331 => "0001101110010100001000",
			2332 => "0000110000001100000100",
			2333 => "0000001010010011100001",
			2334 => "0000001010010011100001",
			2335 => "0000010000011000000100",
			2336 => "0000001010010011100001",
			2337 => "0000000010010011100001",
			2338 => "1111111010010011100001",
			2339 => "0001000101110000000100",
			2340 => "0000011010010011100001",
			2341 => "0001111110111100001000",
			2342 => "0000100011001000000100",
			2343 => "1111111010010011100001",
			2344 => "0000001010010011100001",
			2345 => "0000000111000000010000",
			2346 => "0011000100001000001100",
			2347 => "0011110011001000000100",
			2348 => "1111111010010011100001",
			2349 => "0000011001011000000100",
			2350 => "0000010010010011100001",
			2351 => "1111111010010011100001",
			2352 => "1111111010010011100001",
			2353 => "0011000000110000001100",
			2354 => "0010110111111000001000",
			2355 => "0010111110111100000100",
			2356 => "0000000010010011100001",
			2357 => "1111111010010011100001",
			2358 => "0000000010010011100001",
			2359 => "1111111010010011100001",
			2360 => "0001101110010100011100",
			2361 => "0000100010110100010100",
			2362 => "0000010110000000001000",
			2363 => "0001010011011100000100",
			2364 => "0000000010010110100101",
			2365 => "0000000010010110100101",
			2366 => "0000110101101100000100",
			2367 => "0000000010010110100101",
			2368 => "0010110101101100000100",
			2369 => "0000000010010110100101",
			2370 => "0000000010010110100101",
			2371 => "0000011110100000000100",
			2372 => "0000001010010110100101",
			2373 => "0000000010010110100101",
			2374 => "0000100111010100110000",
			2375 => "0011110011001000011100",
			2376 => "0000010000011000001100",
			2377 => "0000101010001000000100",
			2378 => "0000000010010110100101",
			2379 => "0001010100011000000100",
			2380 => "0000000010010110100101",
			2381 => "0000000010010110100101",
			2382 => "0000101100010000001000",
			2383 => "0001010100000000000100",
			2384 => "0000000010010110100101",
			2385 => "1111111010010110100101",
			2386 => "0001010101101100000100",
			2387 => "0000000010010110100101",
			2388 => "0000000010010110100101",
			2389 => "0001101101111100001000",
			2390 => "0010011010011000000100",
			2391 => "0000001010010110100101",
			2392 => "0000000010010110100101",
			2393 => "0011111100010000000100",
			2394 => "1111111010010110100101",
			2395 => "0011111100000000000100",
			2396 => "0000000010010110100101",
			2397 => "0000000010010110100101",
			2398 => "0001110111001000010100",
			2399 => "0001101000010000010000",
			2400 => "0000011101011100001100",
			2401 => "0000100011000000001000",
			2402 => "0001000011000100000100",
			2403 => "0000001010010110100101",
			2404 => "0000000010010110100101",
			2405 => "0000000010010110100101",
			2406 => "0000000010010110100101",
			2407 => "0000000010010110100101",
			2408 => "1111111010010110100101",
			2409 => "0001100111101000100000",
			2410 => "0010010110101000011100",
			2411 => "0001101011111100001000",
			2412 => "0000000101000100000100",
			2413 => "0000001010011001011011",
			2414 => "0000001010011001011011",
			2415 => "0010110111111000001100",
			2416 => "0000110001110100000100",
			2417 => "0000000010011001011011",
			2418 => "0001000000100000000100",
			2419 => "0000000010011001011011",
			2420 => "0000001010011001011011",
			2421 => "0001011101100000000100",
			2422 => "0000000010011001011011",
			2423 => "1111111010011001011011",
			2424 => "1111111010011001011011",
			2425 => "0011001010000000011000",
			2426 => "0010000000101000010100",
			2427 => "0000111010101100000100",
			2428 => "1111111010011001011011",
			2429 => "0010011110100000001100",
			2430 => "0001110111111000001000",
			2431 => "0011010100000000000100",
			2432 => "0000000010011001011011",
			2433 => "0000001010011001011011",
			2434 => "0000000010011001011011",
			2435 => "1111111010011001011011",
			2436 => "0000010010011001011011",
			2437 => "0001001000110100100000",
			2438 => "0001001000000100010100",
			2439 => "0011011110101100010000",
			2440 => "0001011010010100001000",
			2441 => "0000110111100000000100",
			2442 => "1111111010011001011011",
			2443 => "0000000010011001011011",
			2444 => "0001011001010100000100",
			2445 => "0000010010011001011011",
			2446 => "0000000010011001011011",
			2447 => "1111111010011001011011",
			2448 => "0010101001000100000100",
			2449 => "1111111010011001011011",
			2450 => "0010001001101000000100",
			2451 => "0000011010011001011011",
			2452 => "0000000010011001011011",
			2453 => "1111111010011001011011",
			2454 => "0000000010011001011101",
			2455 => "0000000010011001100001",
			2456 => "0000000010011001100101",
			2457 => "0000000010011001101001",
			2458 => "0000000010011001101101",
			2459 => "0000000010011001110001",
			2460 => "0000000010011001110101",
			2461 => "0000000010011001111001",
			2462 => "0000000010011001111101",
			2463 => "0000000010011010000001",
			2464 => "0000000010011010000101",
			2465 => "0000000010011010001001",
			2466 => "0000000010011010001101",
			2467 => "0000000010011010010001",
			2468 => "0000000010011010010101",
			2469 => "0000000010011010011001",
			2470 => "0000000010011010011101",
			2471 => "0000000010011010100001",
			2472 => "0011001010000000000100",
			2473 => "0000000010011010101101",
			2474 => "0000000010011010101101",
			2475 => "0001111110001100000100",
			2476 => "0000000010011010111001",
			2477 => "0000000010011010111001",
			2478 => "0001110100010100000100",
			2479 => "0000000010011011000101",
			2480 => "0000000010011011000101",
			2481 => "0001100001111000000100",
			2482 => "0000000010011011011001",
			2483 => "0011000011011100000100",
			2484 => "0000000010011011011001",
			2485 => "0000000010011011011001",
			2486 => "0001111110001100001000",
			2487 => "0010110000111000000100",
			2488 => "0000000010011011101101",
			2489 => "0000000010011011101101",
			2490 => "0000000010011011101101",
			2491 => "0001100001111000000100",
			2492 => "0000000010011100000001",
			2493 => "0001101010011000000100",
			2494 => "0000000010011100000001",
			2495 => "0000000010011100000001",
			2496 => "0001101101111100001000",
			2497 => "0001101101011100000100",
			2498 => "0000000010011100010101",
			2499 => "0000000010011100010101",
			2500 => "0000000010011100010101",
			2501 => "0001101110010100000100",
			2502 => "0000000010011100101001",
			2503 => "0001101010011000000100",
			2504 => "0000000010011100101001",
			2505 => "0000000010011100101001",
			2506 => "0001101110010100000100",
			2507 => "0000000010011100111101",
			2508 => "0001101111000000000100",
			2509 => "0000000010011100111101",
			2510 => "0000000010011100111101",
			2511 => "0001111110001100001100",
			2512 => "0011001100110000001000",
			2513 => "0010110000111000000100",
			2514 => "0000000010011101011001",
			2515 => "0000000010011101011001",
			2516 => "0000000010011101011001",
			2517 => "0000000010011101011001",
			2518 => "0001111110001100001100",
			2519 => "0011111001001000000100",
			2520 => "0000000010011101110101",
			2521 => "0011001100110000000100",
			2522 => "0000000010011101110101",
			2523 => "0000000010011101110101",
			2524 => "0000000010011101110101",
			2525 => "0001100001111000001100",
			2526 => "0001101101011100000100",
			2527 => "0000000010011110010001",
			2528 => "0001101011111100000100",
			2529 => "0000000010011110010001",
			2530 => "0000000010011110010001",
			2531 => "0000000010011110010001",
			2532 => "0001110110000100001100",
			2533 => "0011110100011000000100",
			2534 => "0000000010011110101101",
			2535 => "0001101101111100000100",
			2536 => "0000000010011110101101",
			2537 => "0000000010011110101101",
			2538 => "0000000010011110101101",
			2539 => "0001101110010100000100",
			2540 => "0000000010011111001001",
			2541 => "0001101010011000001000",
			2542 => "0001101110010100000100",
			2543 => "0000000010011111001001",
			2544 => "0000000010011111001001",
			2545 => "0000000010011111001001",
			2546 => "0001110110000100001100",
			2547 => "0001101101111100001000",
			2548 => "0001101001011000000100",
			2549 => "0000000010011111101101",
			2550 => "0000000010011111101101",
			2551 => "0000000010011111101101",
			2552 => "0001110111001000000100",
			2553 => "0000000010011111101101",
			2554 => "0000000010011111101101",
			2555 => "0001101011111100001000",
			2556 => "0001101101011100000100",
			2557 => "0000000010100000010001",
			2558 => "0000000010100000010001",
			2559 => "0011000000110000000100",
			2560 => "0000000010100000010001",
			2561 => "0010110000110000000100",
			2562 => "0000000010100000010001",
			2563 => "0000000010100000010001",
			2564 => "0001101101111100001100",
			2565 => "0011111001001000000100",
			2566 => "0000000010100000111101",
			2567 => "0001110110000100000100",
			2568 => "0000000010100000111101",
			2569 => "0000000010100000111101",
			2570 => "0001000110111100000100",
			2571 => "0000000010100000111101",
			2572 => "0001101001100100000100",
			2573 => "0000000010100000111101",
			2574 => "0000000010100000111101",
			2575 => "0011001010000000000100",
			2576 => "0000000010100001100001",
			2577 => "0010100111101100000100",
			2578 => "0000000010100001100001",
			2579 => "0011111100010000001000",
			2580 => "0010111001110100000100",
			2581 => "0000000010100001100001",
			2582 => "0000000010100001100001",
			2583 => "0000000010100001100001",
			2584 => "0001110110000100010000",
			2585 => "0011010100000000000100",
			2586 => "0000000010100010000101",
			2587 => "0001101101111100001000",
			2588 => "0001101001011000000100",
			2589 => "0000000010100010000101",
			2590 => "0000000010100010000101",
			2591 => "0000000010100010000101",
			2592 => "0000000010100010000101",
			2593 => "0001101011111100000100",
			2594 => "0000000010100010101001",
			2595 => "0001001010000100000100",
			2596 => "0000000010100010101001",
			2597 => "0011000000110000000100",
			2598 => "0000000010100010101001",
			2599 => "0010110000110000000100",
			2600 => "0000000010100010101001",
			2601 => "0000000010100010101001",
			2602 => "0011111010111100000100",
			2603 => "0000000010100011001101",
			2604 => "0011000100001000001100",
			2605 => "0011111100111000001000",
			2606 => "0001111110110000000100",
			2607 => "0000000010100011001101",
			2608 => "0000000010100011001101",
			2609 => "0000000010100011001101",
			2610 => "0000000010100011001101",
			2611 => "0001110110000100010000",
			2612 => "0001101101111100001100",
			2613 => "0001101001011000000100",
			2614 => "0000000010100011111001",
			2615 => "0010110000111000000100",
			2616 => "0000000010100011111001",
			2617 => "0000000010100011111001",
			2618 => "0000000010100011111001",
			2619 => "0010111001110100000100",
			2620 => "0000000010100011111001",
			2621 => "0000000010100011111001",
			2622 => "0001110111001000010100",
			2623 => "0000101100010100001000",
			2624 => "0001101011111100000100",
			2625 => "0000000010100100100101",
			2626 => "0000000010100100100101",
			2627 => "0000011101011100001000",
			2628 => "0000000110110100000100",
			2629 => "0000000010100100100101",
			2630 => "0000000010100100100101",
			2631 => "0000000010100100100101",
			2632 => "0000000010100100100101",
			2633 => "0001101101111100010000",
			2634 => "0011111001001000000100",
			2635 => "0000000010100101011001",
			2636 => "0001110110000100001000",
			2637 => "0010100111110100000100",
			2638 => "0000000010100101011001",
			2639 => "0000000010100101011001",
			2640 => "0000000010100101011001",
			2641 => "0010111001110100001000",
			2642 => "0011000000111000000100",
			2643 => "0000000010100101011001",
			2644 => "0000000010100101011001",
			2645 => "0000000010100101011001",
			2646 => "0000011110100000010000",
			2647 => "0011000100000000001100",
			2648 => "0011010011011100000100",
			2649 => "0000000010100110010101",
			2650 => "0001011000111000000100",
			2651 => "0000000010100110010101",
			2652 => "0000000010100110010101",
			2653 => "0000000010100110010101",
			2654 => "0011010010001000001000",
			2655 => "0001101001011000000100",
			2656 => "0000000010100110010101",
			2657 => "0000000010100110010101",
			2658 => "0010011011001100000100",
			2659 => "0000000010100110010101",
			2660 => "0000000010100110010101",
			2661 => "0001101101111100010100",
			2662 => "0011111110110000000100",
			2663 => "0000000010100111001001",
			2664 => "0010100111110100001100",
			2665 => "0001110110000100001000",
			2666 => "0010100100111100000100",
			2667 => "0000000010100111001001",
			2668 => "0000000010100111001001",
			2669 => "0000000010100111001001",
			2670 => "0000000010100111001001",
			2671 => "0001101101011000000100",
			2672 => "0000000010100111001001",
			2673 => "0000000010100111001001",
			2674 => "0011001010000000000100",
			2675 => "0000000010100111110101",
			2676 => "0001100101011100000100",
			2677 => "0000000010100111110101",
			2678 => "0001101001100100001100",
			2679 => "0001101011111100000100",
			2680 => "0000000010100111110101",
			2681 => "0001111010000000000100",
			2682 => "0000000010100111110101",
			2683 => "0000000010100111110101",
			2684 => "0000000010100111110101",
			2685 => "0000010000011000010100",
			2686 => "0011000111111000010000",
			2687 => "0010011100100000000100",
			2688 => "0000000010101000110001",
			2689 => "0010110000111000000100",
			2690 => "0000000010101000110001",
			2691 => "0000011110011100000100",
			2692 => "0000000010101000110001",
			2693 => "0000000010101000110001",
			2694 => "0000000010101000110001",
			2695 => "0001101010011000001000",
			2696 => "0001100001111000000100",
			2697 => "0000000010101000110001",
			2698 => "0000000010101000110001",
			2699 => "0000000010101000110001",
			2700 => "0000101100010100001100",
			2701 => "0001100001000100000100",
			2702 => "0000000010101001101101",
			2703 => "0010100111101100000100",
			2704 => "0000000010101001101101",
			2705 => "0000000010101001101101",
			2706 => "0011000100001000010000",
			2707 => "0000011101011100001100",
			2708 => "0001001101001100001000",
			2709 => "0000100011000000000100",
			2710 => "0000000010101001101101",
			2711 => "0000000010101001101101",
			2712 => "0000000010101001101101",
			2713 => "0000000010101001101101",
			2714 => "0000000010101001101101",
			2715 => "0000101100010100010000",
			2716 => "0001100001000100000100",
			2717 => "0000000010101010110001",
			2718 => "0010100111101100000100",
			2719 => "0000000010101010110001",
			2720 => "0000011100100000000100",
			2721 => "0000000010101010110001",
			2722 => "0000000010101010110001",
			2723 => "0001111110110000010000",
			2724 => "0000011101011100001100",
			2725 => "0001001101001100001000",
			2726 => "0000100011000000000100",
			2727 => "0000000010101010110001",
			2728 => "0000000010101010110001",
			2729 => "0000000010101010110001",
			2730 => "0000000010101010110001",
			2731 => "0000000010101010110001",
			2732 => "0011001010000000010100",
			2733 => "0011111110110000000100",
			2734 => "0000000010101011111101",
			2735 => "0010011001111000001100",
			2736 => "0001110100010100001000",
			2737 => "0011010100000000000100",
			2738 => "0000000010101011111101",
			2739 => "0000000010101011111101",
			2740 => "0000000010101011111101",
			2741 => "0000000010101011111101",
			2742 => "0010011100011000001100",
			2743 => "0001101011111100000100",
			2744 => "0000000010101011111101",
			2745 => "0001111010000000000100",
			2746 => "0000000010101011111101",
			2747 => "0000000010101011111101",
			2748 => "0010011011001100000100",
			2749 => "0000000010101011111101",
			2750 => "0000000010101011111101",
			2751 => "0010010010001100001100",
			2752 => "0000111010101100000100",
			2753 => "0000000010101101001001",
			2754 => "0001111100001000000100",
			2755 => "0000000010101101001001",
			2756 => "0000000010101101001001",
			2757 => "0001101101011000010000",
			2758 => "0000001001101000000100",
			2759 => "0000000010101101001001",
			2760 => "0011000000111000000100",
			2761 => "0000000010101101001001",
			2762 => "0001101011111100000100",
			2763 => "0000000010101101001001",
			2764 => "0000000010101101001001",
			2765 => "0000011101011100001000",
			2766 => "0000011101011100000100",
			2767 => "0000000010101101001001",
			2768 => "0000000010101101001001",
			2769 => "0000000010101101001001",
			2770 => "0001101101111100011100",
			2771 => "0011110010001000010100",
			2772 => "0001100001000100001100",
			2773 => "0000010110000000001000",
			2774 => "0000011110011100000100",
			2775 => "0000000010101110011101",
			2776 => "0000000010101110011101",
			2777 => "0000000010101110011101",
			2778 => "0000011100100000000100",
			2779 => "0000000010101110011101",
			2780 => "0000000010101110011101",
			2781 => "0010111101010100000100",
			2782 => "0000000010101110011101",
			2783 => "0000000010101110011101",
			2784 => "0000101011111000001000",
			2785 => "0010111001110100000100",
			2786 => "0000000010101110011101",
			2787 => "0000000010101110011101",
			2788 => "0011000011011100000100",
			2789 => "0000000010101110011101",
			2790 => "0000000010101110011101",
			2791 => "0000010110000000011000",
			2792 => "0010111110111100000100",
			2793 => "0000000010101111011001",
			2794 => "0001110000101000010000",
			2795 => "0000110010111100000100",
			2796 => "0000000010101111011001",
			2797 => "0011001010000000000100",
			2798 => "0000000010101111011001",
			2799 => "0001011000111100000100",
			2800 => "0000000010101111011001",
			2801 => "0000000010101111011001",
			2802 => "0000000010101111011001",
			2803 => "0000001001101000000100",
			2804 => "0000000010101111011001",
			2805 => "0000000010101111011001",
			2806 => "0001101110010100001100",
			2807 => "0001101001011000000100",
			2808 => "0000000010110000100101",
			2809 => "0011001000111000000100",
			2810 => "0000000010110000100101",
			2811 => "0000000010110000100101",
			2812 => "0011000011011100001000",
			2813 => "0000001000011000000100",
			2814 => "0000000010110000100101",
			2815 => "0000000010110000100101",
			2816 => "0011000100001000010000",
			2817 => "0011101000001100001100",
			2818 => "0000000111000000001000",
			2819 => "0000001011010100000100",
			2820 => "0000000010110000100101",
			2821 => "0000000010110000100101",
			2822 => "0000000010110000100101",
			2823 => "0000000010110000100101",
			2824 => "0000000010110000100101",
			2825 => "0000011110100000010100",
			2826 => "0011111011000000000100",
			2827 => "0000000010110001111001",
			2828 => "0011000100010100001100",
			2829 => "0001100111101000000100",
			2830 => "0000000010110001111001",
			2831 => "0001101010011000000100",
			2832 => "0000000010110001111001",
			2833 => "0000000010110001111001",
			2834 => "0000000010110001111001",
			2835 => "0001010000011100001000",
			2836 => "0010000111110100000100",
			2837 => "0000000010110001111001",
			2838 => "1111111010110001111001",
			2839 => "0010011011001100001100",
			2840 => "0011000100001000001000",
			2841 => "0001010111110000000100",
			2842 => "0000000010110001111001",
			2843 => "0000000010110001111001",
			2844 => "0000000010110001111001",
			2845 => "0000000010110001111001",
			2846 => "0010111010111000011000",
			2847 => "0011001100110000010100",
			2848 => "0001010100000000000100",
			2849 => "0000000010110010101101",
			2850 => "0001111110001100001100",
			2851 => "0001110000110000000100",
			2852 => "0000000010110010101101",
			2853 => "0010011100100000000100",
			2854 => "0000000010110010101101",
			2855 => "0000000010110010101101",
			2856 => "0000000010110010101101",
			2857 => "0000000010110010101101",
			2858 => "0000000010110010101101",
			2859 => "0010101000100100011000",
			2860 => "0010011011001100010100",
			2861 => "0011111011011100001000",
			2862 => "0000010110000000000100",
			2863 => "0000000010110100000001",
			2864 => "0000000010110100000001",
			2865 => "0000001100011100000100",
			2866 => "0000000010110100000001",
			2867 => "0001011010010100000100",
			2868 => "0000001010110100000001",
			2869 => "0000000010110100000001",
			2870 => "0000000010110100000001",
			2871 => "0001100001111000010000",
			2872 => "0001001111100000000100",
			2873 => "0000000010110100000001",
			2874 => "0011000100010100001000",
			2875 => "0000110001110100000100",
			2876 => "0000000010110100000001",
			2877 => "0000000010110100000001",
			2878 => "0000000010110100000001",
			2879 => "1111111010110100000001",
			2880 => "0010000101000100011000",
			2881 => "0001111110001100010000",
			2882 => "0011111110110000000100",
			2883 => "0000000010110101100101",
			2884 => "0010000000001000000100",
			2885 => "0000000010110101100101",
			2886 => "0010000101000100000100",
			2887 => "0000000010110101100101",
			2888 => "0000000010110101100101",
			2889 => "0001101001100100000100",
			2890 => "0000000010110101100101",
			2891 => "0000000010110101100101",
			2892 => "0001101110010100001000",
			2893 => "0001011101100000000100",
			2894 => "0000000010110101100101",
			2895 => "0000000010110101100101",
			2896 => "0000000111000000000100",
			2897 => "0000000010110101100101",
			2898 => "0010010110000000000100",
			2899 => "0000000010110101100101",
			2900 => "0001010100000000000100",
			2901 => "0000000010110101100101",
			2902 => "0001111010000000000100",
			2903 => "0000000010110101100101",
			2904 => "1111111010110101100101",
			2905 => "0000101100010100010100",
			2906 => "0001100001111000010000",
			2907 => "0000100111010000000100",
			2908 => "0000000010110110111001",
			2909 => "0001101011111100001000",
			2910 => "0000011110100000000100",
			2911 => "0000000010110110111001",
			2912 => "0000000010110110111001",
			2913 => "0000000010110110111001",
			2914 => "0000000010110110111001",
			2915 => "0000011101011100010100",
			2916 => "0011000100001000010000",
			2917 => "0010011100100000000100",
			2918 => "0000000010110110111001",
			2919 => "0001001101001100001000",
			2920 => "0000100011000000000100",
			2921 => "0000000010110110111001",
			2922 => "0000000010110110111001",
			2923 => "0000000010110110111001",
			2924 => "0000000010110110111001",
			2925 => "0000000010110110111001",
			2926 => "0001101110010100010000",
			2927 => "0011111110110000000100",
			2928 => "0000000010111000100101",
			2929 => "0000011110100000001000",
			2930 => "0001000100100000000100",
			2931 => "0000001010111000100101",
			2932 => "0000000010111000100101",
			2933 => "0000000010111000100101",
			2934 => "0001000000010000001100",
			2935 => "0001110101101100000100",
			2936 => "0000000010111000100101",
			2937 => "0011001110001100000100",
			2938 => "0000000010111000100101",
			2939 => "0000000010111000100101",
			2940 => "0010010110000000010000",
			2941 => "0010011100100000000100",
			2942 => "0000000010111000100101",
			2943 => "0011000111111000001000",
			2944 => "0000110001110100000100",
			2945 => "0000000010111000100101",
			2946 => "0000000010111000100101",
			2947 => "0000000010111000100101",
			2948 => "0010111001110100000100",
			2949 => "1111111010111000100101",
			2950 => "0010110001101000000100",
			2951 => "0000000010111000100101",
			2952 => "0000000010111000100101",
			2953 => "0010000001110000011100",
			2954 => "0011000100001000011000",
			2955 => "0011111110110000000100",
			2956 => "0000000010111001111001",
			2957 => "0000011001011000010000",
			2958 => "0010000000001000000100",
			2959 => "0000000010111001111001",
			2960 => "0001011001010100001000",
			2961 => "0000000111000000000100",
			2962 => "0000000010111001111001",
			2963 => "0000000010111001111001",
			2964 => "0000000010111001111001",
			2965 => "0000000010111001111001",
			2966 => "0000000010111001111001",
			2967 => "0001101110010100000100",
			2968 => "0000000010111001111001",
			2969 => "0011000000110000000100",
			2970 => "0000000010111001111001",
			2971 => "0010010110000000000100",
			2972 => "0000000010111001111001",
			2973 => "0000000010111001111001",
			2974 => "0010011100110100010000",
			2975 => "0011111010111100000100",
			2976 => "0000000010111011100101",
			2977 => "0010111000111100001000",
			2978 => "0010110000111000000100",
			2979 => "0000000010111011100101",
			2980 => "0000000010111011100101",
			2981 => "0000000010111011100101",
			2982 => "0010001100000100100000",
			2983 => "0011111010010100010000",
			2984 => "0010010010001100000100",
			2985 => "0000000010111011100101",
			2986 => "0001001100001100001000",
			2987 => "0001101001011000000100",
			2988 => "0000000010111011100101",
			2989 => "0000000010111011100101",
			2990 => "0000000010111011100101",
			2991 => "0001111110001100000100",
			2992 => "0000000010111011100101",
			2993 => "0001101001100100001000",
			2994 => "0011111100010100000100",
			2995 => "0000000010111011100101",
			2996 => "0000000010111011100101",
			2997 => "0000000010111011100101",
			2998 => "0010101000100100000100",
			2999 => "0000000010111011100101",
			3000 => "1111111010111011100101",
			3001 => "0001101101111100011100",
			3002 => "0001110110000100011000",
			3003 => "0001101101011100000100",
			3004 => "0000000010111100100001",
			3005 => "0010100111110100010000",
			3006 => "0001011000111100000100",
			3007 => "0000000010111100100001",
			3008 => "0010100011101000001000",
			3009 => "0001000110110100000100",
			3010 => "0000000010111100100001",
			3011 => "0000000010111100100001",
			3012 => "0000000010111100100001",
			3013 => "0000000010111100100001",
			3014 => "0000000010111100100001",
			3015 => "0000000010111100100001",
			3016 => "0001100001111000101000",
			3017 => "0000010110000000001100",
			3018 => "0011111010111100000100",
			3019 => "0000000010111110101101",
			3020 => "0011000111111000000100",
			3021 => "0000001010111110101101",
			3022 => "0000000010111110101101",
			3023 => "0011101000111000001100",
			3024 => "0001100001000100000100",
			3025 => "0000000010111110101101",
			3026 => "0001000101010100000100",
			3027 => "1111111010111110101101",
			3028 => "0000000010111110101101",
			3029 => "0000001100011100000100",
			3030 => "0000000010111110101101",
			3031 => "0011101001110000000100",
			3032 => "0000000010111110101101",
			3033 => "0000010111100100000100",
			3034 => "0000001010111110101101",
			3035 => "0000000010111110101101",
			3036 => "0000000111000000010100",
			3037 => "0001000110111000001100",
			3038 => "0011101001010000001000",
			3039 => "0000110111100000000100",
			3040 => "0000000010111110101101",
			3041 => "0000000010111110101101",
			3042 => "1111111010111110101101",
			3043 => "0011000000001100000100",
			3044 => "0000001010111110101101",
			3045 => "0000000010111110101101",
			3046 => "0000011100100000001000",
			3047 => "0010010000011000000100",
			3048 => "0000000010111110101101",
			3049 => "0000000010111110101101",
			3050 => "1111111010111110101101",
			3051 => "0010011100110100010000",
			3052 => "0011111010111100000100",
			3053 => "0000000011000000100001",
			3054 => "0010111000111100001000",
			3055 => "0010110000111000000100",
			3056 => "0000000011000000100001",
			3057 => "0000000011000000100001",
			3058 => "0000000011000000100001",
			3059 => "0010001100000100100100",
			3060 => "0001000110111000011000",
			3061 => "0001001010000100001100",
			3062 => "0011111010010100000100",
			3063 => "0000000011000000100001",
			3064 => "0001010110110100000100",
			3065 => "0000000011000000100001",
			3066 => "0000000011000000100001",
			3067 => "0010011001111000000100",
			3068 => "0000000011000000100001",
			3069 => "0011111010000100000100",
			3070 => "0000000011000000100001",
			3071 => "0000000011000000100001",
			3072 => "0011001110001100001000",
			3073 => "0011110001001000000100",
			3074 => "0000000011000000100001",
			3075 => "0000000011000000100001",
			3076 => "0000000011000000100001",
			3077 => "0010101000100100000100",
			3078 => "0000000011000000100001",
			3079 => "0000000011000000100001",
			3080 => "0011001010000000100000",
			3081 => "0010011100110100010000",
			3082 => "0011111010111100000100",
			3083 => "0000000011000010101101",
			3084 => "0001001111110000001000",
			3085 => "0001101101111100000100",
			3086 => "0000001011000010101101",
			3087 => "0000000011000010101101",
			3088 => "0000010011000010101101",
			3089 => "0011101011000100001000",
			3090 => "0000010000011000000100",
			3091 => "0000000011000010101101",
			3092 => "1111111011000010101101",
			3093 => "0001100111101000000100",
			3094 => "0000001011000010101101",
			3095 => "0000000011000010101101",
			3096 => "0000000111000000011100",
			3097 => "0011000100001000011000",
			3098 => "0011001000111000001100",
			3099 => "0010011001111000001000",
			3100 => "0011011100110000000100",
			3101 => "0000000011000010101101",
			3102 => "0000000011000010101101",
			3103 => "1111111011000010101101",
			3104 => "0010000111110100000100",
			3105 => "0000000011000010101101",
			3106 => "0000011001011000000100",
			3107 => "0000001011000010101101",
			3108 => "0000000011000010101101",
			3109 => "1111111011000010101101",
			3110 => "0001101011111100000100",
			3111 => "0000000011000010101101",
			3112 => "0010111010000000000100",
			3113 => "0000000011000010101101",
			3114 => "1111111011000010101101",
			3115 => "0000010110000000011100",
			3116 => "0011111110110000001000",
			3117 => "0001100101011100000100",
			3118 => "0000000011000100111001",
			3119 => "0000000011000100111001",
			3120 => "0011000100010100010000",
			3121 => "0000010000011000001000",
			3122 => "0011010100000000000100",
			3123 => "0000000011000100111001",
			3124 => "0000001011000100111001",
			3125 => "0011010011011100000100",
			3126 => "0000000011000100111001",
			3127 => "0000000011000100111001",
			3128 => "0000000011000100111001",
			3129 => "0000000111000000011100",
			3130 => "0010101000100100010100",
			3131 => "0011001000111000010000",
			3132 => "0000001001101000001000",
			3133 => "0011110110100100000100",
			3134 => "0000000011000100111001",
			3135 => "0000000011000100111001",
			3136 => "0011011100101100000100",
			3137 => "0000000011000100111001",
			3138 => "0000000011000100111001",
			3139 => "1111111011000100111001",
			3140 => "0011000000001100000100",
			3141 => "0000001011000100111001",
			3142 => "0000000011000100111001",
			3143 => "0001011001110000000100",
			3144 => "0000000011000100111001",
			3145 => "0010010010001100000100",
			3146 => "0000000011000100111001",
			3147 => "0010100011101000000100",
			3148 => "0000000011000100111001",
			3149 => "1111111011000100111001",
			3150 => "0010101000100100100000",
			3151 => "0010011011001100011100",
			3152 => "0011111011011100001000",
			3153 => "0000010110000000000100",
			3154 => "0000000011000110110101",
			3155 => "0000000011000110110101",
			3156 => "0000001100011100000100",
			3157 => "0000000011000110110101",
			3158 => "0001011010010100001100",
			3159 => "0010100011101000000100",
			3160 => "0000001011000110110101",
			3161 => "0010000101000100000100",
			3162 => "0000000011000110110101",
			3163 => "0000000011000110110101",
			3164 => "0000000011000110110101",
			3165 => "0000000011000110110101",
			3166 => "0010011100110100011000",
			3167 => "0001100001111000010000",
			3168 => "0001110100010100001100",
			3169 => "0011111101010100000100",
			3170 => "0000000011000110110101",
			3171 => "0001001101110100000100",
			3172 => "0000000011000110110101",
			3173 => "0000000011000110110101",
			3174 => "0000000011000110110101",
			3175 => "0011111111011100000100",
			3176 => "0000000011000110110101",
			3177 => "0000000011000110110101",
			3178 => "0001010100000000000100",
			3179 => "0000000011000110110101",
			3180 => "1111111011000110110101",
			3181 => "0001100111101000011100",
			3182 => "0000011110100000011000",
			3183 => "0001101110010100010000",
			3184 => "0011000100010100001100",
			3185 => "0011110111001000000100",
			3186 => "0000000011001001000001",
			3187 => "0010011001111000000100",
			3188 => "0000001011001001000001",
			3189 => "0000000011001001000001",
			3190 => "0000010011001001000001",
			3191 => "0000101110010000000100",
			3192 => "1111111011001001000001",
			3193 => "0000001011001001000001",
			3194 => "1111111011001001000001",
			3195 => "0001111110111100001100",
			3196 => "0000100011001000000100",
			3197 => "1111111011001001000001",
			3198 => "0011110110110100000100",
			3199 => "0000001011001001000001",
			3200 => "0000001011001001000001",
			3201 => "0010100011101000010000",
			3202 => "0010110110100100001100",
			3203 => "0010110100001000000100",
			3204 => "1111111011001001000001",
			3205 => "0000101100000000000100",
			3206 => "0000101011001001000001",
			3207 => "0000000011001001000001",
			3208 => "1111111011001001000001",
			3209 => "0011000000110000001100",
			3210 => "0000110011010000001000",
			3211 => "0000110001110100000100",
			3212 => "1111111011001001000001",
			3213 => "0000001011001001000001",
			3214 => "1111111011001001000001",
			3215 => "1111111011001001000001",
			3216 => "0001100001111000100100",
			3217 => "0000010110000000010000",
			3218 => "0011111010111100000100",
			3219 => "0000000011001011010101",
			3220 => "0001110000101000001000",
			3221 => "0001101110010100000100",
			3222 => "0000001011001011010101",
			3223 => "0000000011001011010101",
			3224 => "0000000011001011010101",
			3225 => "0011110100010000001000",
			3226 => "0010010010001100000100",
			3227 => "0000000011001011010101",
			3228 => "1111111011001011010101",
			3229 => "0000110101110100001000",
			3230 => "0011111010010100000100",
			3231 => "0000000011001011010101",
			3232 => "0000001011001011010101",
			3233 => "0000000011001011010101",
			3234 => "0001000110101100001100",
			3235 => "0000001011010100000100",
			3236 => "1111111011001011010101",
			3237 => "0011101110101000000100",
			3238 => "0000000011001011010101",
			3239 => "0000001011001011010101",
			3240 => "0001111110111100011000",
			3241 => "0010011110100000010100",
			3242 => "0011011000111100001100",
			3243 => "0001111110111100001000",
			3244 => "0011010100000000000100",
			3245 => "0000000011001011010101",
			3246 => "0000000011001011010101",
			3247 => "0000000011001011010101",
			3248 => "0000011110011100000100",
			3249 => "0000000011001011010101",
			3250 => "0000000011001011010101",
			3251 => "0000000011001011010101",
			3252 => "1111111011001011010101",
			3253 => "0000010000011000010000",
			3254 => "0011111110110000000100",
			3255 => "0000000011001101011001",
			3256 => "0001011100101000001000",
			3257 => "0011010100000000000100",
			3258 => "0000000011001101011001",
			3259 => "0000001011001101011001",
			3260 => "0000000011001101011001",
			3261 => "0000001000110000101000",
			3262 => "0001000110111000011100",
			3263 => "0001001010000100010000",
			3264 => "0011111011000000000100",
			3265 => "0000000011001101011001",
			3266 => "0001110110000100001000",
			3267 => "0010000000001000000100",
			3268 => "0000000011001101011001",
			3269 => "0000000011001101011001",
			3270 => "0000000011001101011001",
			3271 => "0001110111001000001000",
			3272 => "0000011110100000000100",
			3273 => "0000000011001101011001",
			3274 => "1111111011001101011001",
			3275 => "0000000011001101011001",
			3276 => "0011001110001100001000",
			3277 => "0000001000101100000100",
			3278 => "0000000011001101011001",
			3279 => "0000000011001101011001",
			3280 => "0000000011001101011001",
			3281 => "0001101011111100000100",
			3282 => "0000000011001101011001",
			3283 => "0001010100000000000100",
			3284 => "0000000011001101011001",
			3285 => "1111111011001101011001",
			3286 => "0000010000011000010100",
			3287 => "0000011110011100000100",
			3288 => "0000000011001111001101",
			3289 => "0011000111111000001100",
			3290 => "0011111010111100000100",
			3291 => "0000000011001111001101",
			3292 => "0011010100000000000100",
			3293 => "0000000011001111001101",
			3294 => "0000001011001111001101",
			3295 => "0000000011001111001101",
			3296 => "0010000001110000100000",
			3297 => "0011000100001000011100",
			3298 => "0011100100000000001000",
			3299 => "0001001000110100000100",
			3300 => "0000000011001111001101",
			3301 => "0000000011001111001101",
			3302 => "0000011101011100010000",
			3303 => "0001110111001000001000",
			3304 => "0001100001111000000100",
			3305 => "0000000011001111001101",
			3306 => "0000000011001111001101",
			3307 => "0000011101011100000100",
			3308 => "0000000011001111001101",
			3309 => "0000001011001111001101",
			3310 => "0000000011001111001101",
			3311 => "0000000011001111001101",
			3312 => "0001101110010100000100",
			3313 => "0000000011001111001101",
			3314 => "1111111011001111001101",
			3315 => "0000010000011000010000",
			3316 => "0011111011000000000100",
			3317 => "0000000011010001010001",
			3318 => "0001011100101000001000",
			3319 => "0011010100000000000100",
			3320 => "0000000011010001010001",
			3321 => "0000001011010001010001",
			3322 => "0000000011010001010001",
			3323 => "0000001000110000101000",
			3324 => "0010011011001100011100",
			3325 => "0010011100011000010100",
			3326 => "0001100001111000010000",
			3327 => "0011101011000100001000",
			3328 => "0011010110000100000100",
			3329 => "0000000011010001010001",
			3330 => "0000000011010001010001",
			3331 => "0001010110100100000100",
			3332 => "0000000011010001010001",
			3333 => "0000000011010001010001",
			3334 => "0000000011010001010001",
			3335 => "0011011110101100000100",
			3336 => "0000000011010001010001",
			3337 => "0000000011010001010001",
			3338 => "0010101001000100000100",
			3339 => "0000000011010001010001",
			3340 => "0010011001111100000100",
			3341 => "0000000011010001010001",
			3342 => "0000000011010001010001",
			3343 => "0001101011111100000100",
			3344 => "0000000011010001010001",
			3345 => "0001010100000000000100",
			3346 => "0000000011010001010001",
			3347 => "1111111011010001010001",
			3348 => "0001100111101000100000",
			3349 => "0010011001111000011100",
			3350 => "0011111101010100001000",
			3351 => "0001110000110000000100",
			3352 => "0000000011010011011101",
			3353 => "1111111011010011011101",
			3354 => "0000100101110100000100",
			3355 => "0000010011010011011101",
			3356 => "0011000111111000001100",
			3357 => "0001101110010100000100",
			3358 => "0000001011010011011101",
			3359 => "0000101110010000000100",
			3360 => "1111111011010011011101",
			3361 => "0000001011010011011101",
			3362 => "1111111011010011011101",
			3363 => "1111111011010011011101",
			3364 => "0001111110111100001100",
			3365 => "0000100011001000000100",
			3366 => "1111111011010011011101",
			3367 => "0011110110110100000100",
			3368 => "0000001011010011011101",
			3369 => "0000001011010011011101",
			3370 => "0011000000111000001000",
			3371 => "0010001110111100000100",
			3372 => "0000000011010011011101",
			3373 => "0000000011010011011101",
			3374 => "0001001000110100010000",
			3375 => "0001001000000100000100",
			3376 => "1111111011010011011101",
			3377 => "0010000001110000000100",
			3378 => "1111111011010011011101",
			3379 => "0010001100000100000100",
			3380 => "0000011011010011011101",
			3381 => "1111111011010011011101",
			3382 => "1111111011010011011101",
			3383 => "0000010000011000011000",
			3384 => "0011000100010100010100",
			3385 => "0000111010101100001000",
			3386 => "0001110000110000000100",
			3387 => "0000000011010101011001",
			3388 => "0000000011010101011001",
			3389 => "0001001111110000001000",
			3390 => "0000101110101000000100",
			3391 => "0000000011010101011001",
			3392 => "0000001011010101011001",
			3393 => "0000010011010101011001",
			3394 => "1111111011010101011001",
			3395 => "0010000001110000100100",
			3396 => "0011000100001000100000",
			3397 => "0011101101010100001100",
			3398 => "0010011001111000001000",
			3399 => "0000110000101000000100",
			3400 => "0000000011010101011001",
			3401 => "0000001011010101011001",
			3402 => "1111111011010101011001",
			3403 => "0000011101011100010000",
			3404 => "0000000110001000001000",
			3405 => "0010110001111100000100",
			3406 => "0000001011010101011001",
			3407 => "1111111011010101011001",
			3408 => "0000101110010000000100",
			3409 => "0000000011010101011001",
			3410 => "0000001011010101011001",
			3411 => "0000000011010101011001",
			3412 => "1111111011010101011001",
			3413 => "1111111011010101011001",
			3414 => "0001101110010100100000",
			3415 => "0001010100011000011100",
			3416 => "0000100001001000001100",
			3417 => "0000110100000000000100",
			3418 => "1111111011010111111101",
			3419 => "0000011110100000000100",
			3420 => "0000001011010111111101",
			3421 => "0000000011010111111101",
			3422 => "0000011110100000001100",
			3423 => "0000010110000000000100",
			3424 => "0000001011010111111101",
			3425 => "0001101011111100000100",
			3426 => "0000001011010111111101",
			3427 => "0000000011010111111101",
			3428 => "0000000011010111111101",
			3429 => "1111111011010111111101",
			3430 => "0010011110100000010000",
			3431 => "0000101000101000001100",
			3432 => "0001001111110100001000",
			3433 => "0000101110010000000100",
			3434 => "1111111011010111111101",
			3435 => "0000001011010111111101",
			3436 => "1111111011010111111101",
			3437 => "0000100011010111111101",
			3438 => "0001000110101100010000",
			3439 => "0010000110011000000100",
			3440 => "1111111011010111111101",
			3441 => "0011101110101000000100",
			3442 => "0000000011010111111101",
			3443 => "0010011001111100000100",
			3444 => "0000001011010111111101",
			3445 => "0000000011010111111101",
			3446 => "0010000001110000010000",
			3447 => "0010010100111100001100",
			3448 => "0000101000001100001000",
			3449 => "0001000101000000000100",
			3450 => "1111111011010111111101",
			3451 => "0000000011010111111101",
			3452 => "0000001011010111111101",
			3453 => "1111111011010111111101",
			3454 => "1111111011010111111101",
			3455 => "0001100001111000101100",
			3456 => "0000100101001000100000",
			3457 => "0010100011101000011000",
			3458 => "0011111110110000000100",
			3459 => "0000000011011010010001",
			3460 => "0000010111100100010000",
			3461 => "0010101010100000001000",
			3462 => "0010000000001000000100",
			3463 => "0000000011011010010001",
			3464 => "0000001011011010010001",
			3465 => "0001110100010100000100",
			3466 => "0000000011011010010001",
			3467 => "0000000011011010010001",
			3468 => "0000000011011010010001",
			3469 => "0001101011111100000100",
			3470 => "0000000011011010010001",
			3471 => "1111111011011010010001",
			3472 => "0001110000101000001000",
			3473 => "0000011110100000000100",
			3474 => "0000001011011010010001",
			3475 => "0000000011011010010001",
			3476 => "0000000011011010010001",
			3477 => "0000101110110100000100",
			3478 => "1111111011011010010001",
			3479 => "0011000100001000011000",
			3480 => "0000000111000000010000",
			3481 => "0010111001110100001000",
			3482 => "0011110010000100000100",
			3483 => "0000000011011010010001",
			3484 => "0000000011011010010001",
			3485 => "0010110001101000000100",
			3486 => "0000001011011010010001",
			3487 => "0000000011011010010001",
			3488 => "0010111011000100000100",
			3489 => "0000000011011010010001",
			3490 => "1111111011011010010001",
			3491 => "1111111011011010010001",
			3492 => "0001100111101000100100",
			3493 => "0000011110100000011000",
			3494 => "0000100101110100000100",
			3495 => "0000011011011100110101",
			3496 => "0000011110011100000100",
			3497 => "1111111011011100110101",
			3498 => "0000100111100000001000",
			3499 => "0001101110010100000100",
			3500 => "0000001011011100110101",
			3501 => "1111111011011100110101",
			3502 => "0000110000001100000100",
			3503 => "0000001011011100110101",
			3504 => "0000010011011100110101",
			3505 => "0000011110100000001000",
			3506 => "0000011110100000000100",
			3507 => "1111111011011100110101",
			3508 => "0000000011011100110101",
			3509 => "1111111011011100110101",
			3510 => "0001111110111100001100",
			3511 => "0000100011001000000100",
			3512 => "1111111011011100110101",
			3513 => "0010100001010100000100",
			3514 => "0000010011011100110101",
			3515 => "0000001011011100110101",
			3516 => "0001000101110000000100",
			3517 => "0000010011011100110101",
			3518 => "0001001000110100010000",
			3519 => "0001111110110000001100",
			3520 => "0011010101100100000100",
			3521 => "1111111011011100110101",
			3522 => "0010000110011100000100",
			3523 => "0000010011011100110101",
			3524 => "0001000011011100110101",
			3525 => "1111111011011100110101",
			3526 => "0001011001110000001100",
			3527 => "0011011000111000000100",
			3528 => "1111111011011100110101",
			3529 => "0001011000111100000100",
			3530 => "0000000011011100110101",
			3531 => "1111111011011100110101",
			3532 => "1111111011011100110101",
			3533 => "0001100111101000011100",
			3534 => "0010010110101000011000",
			3535 => "0000100010110100001100",
			3536 => "0001101011111100001000",
			3537 => "0000110100000000000100",
			3538 => "0000000011011111001001",
			3539 => "0000001011011111001001",
			3540 => "1111111011011111001001",
			3541 => "0011000111111000001000",
			3542 => "0001101110010100000100",
			3543 => "0000001011011111001001",
			3544 => "0000000011011111001001",
			3545 => "0000000011011111001001",
			3546 => "1111111011011111001001",
			3547 => "0001000101110000000100",
			3548 => "0000010011011111001001",
			3549 => "0000000111000000010100",
			3550 => "0011000100001000010000",
			3551 => "0011110011001000000100",
			3552 => "1111111011011111001001",
			3553 => "0000011001011000001000",
			3554 => "0001101101111100000100",
			3555 => "0000000011011111001001",
			3556 => "0000010011011111001001",
			3557 => "1111111011011111001001",
			3558 => "1111111011011111001001",
			3559 => "0001111110111100001000",
			3560 => "0000100011001000000100",
			3561 => "1111111011011111001001",
			3562 => "0000001011011111001001",
			3563 => "0011000000110000001100",
			3564 => "0011100001110100001000",
			3565 => "0011010100000000000100",
			3566 => "0000000011011111001001",
			3567 => "0000000011011111001001",
			3568 => "1111111011011111001001",
			3569 => "1111111011011111001001",
			3570 => "0001100111101000100000",
			3571 => "0000011110100000011100",
			3572 => "0011111101010100001000",
			3573 => "0001110000110000000100",
			3574 => "0000000011100001110101",
			3575 => "1111111011100001110101",
			3576 => "0001101110010100001000",
			3577 => "0001000010000000000100",
			3578 => "0000010011100001110101",
			3579 => "0000001011100001110101",
			3580 => "0001110100010100001000",
			3581 => "0001001111100000000100",
			3582 => "0000000011100001110101",
			3583 => "0000001011100001110101",
			3584 => "1111111011100001110101",
			3585 => "1111111011100001110101",
			3586 => "0001111110111100001100",
			3587 => "0011111110110000000100",
			3588 => "1111111011100001110101",
			3589 => "0000010000011000000100",
			3590 => "0000001011100001110101",
			3591 => "1111111011100001110101",
			3592 => "0011000000111000001000",
			3593 => "0010001110111100000100",
			3594 => "0000000011100001110101",
			3595 => "0000000011100001110101",
			3596 => "0001001000110100011000",
			3597 => "0001001000000100001100",
			3598 => "0011000100001000001000",
			3599 => "0011000000001100000100",
			3600 => "1111111011100001110101",
			3601 => "0000001011100001110101",
			3602 => "1111111011100001110101",
			3603 => "0011000000001100001000",
			3604 => "0011000000101000000100",
			3605 => "0000000011100001110101",
			3606 => "0000010011100001110101",
			3607 => "1111111011100001110101",
			3608 => "0011001010000000001000",
			3609 => "0011001010000000000100",
			3610 => "1111111011100001110101",
			3611 => "0000001011100001110101",
			3612 => "1111111011100001110101",
			3613 => "0011001010000000101000",
			3614 => "0011111010111100000100",
			3615 => "1111111011100101100011",
			3616 => "0000010110000000010100",
			3617 => "0000101110000100001100",
			3618 => "0010100110011000000100",
			3619 => "0000010011100101100011",
			3620 => "0000001100001000000100",
			3621 => "1111111011100101100011",
			3622 => "0000000011100101100011",
			3623 => "0000000100000100000100",
			3624 => "0000010011100101100011",
			3625 => "0000010011100101100011",
			3626 => "0010101000100100001000",
			3627 => "0001011101100000000100",
			3628 => "0000010011100101100011",
			3629 => "0000000011100101100011",
			3630 => "0001000011011000000100",
			3631 => "1111111011100101100011",
			3632 => "0000000011100101100011",
			3633 => "0001110100010100011100",
			3634 => "0010100111110100001000",
			3635 => "0000101101000100000100",
			3636 => "0000000011100101100011",
			3637 => "0000010011100101100011",
			3638 => "0000101010001000001100",
			3639 => "0010111010000000001000",
			3640 => "0001010100000000000100",
			3641 => "1111111011100101100011",
			3642 => "0000000011100101100011",
			3643 => "1111111011100101100011",
			3644 => "0000010000011000000100",
			3645 => "0000001011100101100011",
			3646 => "1111111011100101100011",
			3647 => "0000100001001000010100",
			3648 => "0010010010001100001000",
			3649 => "0001000000010100000100",
			3650 => "0000010011100101100011",
			3651 => "0000000011100101100011",
			3652 => "0011111010011100000100",
			3653 => "1111111011100101100011",
			3654 => "0001011000011000000100",
			3655 => "0000010011100101100011",
			3656 => "1111111011100101100011",
			3657 => "0010000101000100010100",
			3658 => "0001111110110000010000",
			3659 => "0000101110010000001000",
			3660 => "0010101010100000000100",
			3661 => "0000001011100101100011",
			3662 => "1111111011100101100011",
			3663 => "0011011011110100000100",
			3664 => "0000111011100101100011",
			3665 => "0000000011100101100011",
			3666 => "1111111011100101100011",
			3667 => "0011011000111100001000",
			3668 => "0001011000111000000100",
			3669 => "1111111011100101100011",
			3670 => "0000000011100101100011",
			3671 => "1111111011100101100011",
			others => (others => '0')
		);
		initial_addr_2 <= std_logic_vector(to_unsigned(1192, initial_addr_2'length));
		initial_addr_3 <= std_logic_vector(to_unsigned(2454, initial_addr_3'length));
	end generate gen_rom_15;

	process (Clk)
	begin
		if rising_edge(Clk) then
			if (Re = '1') then
				-- Read from Addr
				Dout <= bank(to_integer(unsigned(Addr)));
			else
				Dout <= (others => '0');
			end if;
		end if;
	end process;
end Behavioral;
