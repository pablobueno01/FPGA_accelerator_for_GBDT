-------------------------------------------------------------------------------
-- VHDL test file for 'image.vhd'
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 13;
            NUM_FEATURES:  positive := 16);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
            --  Load_trees: in std_logic;
            --  Valid_node: in std_logic;
            --  Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
            --  Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    -- signal Load_trees:    std_logic := '0';
    -- signal Valid_node:    std_logic := '0';
    -- signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
    --                                        0) := (others => '0');
    -- signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 --Load_trees    => Load_trees,
                 --Valid_node    => Valid_node,
                 --Addr          => Addr,
                 --Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        
        
        -- LOAD FEATURES
        -----------------------------------------------------------------------
        

		-- PIXELS OF CLASS 0
		---------------------
		class_label <= std_logic_vector(to_unsigned(0, class_label'length));

		-- PIXEL 0
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000100111010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 1
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000011010101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000001111001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 2
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000101000111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 3
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100001101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 4
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 5
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 6
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000101001000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 7
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 8
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 9
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 10
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 11
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101000011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 12
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000101000001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 13
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 14
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100100100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000010001000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 15
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100001001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001001010";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 16
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 17
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000100100010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 18
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100100000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 19
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 20
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100100010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 21
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 22
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 23
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 24
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 25
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 26
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000101001010";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011001011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 27
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 28
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100111000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 29
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001001101";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 30
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 31
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000011101101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001111110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 32
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 33
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 34
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101001010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 35
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000001001111";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 36
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 37
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 38
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 39
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000101000101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 40
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000100011101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 41
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 42
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000000";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 43
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001001010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 44
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 45
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 46
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 47
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100110011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 48
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 49
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 50
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 51
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 52
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 53
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101001000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 54
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001010011";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 55
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 56
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011101001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000011011110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010000101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000001110010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 57
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 58
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 59
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100000111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 60
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 61
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100000011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000001111001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 62
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000010010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000001100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000001101110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 63
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 64
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100011000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 65
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 66
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 67
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 68
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 69
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100111000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 70
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100100001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 71
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000011010010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010000010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000001110001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 72
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 73
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 74
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100100001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 75
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 76
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 77
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 78
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000001010110";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 79
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000011000111";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 80
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 81
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101011000";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000011010001";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 82
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000101001001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 83
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 84
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001111011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000001101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 85
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111011";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 86
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 87
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 88
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 89
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100100010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 90
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100111100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 91
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000100100000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000001010000";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 92
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101010000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011001101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 93
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000001001111";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 94
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 95
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100110010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 96
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 97
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100110011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 98
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000001011";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000010100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000001110011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000001011111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 99
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 100
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100001001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 101
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100111101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 102
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000101001111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011001101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 103
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 104
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 105
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 106
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001110110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000001100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 107
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100010011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 108
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000001111";
		wait for Clk_period;
		Features_din <= "0000000100110011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 109
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 110
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000011010011";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 111
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100010001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010000010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 112
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100111111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000011000000";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 113
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100011000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 114
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000011111000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000001111101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 115
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 116
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001111111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001101111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 117
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 118
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100011011";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001101";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 119
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 120
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 121
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 122
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000011111011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010001011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 123
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001111000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 124
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 125
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000100110011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 126
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011001100";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 127
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000101010001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000011011000";
		wait for Clk_period;
		Features_din <= "0000000001010010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 128
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100010110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 129
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100111011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 130
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000101001000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 131
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000100010101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010001011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 132
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 133
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101100011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101010101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011010100";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 134
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 135
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100001110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000001010000";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 136
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100011011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010000111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 137
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 138
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100001110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 139
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 140
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 141
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 142
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 143
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 144
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 145
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 146
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100111010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011001100";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 147
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 148
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 149
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000011000001";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 150
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011111111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000011110100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000001111110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 151
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100010000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 152
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000101000011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 153
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100111111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 154
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 155
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001001111";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 156
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 157
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 158
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 159
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011001111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 160
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100011101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 161
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011100010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000011011000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010001011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000001111010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010011000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 162
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 163
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 164
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 165
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100111011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 166
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011000000";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 167
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 168
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 169
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 170
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 171
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100111100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000011000111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 172
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 173
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 174
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100010101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 175
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100010010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 176
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101001010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 177
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100110010";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 178
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101100011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101010111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 179
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100001011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 180
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 181
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 182
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 183
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 184
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 185
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010000100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 186
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 187
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 188
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100101101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 189
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100100011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 190
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 191
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100111010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 192
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100000000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001111011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 193
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010001";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 194
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100010111";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000001010100";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 195
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100001001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 196
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100111010";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000011000000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 197
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000001111111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 198
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 199
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101000101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 200
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000101000111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 201
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000010110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001110111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000001100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 202
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 203
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 204
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 205
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101001110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000011001100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 206
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 207
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 208
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 209
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 210
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000011111010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 211
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 212
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 213
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 214
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000101001000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 215
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 216
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 217
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 218
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 219
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100010010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 220
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101100001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101010011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011001111";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 221
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100010010";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010000101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 222
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 223
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100111010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 224
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 225
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 226
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 227
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 228
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 229
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000011111101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000001111011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 230
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 231
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 232
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000101001110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000011001101";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 233
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 234
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 235
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100000010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 236
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 237
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 238
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000101001000";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001001010";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 239
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100010110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001001010";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 240
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 241
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 242
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100000010";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010000000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 243
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 244
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 245
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000010";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 246
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000101001011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 247
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100100010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 248
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101101";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000001010001";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 249
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 250
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 251
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 252
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 253
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 254
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 255
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 256
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 257
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 258
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000100011011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010001010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 259
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 260
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 261
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 262
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000001111";
		wait for Clk_period;
		Features_din <= "0000000101000111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000011001011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 263
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000001010001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 264
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 265
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100011101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 266
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100100110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 267
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000011110010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 268
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010001";
		wait for Clk_period;
		Features_din <= "0000000100010100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010000101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 269
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101001001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000011000111";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 270
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 271
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 272
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000100100001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 273
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 274
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100000011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010000110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 275
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101001110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000011010000";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 276
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 277
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 278
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000001101100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000001011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000001111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 279
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000011000111";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 280
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100000001";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000001111010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 281
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 282
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 283
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011111010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000011110000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000001111110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 284
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000001010001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 285
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000101000110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011001110";
		wait for Clk_period;
		Features_din <= "0000000001010000";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 286
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100001011";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000010001010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 287
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000001110011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000001100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000001111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 288
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100000010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000001110110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010100101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 289
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 290
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000001111";
		wait for Clk_period;
		Features_din <= "0000000011101010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000010000001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010010110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 291
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100111101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 292
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010111000";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 293
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 294
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 295
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100100010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 296
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 297
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 298
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001001101";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 299
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000101000110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000011000100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 300
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 301
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000011011100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000010001011";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000001110110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010011101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 302
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100001110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 303
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000011001010";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 304
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011000";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 305
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 306
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101000001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010100110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 307
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000010010100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 308
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000010110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000010100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010000010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001110000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 309
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101000000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 310
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010111101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 311
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 312
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000010001110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 313
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100000110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010100010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 314
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 315
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 316
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 317
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101001010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000011010000";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010110001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 318
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100001101";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 319
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100010110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 320
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100001011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 321
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001001010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 322
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100010000";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010101100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 323
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100001111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010010110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 324
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 325
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010111110";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 326
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100111011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 327
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100011010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010101111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 328
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 329
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101011011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000101001100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001001110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 330
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 331
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 332
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000010111011";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 333
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101101000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000101011000";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011010100";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011101110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 334
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100111100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 335
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100011001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 336
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000100100011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010111001";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010011011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 337
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010100000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 338
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100011011";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000011";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 339
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010111011";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 340
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100100101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 341
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101000010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011001000";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000010101001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 342
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100100000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 343
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 344
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100111001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011000001";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 345
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100100111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 346
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000100111000";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000011000001";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 347
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000010011100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 348
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000100011111";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000010110000";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 349
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000100110100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000011000011";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 350
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100011110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010001101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 351
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000101000011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 352
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100101111";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000001001001";
		wait for Clk_period;
		Features_din <= "0000000010101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010010101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 353
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101011";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000010110010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 354
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000100111110";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 355
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000101000111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010111010";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 356
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000100111100";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010111111";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000010100011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 357
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100010011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010100001";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010001000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 358
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100010000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010011111";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010000111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 359
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000100101001";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 360
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010110011";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010011001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 361
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000011010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010101";
		wait for Clk_period;
		Features_din <= "0000000011001110";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000001111101";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000001101100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010001010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 362
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101101001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000101011001";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000011011000";
		wait for Clk_period;
		Features_din <= "0000000001001011";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000010110110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011110000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 363
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100101001";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100011101";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000001011100";
		wait for Clk_period;
		Features_din <= "0000000010100101";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000001010010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 364
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100010110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 365
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000100110010";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000011000101";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 366
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000111110";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001001000";
		wait for Clk_period;
		Features_din <= "0000000010110111";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011010";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 367
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000101001001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001000101";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010101000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011100011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 368
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101001110";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000101000001";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000011000110";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000010100111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 369
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110100";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010110";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010110101";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 370
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101000010";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000100110110";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010111100";
		wait for Clk_period;
		Features_din <= "0000000001000110";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010011110";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011010011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 371
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011000";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010101010";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010010011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 372
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100000011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000011111000";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000001000100";
		wait for Clk_period;
		Features_din <= "0000000010001100";
		wait for Clk_period;
		Features_din <= "0000000000110001";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000100100";
		wait for Clk_period;
		Features_din <= "0000000000111010";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000001110111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010011110";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 373
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100100111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100011100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000010101101";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100011";
		wait for Clk_period;
		Features_din <= "0000000000110011";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000000011000";
		wait for Clk_period;
		Features_din <= "0000000010001111";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000001";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 374
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010011";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101000100";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000110101";
		wait for Clk_period;
		Features_din <= "0000000001000010";
		wait for Clk_period;
		Features_din <= "0000000011000010";
		wait for Clk_period;
		Features_din <= "0000000001001100";
		wait for Clk_period;
		Features_din <= "0000000000110110";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000001000001";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 375
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010111";
		wait for Clk_period;
		Features_din <= "0000000100101000";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000001000000";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000010010001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000100";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 376
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100110111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010110100";
		wait for Clk_period;
		Features_din <= "0000000000111101";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011111";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010011000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011001000";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 377
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100011101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100010010";
		wait for Clk_period;
		Features_din <= "0000000000101101";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000110100";
		wait for Clk_period;
		Features_din <= "0000000010100100";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000110010";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011101";
		wait for Clk_period;
		Features_din <= "0000000000011100";
		wait for Clk_period;
		Features_din <= "0000000010001001";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010111011";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 378
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000101010101";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000101000111";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101001";
		wait for Clk_period;
		Features_din <= "0000000000111011";
		wait for Clk_period;
		Features_din <= "0000000011001001";
		wait for Clk_period;
		Features_din <= "0000000001000111";
		wait for Clk_period;
		Features_din <= "0000000000101110";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000111000";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000000100111";
		wait for Clk_period;
		Features_din <= "0000000000100110";
		wait for Clk_period;
		Features_din <= "0000000010101011";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011011111";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 379
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100111000";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000010011";
		wait for Clk_period;
		Features_din <= "0000000100101010";
		wait for Clk_period;
		Features_din <= "0000000000101111";
		wait for Clk_period;
		Features_din <= "0000000000101010";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000010101110";
		wait for Clk_period;
		Features_din <= "0000000000111001";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000100101";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000011010";
		wait for Clk_period;
		Features_din <= "0000000000011011";
		wait for Clk_period;
		Features_din <= "0000000000011110";
		wait for Clk_period;
		Features_din <= "0000000010010000";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000011000101";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXEL 380
		-- Load and valid features flags
		Load_features <= '1';
		Valid_feature <= '1';

		Features_din <= "0000000100010111";
		wait for Clk_period;

		-- Reset load flag
		Load_features <= '0';

		Features_din <= "0000000000011001";
		wait for Clk_period;
		Features_din <= "0000000100001100";
		wait for Clk_period;
		Features_din <= "0000000000110000";
		wait for Clk_period;
		Features_din <= "0000000000101100";
		wait for Clk_period;
		Features_din <= "0000000000111111";
		wait for Clk_period;
		Features_din <= "0000000010011101";
		wait for Clk_period;
		Features_din <= "0000000000111100";
		wait for Clk_period;
		Features_din <= "0000000000101000";
		wait for Clk_period;
		Features_din <= "0000000000101011";
		wait for Clk_period;
		Features_din <= "0000000000110111";
		wait for Clk_period;
		Features_din <= "0000000000100001";
		wait for Clk_period;
		Features_din <= "0000000000100010";
		wait for Clk_period;
		Features_din <= "0000000000100000";
		wait for Clk_period;
		Features_din <= "0000000010000100";
		wait for Clk_period;

		last_feature <= '1';
		pc_count     <= '1'; -- count pixel
		Features_din <= "0000000010110010";
		wait for Clk_period;

		-- Reset count, last and valid flags
		pc_count      <= '0';
		Last_feature  <= '0';
		Valid_feature <= '0';

		-- Wait until inference is complete
		wait until Finish = '1';

		wait for Clk_period * 1/2;

		if Dout = class_label then
			hc_count <= '1';
		end if;

		wait for Clk_period;
		hc_count <= '0';

		-- PIXELS OF CLASS 1
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(1, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 2
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(2, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 3
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(3, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000101001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 4
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(4, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000101010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000101010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 5
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(5, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000101001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000101011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000110000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000101001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000101001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000101011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100111101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000101010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 6
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(6, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000101000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000101010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000101001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000101010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000101100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000101010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000100011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000101100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000100110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000101011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000101001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 7
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(7, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 202
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 203
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 204
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 205
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 206
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 207
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 208
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 209
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 210
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 211
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 212
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 213
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 214
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 215
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 8
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(8, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 202
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 203
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 204
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 205
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 206
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 207
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 208
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 209
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 210
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 211
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 212
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 213
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 214
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 215
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 216
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 217
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 218
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 219
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 220
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 221
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 222
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 223
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 224
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 225
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 226
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 227
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 228
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 229
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 230
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 231
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 232
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 233
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 234
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 235
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 236
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 237
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 238
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 239
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 240
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 241
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 242
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 243
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 244
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 245
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 246
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 247
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 248
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 249
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 250
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 251
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 252
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 253
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000100001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 254
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 255
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 256
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 257
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 258
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 259
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 9
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(9, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "1111111111111100";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "1111111111111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "1111111111111100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "1111111111111110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 10
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(10, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011000100";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000011000001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000100001110";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001110";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000011000011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011010000";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000100000001";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000011010001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010101110";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000011000101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011001100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011101011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011110111";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010101101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011100101";
--		wait for Clk_period;
--		Features_din <= "0000000010110000";
--		wait for Clk_period;
--		Features_din <= "0000000011001000";
--		wait for Clk_period;
--		Features_din <= "0000000011111010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000010111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011101";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000010100001";
--		wait for Clk_period;
--		Features_din <= "0000000011001010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100111";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000011011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011110011";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000010110011";
--		wait for Clk_period;
--		Features_din <= "0000000011001011";
--		wait for Clk_period;
--		Features_din <= "0000000011111101";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000010111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011010110";
--		wait for Clk_period;
--		Features_din <= "0000000010101000";
--		wait for Clk_period;
--		Features_din <= "0000000011000010";
--		wait for Clk_period;
--		Features_din <= "0000000011110010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000010110111";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011010111";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000011011100";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000010100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010110101";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011001001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011100010";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000010010011";
--		wait for Clk_period;
--		Features_din <= "0000000010111100";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000010000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000100001010";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000010001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--		Features_din <= "0000000010000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110110";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--		Features_din <= "0000000011010011";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000100000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011110101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 202
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000010011110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 203
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 204
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011011001";
--		wait for Clk_period;
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--		Features_din <= "0000000010110100";
--		wait for Clk_period;
--		Features_din <= "0000000011100000";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 205
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000011010100";
--		wait for Clk_period;
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010100101";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 206
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000011000111";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 207
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000011001101";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000010111011";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 208
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000011001111";
--		wait for Clk_period;
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101111";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000010000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 209
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000011110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000011100110";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--		Features_din <= "0000000010001011";
--		wait for Clk_period;
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000010000011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 11
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(11, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000001111100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000010001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000010000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000000001";
--		wait for Clk_period;
--		Features_din <= "1111111111111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000010100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000001100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000001011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "1111111111111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "1111111111111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001110010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000010011001";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "1111111111111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "1111111111111101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000010011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "1111111111111101";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001111000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 202
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 203
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 204
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 205
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 206
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 207
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 208
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 209
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000010001010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 210
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 211
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 212
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 213
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 214
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 215
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 216
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 217
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 218
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 219
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 220
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000010000010";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--		Features_din <= "0000000001000010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 221
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 222
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000001000011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 223
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 224
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 225
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 226
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 227
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 228
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 229
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000000100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 230
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000010010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000010";
--		wait for Clk_period;
--		Features_din <= "0000000010001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000001011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 231
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 232
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 233
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 234
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000111110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 235
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 236
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 237
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 238
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 239
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000001001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 240
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 241
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001000110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 242
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001110101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001110000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 243
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000001000100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 244
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000001101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 245
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001000000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000111100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 246
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001001000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000001000101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 247
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001011000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000001010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000111011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 248
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 249
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 250
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 251
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000001010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000001010000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXELS OF CLASS 12
--		---------------------
--		class_label <= std_logic_vector(to_unsigned(12, class_label'length));
--
--		-- PIXEL 0
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 1
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 2
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 3
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 4
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 5
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 6
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 7
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 8
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 9
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 10
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 11
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 12
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 13
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 14
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 15
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 16
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 17
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 18
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 19
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 20
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 21
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 22
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 23
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 24
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 25
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 26
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 27
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 28
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 29
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 30
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 31
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 32
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 33
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 34
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 35
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 36
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 37
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 38
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 39
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 40
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 41
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 42
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 43
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 44
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 45
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 46
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 47
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 48
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 49
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 50
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 51
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 52
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 53
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 54
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 55
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 56
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 57
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 58
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 59
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 60
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 61
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 62
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 63
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 64
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 65
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 66
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 67
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 68
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 69
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 70
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 71
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 72
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 73
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 74
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 75
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 76
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 77
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 78
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 79
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 80
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 81
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 82
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 83
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 84
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 85
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 86
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 87
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 88
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 89
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 90
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 91
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 92
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 93
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 94
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 95
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 96
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 97
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 98
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 99
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 100
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 101
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 102
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 103
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 104
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 105
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 106
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 107
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 108
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 109
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 110
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 111
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 112
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 113
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 114
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 115
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 116
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 117
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 118
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 119
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 120
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 121
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 122
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 123
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 124
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 125
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 126
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 127
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 128
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 129
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 130
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 131
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 132
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 133
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 134
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 135
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 136
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 137
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 138
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 139
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 140
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 141
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 142
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 143
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 144
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 145
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 146
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 147
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 148
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 149
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 150
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 151
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 152
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 153
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 154
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 155
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 156
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 157
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 158
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 159
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 160
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 161
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 162
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 163
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 164
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 165
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 166
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 167
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 168
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 169
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 170
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 171
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 172
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 173
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 174
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 175
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 176
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 177
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 178
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 179
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 180
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 181
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 182
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 183
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 184
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 185
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 186
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 187
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 188
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 189
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 190
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 191
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 192
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 193
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 194
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 195
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 196
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 197
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 198
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 199
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 200
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 201
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 202
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 203
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 204
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 205
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 206
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 207
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 208
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 209
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 210
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 211
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 212
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 213
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 214
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 215
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 216
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 217
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 218
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 219
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 220
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 221
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 222
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 223
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 224
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 225
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 226
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 227
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 228
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 229
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 230
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 231
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 232
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 233
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 234
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 235
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 236
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 237
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 238
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 239
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000111010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000111101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 240
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 241
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 242
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 243
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 244
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 245
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 246
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 247
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 248
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 249
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 250
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 251
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 252
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 253
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 254
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 255
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 256
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 257
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 258
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 259
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 260
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 261
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 262
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 263
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 264
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 265
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 266
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 267
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 268
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 269
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 270
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 271
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 272
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 273
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 274
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 275
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 276
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 277
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 278
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 279
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 280
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 281
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 282
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 283
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 284
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 285
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 286
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 287
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 288
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 289
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 290
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 291
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 292
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 293
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 294
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 295
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 296
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 297
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 298
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 299
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 300
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 301
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 302
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 303
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 304
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 305
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 306
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 307
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 308
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 309
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 310
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 311
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 312
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 313
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 314
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 315
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 316
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 317
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 318
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 319
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 320
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 321
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 322
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 323
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 324
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 325
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 326
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 327
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 328
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 329
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 330
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 331
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 332
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 333
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 334
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 335
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 336
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 337
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 338
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 339
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 340
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 341
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 342
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 343
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 344
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 345
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 346
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 347
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 348
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 349
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 350
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 351
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 352
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 353
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 354
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 355
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 356
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 357
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 358
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 359
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 360
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 361
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 362
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 363
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 364
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 365
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 366
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 367
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 368
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 369
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 370
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 371
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 372
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 373
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 374
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 375
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 376
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 377
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 378
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 379
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 380
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 381
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 382
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 383
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 384
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 385
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 386
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 387
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 388
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 389
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 390
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 391
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 392
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 393
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 394
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 395
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 396
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 397
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 398
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 399
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 400
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 401
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 402
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 403
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 404
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 405
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 406
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 407
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 408
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 409
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 410
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 411
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 412
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 413
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 414
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 415
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 416
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 417
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 418
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 419
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 420
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000110";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 421
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000111000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 422
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 423
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 424
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 425
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 426
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 427
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 428
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 429
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 430
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 431
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 432
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 433
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 434
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 435
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 436
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 437
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 438
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 439
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 440
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 441
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 442
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 443
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 444
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 445
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000110100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101101";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 446
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 447
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110101";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 448
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 449
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 450
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000110110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000110010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 451
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 452
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 453
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 454
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 455
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000001100";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 456
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000001001";
--		wait for Clk_period;
--		Features_din <= "0000000000001000";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000001011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 457
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100111";
--		wait for Clk_period;
--		Features_din <= "0000000000110000";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 458
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000001101";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 459
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000101110";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011101";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 460
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000001110";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000010111";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000011110";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 461
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--		Features_din <= "0000000000110111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000110011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--		Features_din <= "0000000000101000";
--		wait for Clk_period;
--		Features_din <= "0000000000100010";
--		wait for Clk_period;
--		Features_din <= "0000000000100110";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100100";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 462
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000000111";
--		wait for Clk_period;
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--		Features_din <= "0000000000001111";
--		wait for Clk_period;
--		Features_din <= "0000000000010000";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000010100";
--		wait for Clk_period;
--		Features_din <= "0000000000101010";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000010010";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011100";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000010101";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000010011";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
--		-- PIXEL 463
--		-- Load and valid features flags
--		Load_features <= '1';
--		Valid_feature <= '1';
--
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset load flag
--		Load_features <= '0';
--
--		Features_din <= "0000000000010001";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000011000";
--		wait for Clk_period;
--		Features_din <= "0000000000010110";
--		wait for Clk_period;
--		Features_din <= "0000000000011010";
--		wait for Clk_period;
--		Features_din <= "0000000000011111";
--		wait for Clk_period;
--		Features_din <= "0000000000101111";
--		wait for Clk_period;
--		Features_din <= "0000000000100101";
--		wait for Clk_period;
--		Features_din <= "0000000000101011";
--		wait for Clk_period;
--		Features_din <= "0000000000011001";
--		wait for Clk_period;
--		Features_din <= "0000000000100001";
--		wait for Clk_period;
--		Features_din <= "0000000000100011";
--		wait for Clk_period;
--		Features_din <= "0000000000011011";
--		wait for Clk_period;
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		last_feature <= '1';
--		pc_count     <= '1'; -- count pixel
--		Features_din <= "0000000000100000";
--		wait for Clk_period;
--
--		-- Reset count, last and valid flags
--		pc_count      <= '0';
--		Last_feature  <= '0';
--		Valid_feature <= '0';
--
--		-- Wait until inference is complete
--		wait until Finish = '1';
--
--		wait for Clk_period * 1/2;
--
--		if Dout = class_label then
--			hc_count <= '1';
--		end if;
--
--		wait for Clk_period;
--		hc_count <= '0';
--
		wait;
	end process;
end;
